
module mult_N128_CC1 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
         n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
         n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041,
         n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
         n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057,
         n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
         n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
         n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081,
         n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
         n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097,
         n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
         n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
         n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
         n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129,
         n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
         n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
         n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153,
         n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
         n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
         n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177,
         n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185,
         n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
         n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201,
         n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
         n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217,
         n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
         n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233,
         n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241,
         n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249,
         n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257,
         n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
         n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273,
         n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
         n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289,
         n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297,
         n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305,
         n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313,
         n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321,
         n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329,
         n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337,
         n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345,
         n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353,
         n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361,
         n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369,
         n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377,
         n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385,
         n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393,
         n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401,
         n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409,
         n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417,
         n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
         n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433,
         n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441,
         n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449,
         n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457,
         n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465,
         n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473,
         n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481,
         n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489,
         n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497,
         n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505,
         n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513,
         n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521,
         n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529,
         n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537,
         n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545,
         n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553,
         n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561,
         n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569,
         n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577,
         n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585,
         n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593,
         n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601,
         n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609,
         n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617,
         n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625,
         n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633,
         n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641,
         n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649,
         n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657,
         n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665,
         n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673,
         n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681,
         n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689,
         n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697,
         n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705,
         n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713,
         n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721,
         n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729,
         n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737,
         n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745,
         n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753,
         n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761,
         n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769,
         n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777,
         n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
         n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793,
         n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801,
         n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809,
         n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817,
         n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825,
         n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833,
         n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
         n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849,
         n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
         n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865,
         n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873,
         n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
         n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889,
         n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897,
         n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905,
         n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
         n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921,
         n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929,
         n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937,
         n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945,
         n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953,
         n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961,
         n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969,
         n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977,
         n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985,
         n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993,
         n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
         n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
         n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017,
         n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025,
         n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033,
         n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041,
         n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049,
         n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057,
         n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065,
         n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073,
         n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081,
         n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089,
         n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097,
         n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105,
         n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113,
         n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121,
         n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
         n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137,
         n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145,
         n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153,
         n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161,
         n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169,
         n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177,
         n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185,
         n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193,
         n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201,
         n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209,
         n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217,
         n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225,
         n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233,
         n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241,
         n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249,
         n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257,
         n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265,
         n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273,
         n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281,
         n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289,
         n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297,
         n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305,
         n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313,
         n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321,
         n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329,
         n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337,
         n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
         n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353,
         n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
         n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369,
         n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377,
         n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385,
         n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393,
         n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401,
         n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409,
         n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
         n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425,
         n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
         n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441,
         n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449,
         n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457,
         n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465,
         n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473,
         n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481,
         n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
         n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497,
         n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
         n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513,
         n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521,
         n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529,
         n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537,
         n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545,
         n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553,
         n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
         n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569,
         n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577,
         n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585,
         n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593,
         n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601,
         n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609,
         n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617,
         n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625,
         n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
         n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641,
         n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649,
         n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657,
         n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665,
         n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673,
         n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681,
         n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689,
         n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697,
         n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
         n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713,
         n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721,
         n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729,
         n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737,
         n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745,
         n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753,
         n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761,
         n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769,
         n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
         n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785,
         n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
         n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801,
         n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809,
         n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817,
         n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825,
         n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833,
         n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841,
         n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
         n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857,
         n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865,
         n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873,
         n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881,
         n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889,
         n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897,
         n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905,
         n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913,
         n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
         n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929,
         n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
         n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945,
         n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953,
         n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961,
         n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969,
         n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977,
         n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985,
         n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993,
         n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001,
         n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009,
         n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017,
         n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025,
         n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033,
         n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041,
         n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049,
         n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057,
         n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065,
         n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073,
         n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
         n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089,
         n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097,
         n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105,
         n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113,
         n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121,
         n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129,
         n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137,
         n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145,
         n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153,
         n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161,
         n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169,
         n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177,
         n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185,
         n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193,
         n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201,
         n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209,
         n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217,
         n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225,
         n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233,
         n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241,
         n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
         n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257,
         n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265,
         n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273,
         n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281,
         n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289,
         n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297,
         n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305,
         n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313,
         n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
         n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329,
         n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337,
         n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345,
         n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353,
         n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361,
         n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369,
         n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377,
         n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385,
         n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393,
         n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401,
         n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409,
         n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417,
         n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425,
         n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433,
         n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
         n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449,
         n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457,
         n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465,
         n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473,
         n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481,
         n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489,
         n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497,
         n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505,
         n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
         n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521,
         n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529,
         n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
         n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545,
         n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553,
         n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561,
         n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
         n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577,
         n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
         n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593,
         n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601,
         n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
         n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
         n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625,
         n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633,
         n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
         n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649,
         n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657,
         n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665,
         n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673,
         n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681,
         n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689,
         n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697,
         n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705,
         n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713,
         n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721,
         n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729,
         n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737,
         n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745,
         n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753,
         n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761,
         n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769,
         n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777,
         n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785,
         n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793,
         n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801,
         n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809,
         n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817,
         n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825,
         n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833,
         n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841,
         n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849,
         n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857,
         n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865,
         n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873,
         n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881,
         n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889,
         n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897,
         n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905,
         n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913,
         n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921,
         n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929,
         n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937,
         n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945,
         n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953,
         n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961,
         n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969,
         n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977,
         n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985,
         n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993,
         n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
         n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009,
         n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017,
         n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025,
         n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033,
         n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041,
         n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049,
         n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057,
         n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065,
         n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073,
         n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081,
         n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089,
         n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097,
         n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105,
         n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113,
         n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121,
         n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129,
         n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137,
         n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145,
         n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153,
         n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161,
         n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169,
         n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177,
         n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185,
         n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193,
         n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201,
         n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209,
         n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217,
         n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225,
         n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233,
         n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241,
         n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249,
         n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257,
         n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265,
         n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273,
         n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281,
         n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289,
         n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297,
         n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305,
         n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313,
         n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321,
         n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329,
         n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337,
         n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345,
         n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353,
         n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361,
         n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369,
         n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377,
         n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385,
         n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393,
         n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401,
         n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409,
         n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417,
         n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425,
         n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
         n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441,
         n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449,
         n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457,
         n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465,
         n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473,
         n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481,
         n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489,
         n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497,
         n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505,
         n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513,
         n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521,
         n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529,
         n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537,
         n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545,
         n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553,
         n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561,
         n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569,
         n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577,
         n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585,
         n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593,
         n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601,
         n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609,
         n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617,
         n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625,
         n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633,
         n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641,
         n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649,
         n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657,
         n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665,
         n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673,
         n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681,
         n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689,
         n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697,
         n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705,
         n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713,
         n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721,
         n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729,
         n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737,
         n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745,
         n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753,
         n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761,
         n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769,
         n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777,
         n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785,
         n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793,
         n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801,
         n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809,
         n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817,
         n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825,
         n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833,
         n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841,
         n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849,
         n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857,
         n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865,
         n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873,
         n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
         n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889,
         n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897,
         n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905,
         n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913,
         n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921,
         n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929,
         n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
         n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945,
         n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953,
         n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961,
         n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969,
         n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977,
         n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985,
         n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993,
         n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001,
         n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009,
         n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017,
         n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025,
         n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033,
         n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041,
         n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049,
         n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057,
         n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065,
         n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073,
         n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081,
         n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089,
         n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097,
         n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105,
         n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113,
         n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121,
         n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129,
         n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137,
         n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145,
         n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153,
         n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161,
         n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169,
         n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177,
         n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185,
         n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193,
         n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201,
         n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209,
         n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217,
         n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225,
         n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233,
         n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
         n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249,
         n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257,
         n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265,
         n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273,
         n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281,
         n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289,
         n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297,
         n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305,
         n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
         n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321,
         n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329,
         n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337,
         n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345,
         n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353,
         n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361,
         n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369,
         n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377,
         n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
         n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393,
         n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401,
         n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409,
         n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417,
         n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425,
         n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433,
         n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441,
         n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449,
         n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
         n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465,
         n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473,
         n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481,
         n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489,
         n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497,
         n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505,
         n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513,
         n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521,
         n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
         n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537,
         n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545,
         n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
         n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561,
         n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569,
         n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577,
         n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585,
         n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593,
         n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
         n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609,
         n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617,
         n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625,
         n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633,
         n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641,
         n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649,
         n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657,
         n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665,
         n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
         n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681,
         n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689,
         n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697,
         n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705,
         n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713,
         n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721,
         n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729,
         n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737,
         n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
         n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753,
         n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761,
         n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769,
         n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777,
         n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785,
         n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793,
         n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801,
         n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809,
         n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817,
         n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825,
         n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833,
         n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841,
         n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849,
         n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857,
         n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865,
         n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873,
         n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881,
         n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889,
         n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897,
         n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905,
         n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913,
         n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921,
         n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929,
         n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937,
         n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945,
         n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953,
         n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961,
         n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969,
         n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977,
         n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985,
         n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993,
         n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001,
         n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009,
         n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017,
         n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025,
         n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033,
         n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041,
         n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049,
         n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
         n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065,
         n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073,
         n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081,
         n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
         n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097,
         n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
         n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113,
         n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121,
         n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
         n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137,
         n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145,
         n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153,
         n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
         n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169,
         n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
         n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185,
         n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193,
         n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
         n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209,
         n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217,
         n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225,
         n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233,
         n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241,
         n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249,
         n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257,
         n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265,
         n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273,
         n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281,
         n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289,
         n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297,
         n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305,
         n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313,
         n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
         n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329,
         n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337,
         n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345,
         n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353,
         n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361,
         n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369,
         n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
         n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385,
         n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
         n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401,
         n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409,
         n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417,
         n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425,
         n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433,
         n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441,
         n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449,
         n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457,
         n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465,
         n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473,
         n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481,
         n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489,
         n47490, n47491, n47492;

  XOR U1 ( .A(n27423), .B(n27905), .Z(n27427) );
  XOR U2 ( .A(n27438), .B(n27902), .Z(n27442) );
  XOR U3 ( .A(n26954), .B(n27412), .Z(n26958) );
  XOR U4 ( .A(n24913), .B(n25397), .Z(n24917) );
  XOR U5 ( .A(n26472), .B(n26912), .Z(n26476) );
  XOR U6 ( .A(n25976), .B(n26410), .Z(n25980) );
  XNOR U7 ( .A(n25982), .B(n25471), .Z(n25473) );
  XOR U8 ( .A(n22777), .B(n23284), .Z(n22781) );
  XOR U9 ( .A(n25483), .B(n25899), .Z(n25487) );
  XOR U10 ( .A(n23916), .B(n24338), .Z(n23920) );
  XOR U11 ( .A(n24456), .B(n24861), .Z(n24460) );
  XOR U12 ( .A(n21114), .B(n21638), .Z(n21118) );
  XOR U13 ( .A(n23936), .B(n24334), .Z(n23940) );
  XOR U14 ( .A(n22872), .B(n23264), .Z(n22876) );
  XOR U15 ( .A(n21764), .B(n22174), .Z(n21768) );
  XOR U16 ( .A(n20607), .B(n21066), .Z(n20611) );
  XOR U17 ( .A(n20642), .B(n21059), .Z(n20646) );
  XOR U18 ( .A(n22353), .B(n22715), .Z(n22357) );
  XOR U19 ( .A(n21814), .B(n22164), .Z(n21818) );
  XOR U20 ( .A(n21264), .B(n21608), .Z(n21268) );
  XOR U21 ( .A(n20717), .B(n21043), .Z(n20721) );
  XOR U22 ( .A(n19592), .B(n19900), .Z(n19596) );
  XNOR U23 ( .A(n27912), .B(n27426), .Z(n27428) );
  XOR U24 ( .A(n25946), .B(n26416), .Z(n25950) );
  XOR U25 ( .A(n27443), .B(n27901), .Z(n27447) );
  XOR U26 ( .A(n26437), .B(n26921), .Z(n26441) );
  XNOR U27 ( .A(n26965), .B(n26465), .Z(n26467) );
  XOR U28 ( .A(n24943), .B(n25391), .Z(n24947) );
  XOR U29 ( .A(n29359), .B(n29793), .Z(n29363) );
  XOR U30 ( .A(n26477), .B(n26911), .Z(n26481) );
  XOR U31 ( .A(n23856), .B(n24350), .Z(n23860) );
  XOR U32 ( .A(n25473), .B(n25901), .Z(n25477) );
  XOR U33 ( .A(n25453), .B(n25906), .Z(n25457) );
  XNOR U34 ( .A(n25479), .B(n24961), .Z(n24963) );
  XOR U35 ( .A(n30733), .B(n31149), .Z(n30737) );
  XOR U36 ( .A(n22782), .B(n23283), .Z(n22786) );
  XOR U37 ( .A(n22807), .B(n23278), .Z(n22811) );
  XOR U38 ( .A(n25488), .B(n25898), .Z(n25492) );
  XOR U39 ( .A(n23921), .B(n24337), .Z(n23925) );
  XOR U40 ( .A(n23876), .B(n24346), .Z(n23880) );
  XOR U41 ( .A(n23360), .B(n23812), .Z(n23364) );
  XNOR U42 ( .A(n24984), .B(n24459), .Z(n24461) );
  XOR U43 ( .A(n32053), .B(n32451), .Z(n32057) );
  XOR U44 ( .A(n22288), .B(n22729), .Z(n22292) );
  XOR U45 ( .A(n21099), .B(n21641), .Z(n21103) );
  XOR U46 ( .A(n21144), .B(n21632), .Z(n21148) );
  XOR U47 ( .A(n23410), .B(n23802), .Z(n23414) );
  XOR U48 ( .A(n22847), .B(n23270), .Z(n22851) );
  XOR U49 ( .A(n19975), .B(n20511), .Z(n19979) );
  XOR U50 ( .A(n19955), .B(n20515), .Z(n19959) );
  XNOR U51 ( .A(n23416), .B(n22875), .Z(n22877) );
  XOR U52 ( .A(n24471), .B(n24857), .Z(n24475) );
  XOR U53 ( .A(n33319), .B(n33699), .Z(n33323) );
  XOR U54 ( .A(n21204), .B(n21620), .Z(n21208) );
  XOR U55 ( .A(n20035), .B(n20499), .Z(n20039) );
  XOR U56 ( .A(n20015), .B(n20503), .Z(n20019) );
  XOR U57 ( .A(n22887), .B(n23261), .Z(n22891) );
  XOR U58 ( .A(n21234), .B(n21614), .Z(n21238) );
  XOR U59 ( .A(n34531), .B(n34893), .Z(n34535) );
  XOR U60 ( .A(n21804), .B(n22166), .Z(n21808) );
  XOR U61 ( .A(n20652), .B(n21057), .Z(n20656) );
  XOR U62 ( .A(n35689), .B(n36033), .Z(n35693) );
  XOR U63 ( .A(n20702), .B(n21046), .Z(n20706) );
  XOR U64 ( .A(n21819), .B(n22163), .Z(n21823) );
  XOR U65 ( .A(n20682), .B(n21051), .Z(n20686) );
  XOR U66 ( .A(n36793), .B(n37119), .Z(n36797) );
  XOR U67 ( .A(n19577), .B(n19903), .Z(n19581) );
  XOR U68 ( .A(n20722), .B(n21042), .Z(n20726) );
  XOR U69 ( .A(n37843), .B(n38151), .Z(n37847) );
  XOR U70 ( .A(n19597), .B(n19899), .Z(n19601) );
  XOR U71 ( .A(n38839), .B(n39129), .Z(n38843) );
  XOR U72 ( .A(n39781), .B(n40053), .Z(n39785) );
  XOR U73 ( .A(n40669), .B(n40923), .Z(n40673) );
  XOR U74 ( .A(n41503), .B(n41739), .Z(n41507) );
  XOR U75 ( .A(n42283), .B(n42501), .Z(n42287) );
  XOR U76 ( .A(n43009), .B(n43209), .Z(n43013) );
  XOR U77 ( .A(n43681), .B(n43863), .Z(n43685) );
  XOR U78 ( .A(n44299), .B(n44463), .Z(n44303) );
  XOR U79 ( .A(n44863), .B(n45009), .Z(n44867) );
  XOR U80 ( .A(n45373), .B(n45501), .Z(n45377) );
  XOR U81 ( .A(n45829), .B(n45939), .Z(n45833) );
  XOR U82 ( .A(n46231), .B(n46323), .Z(n46235) );
  XOR U83 ( .A(n46579), .B(n46653), .Z(n46583) );
  XOR U84 ( .A(n46873), .B(n46929), .Z(n46877) );
  XOR U85 ( .A(n47113), .B(n47151), .Z(n47117) );
  XOR U86 ( .A(n27916), .B(n28386), .Z(n27920) );
  XOR U87 ( .A(n26939), .B(n27415), .Z(n26943) );
  XOR U88 ( .A(n25921), .B(n26421), .Z(n25925) );
  XOR U89 ( .A(n25951), .B(n26415), .Z(n25955) );
  XOR U90 ( .A(n27936), .B(n28382), .Z(n27940) );
  XOR U91 ( .A(n26964), .B(n27410), .Z(n26968) );
  XOR U92 ( .A(n26467), .B(n26913), .Z(n26471) );
  XOR U93 ( .A(n25418), .B(n25913), .Z(n25422) );
  XOR U94 ( .A(n24361), .B(n24882), .Z(n24365) );
  XOR U95 ( .A(n24386), .B(n24877), .Z(n24390) );
  XOR U96 ( .A(n24416), .B(n24871), .Z(n24420) );
  XOR U97 ( .A(n29364), .B(n29792), .Z(n29368) );
  XOR U98 ( .A(n26979), .B(n27407), .Z(n26983) );
  XOR U99 ( .A(n25981), .B(n26409), .Z(n25985) );
  XNOR U100 ( .A(n25987), .B(n25476), .Z(n25478) );
  XOR U101 ( .A(n24928), .B(n25394), .Z(n24932) );
  XOR U102 ( .A(n23300), .B(n23824), .Z(n23304) );
  XOR U103 ( .A(n23846), .B(n24352), .Z(n23850) );
  XNOR U104 ( .A(n25997), .B(n25486), .Z(n25488) );
  XOR U105 ( .A(n22228), .B(n22741), .Z(n22232) );
  XOR U106 ( .A(n24431), .B(n24868), .Z(n24435) );
  XOR U107 ( .A(n30738), .B(n31148), .Z(n30742) );
  XNOR U108 ( .A(n26002), .B(n25491), .Z(n25493) );
  XNOR U109 ( .A(n24979), .B(n24454), .Z(n24456) );
  XOR U110 ( .A(n23380), .B(n23808), .Z(n23384) );
  XOR U111 ( .A(n23335), .B(n23817), .Z(n23339) );
  XOR U112 ( .A(n22258), .B(n22735), .Z(n22262) );
  XOR U113 ( .A(n21659), .B(n22195), .Z(n21663) );
  XOR U114 ( .A(n21119), .B(n21637), .Z(n21123) );
  XOR U115 ( .A(n22822), .B(n23275), .Z(n22826) );
  XOR U116 ( .A(n32058), .B(n32450), .Z(n32062) );
  XOR U117 ( .A(n24466), .B(n24858), .Z(n24470) );
  XOR U118 ( .A(n22293), .B(n22728), .Z(n22297) );
  XOR U119 ( .A(n21714), .B(n22184), .Z(n21718) );
  XOR U120 ( .A(n23946), .B(n24332), .Z(n23950) );
  XOR U121 ( .A(n21174), .B(n21626), .Z(n21178) );
  XOR U122 ( .A(n19397), .B(n19939), .Z(n19401) );
  XOR U123 ( .A(n19960), .B(n20514), .Z(n19964) );
  XOR U124 ( .A(n20005), .B(n20505), .Z(n20009) );
  XOR U125 ( .A(n19985), .B(n20509), .Z(n19989) );
  XOR U126 ( .A(n22882), .B(n23262), .Z(n22886) );
  XOR U127 ( .A(n33324), .B(n33698), .Z(n33328) );
  XOR U128 ( .A(n22308), .B(n22725), .Z(n22312) );
  XOR U129 ( .A(n20567), .B(n21074), .Z(n20571) );
  XOR U130 ( .A(n20637), .B(n21060), .Z(n20641) );
  XOR U131 ( .A(n19457), .B(n19927), .Z(n19461) );
  XOR U132 ( .A(n20020), .B(n20502), .Z(n20024) );
  XOR U133 ( .A(n20667), .B(n21054), .Z(n20671) );
  XOR U134 ( .A(n20045), .B(n20497), .Z(n20049) );
  XOR U135 ( .A(n21784), .B(n22170), .Z(n21788) );
  XOR U136 ( .A(n34536), .B(n34892), .Z(n34540) );
  XOR U137 ( .A(n22358), .B(n22714), .Z(n22362) );
  XOR U138 ( .A(n19492), .B(n19920), .Z(n19496) );
  XOR U139 ( .A(n19522), .B(n19914), .Z(n19526) );
  XOR U140 ( .A(n20085), .B(n20489), .Z(n20089) );
  XOR U141 ( .A(n35694), .B(n36032), .Z(n35698) );
  XOR U142 ( .A(n22373), .B(n22711), .Z(n22377) );
  XOR U143 ( .A(n21269), .B(n21607), .Z(n21273) );
  XOR U144 ( .A(n19552), .B(n19908), .Z(n19556) );
  XOR U145 ( .A(n20115), .B(n20483), .Z(n20119) );
  XOR U146 ( .A(n20145), .B(n20477), .Z(n20149) );
  XOR U147 ( .A(n36798), .B(n37118), .Z(n36802) );
  XNOR U148 ( .A(n21290), .B(n20725), .Z(n20727) );
  XOR U149 ( .A(n19582), .B(n19902), .Z(n19586) );
  XOR U150 ( .A(n37848), .B(n38150), .Z(n37852) );
  XOR U151 ( .A(n19602), .B(n19898), .Z(n19606) );
  XOR U152 ( .A(n38844), .B(n39128), .Z(n38848) );
  XOR U153 ( .A(n39786), .B(n40052), .Z(n39790) );
  XOR U154 ( .A(n40674), .B(n40922), .Z(n40678) );
  XOR U155 ( .A(n5035), .B(n5712), .Z(n5039) );
  XOR U156 ( .A(n41508), .B(n41738), .Z(n41512) );
  XOR U157 ( .A(n42288), .B(n42500), .Z(n42292) );
  XOR U158 ( .A(n43014), .B(n43208), .Z(n43018) );
  XOR U159 ( .A(n10917), .B(n11112), .Z(n10921) );
  XOR U160 ( .A(n43686), .B(n43862), .Z(n43690) );
  XOR U161 ( .A(n9603), .B(n9774), .Z(n9607) );
  XOR U162 ( .A(n44304), .B(n44462), .Z(n44308) );
  XOR U163 ( .A(n44868), .B(n45008), .Z(n44872) );
  XOR U164 ( .A(n8270), .B(n8411), .Z(n8274) );
  XOR U165 ( .A(n45378), .B(n45500), .Z(n45382) );
  XOR U166 ( .A(n6903), .B(n7026), .Z(n6907) );
  XOR U167 ( .A(n45834), .B(n45938), .Z(n45838) );
  XOR U168 ( .A(n46236), .B(n46322), .Z(n46240) );
  XOR U169 ( .A(n46584), .B(n46652), .Z(n46588) );
  XOR U170 ( .A(n47161), .B(n47216), .Z(n47165) );
  XOR U171 ( .A(n46878), .B(n46928), .Z(n46882) );
  XOR U172 ( .A(n47123), .B(n47149), .Z(n47127) );
  XOR U173 ( .A(n27428), .B(n27904), .Z(n27432) );
  XOR U174 ( .A(n27926), .B(n28384), .Z(n27930) );
  XOR U175 ( .A(n26457), .B(n26916), .Z(n26461) );
  XNOR U176 ( .A(n27932), .B(n27446), .Z(n27448) );
  XOR U177 ( .A(n29803), .B(n30255), .Z(n29807) );
  XOR U178 ( .A(n28879), .B(n29331), .Z(n28883) );
  XOR U179 ( .A(n25433), .B(n25910), .Z(n25437) );
  XOR U180 ( .A(n25931), .B(n26419), .Z(n25935) );
  XNOR U181 ( .A(n26970), .B(n26470), .Z(n26472) );
  XOR U182 ( .A(n28418), .B(n28858), .Z(n28422) );
  XOR U183 ( .A(n27458), .B(n27898), .Z(n27462) );
  XNOR U184 ( .A(n26975), .B(n26475), .Z(n26477) );
  XOR U185 ( .A(n24366), .B(n24881), .Z(n24370) );
  XOR U186 ( .A(n30718), .B(n31152), .Z(n30722) );
  XOR U187 ( .A(n29818), .B(n30252), .Z(n29822) );
  XOR U188 ( .A(n24923), .B(n25395), .Z(n24927) );
  XOR U189 ( .A(n24903), .B(n25399), .Z(n24907) );
  XOR U190 ( .A(n23320), .B(n23820), .Z(n23324) );
  XOR U191 ( .A(n22752), .B(n23289), .Z(n22756) );
  XOR U192 ( .A(n23886), .B(n24344), .Z(n23890) );
  XOR U193 ( .A(n29369), .B(n29791), .Z(n29373) );
  XOR U194 ( .A(n28433), .B(n28855), .Z(n28437) );
  XOR U195 ( .A(n27473), .B(n27895), .Z(n27477) );
  XOR U196 ( .A(n26487), .B(n26909), .Z(n26491) );
  XOR U197 ( .A(n24426), .B(n24869), .Z(n24430) );
  XOR U198 ( .A(n32461), .B(n32877), .Z(n32465) );
  XOR U199 ( .A(n31609), .B(n32025), .Z(n31613) );
  XOR U200 ( .A(n24938), .B(n25392), .Z(n24942) );
  XOR U201 ( .A(n24963), .B(n25386), .Z(n24967) );
  XOR U202 ( .A(n21674), .B(n22192), .Z(n21678) );
  XOR U203 ( .A(n22767), .B(n23286), .Z(n22771) );
  XOR U204 ( .A(n21654), .B(n22196), .Z(n21658) );
  XOR U205 ( .A(n31184), .B(n31588), .Z(n31188) );
  XOR U206 ( .A(n30296), .B(n30700), .Z(n30300) );
  XOR U207 ( .A(n29384), .B(n29788), .Z(n29388) );
  XOR U208 ( .A(n28448), .B(n28852), .Z(n28452) );
  XOR U209 ( .A(n27488), .B(n27892), .Z(n27492) );
  XOR U210 ( .A(n26502), .B(n26906), .Z(n26506) );
  XOR U211 ( .A(n25493), .B(n25897), .Z(n25497) );
  XOR U212 ( .A(n23926), .B(n24336), .Z(n23930) );
  XOR U213 ( .A(n22837), .B(n23272), .Z(n22841) );
  XOR U214 ( .A(n22238), .B(n22739), .Z(n22242) );
  XOR U215 ( .A(n23365), .B(n23811), .Z(n23369) );
  XOR U216 ( .A(n22263), .B(n22734), .Z(n22267) );
  XOR U217 ( .A(n33304), .B(n33702), .Z(n33308) );
  XOR U218 ( .A(n32476), .B(n32874), .Z(n32480) );
  XOR U219 ( .A(n22797), .B(n23280), .Z(n22801) );
  XNOR U220 ( .A(n24995), .B(n24469), .Z(n24471) );
  XOR U221 ( .A(n21104), .B(n21640), .Z(n21108) );
  XOR U222 ( .A(n32063), .B(n32449), .Z(n32067) );
  XOR U223 ( .A(n31199), .B(n31585), .Z(n31203) );
  XOR U224 ( .A(n30311), .B(n30697), .Z(n30315) );
  XOR U225 ( .A(n29399), .B(n29785), .Z(n29403) );
  XOR U226 ( .A(n28463), .B(n28849), .Z(n28467) );
  XOR U227 ( .A(n27503), .B(n27889), .Z(n27507) );
  XOR U228 ( .A(n26517), .B(n26903), .Z(n26521) );
  XOR U229 ( .A(n25508), .B(n25894), .Z(n25512) );
  XOR U230 ( .A(n21129), .B(n21635), .Z(n21133) );
  XOR U231 ( .A(n19377), .B(n19943), .Z(n19381) );
  XOR U232 ( .A(n22278), .B(n22731), .Z(n22282) );
  XOR U233 ( .A(n20582), .B(n21071), .Z(n20586) );
  XOR U234 ( .A(n22877), .B(n23263), .Z(n22881) );
  XOR U235 ( .A(n34516), .B(n34896), .Z(n34520) );
  XOR U236 ( .A(n33724), .B(n34104), .Z(n33728) );
  XOR U237 ( .A(n23405), .B(n23803), .Z(n23409) );
  XOR U238 ( .A(n21744), .B(n22178), .Z(n21748) );
  XOR U239 ( .A(n21699), .B(n22187), .Z(n21703) );
  XOR U240 ( .A(n19402), .B(n19938), .Z(n19406) );
  XOR U241 ( .A(n21159), .B(n21629), .Z(n21163) );
  XOR U242 ( .A(n21769), .B(n22173), .Z(n21773) );
  XOR U243 ( .A(n20612), .B(n21065), .Z(n20616) );
  XOR U244 ( .A(n19970), .B(n20512), .Z(n19974) );
  XOR U245 ( .A(n33329), .B(n33697), .Z(n33333) );
  XOR U246 ( .A(n32501), .B(n32869), .Z(n32505) );
  XOR U247 ( .A(n31649), .B(n32017), .Z(n31653) );
  XOR U248 ( .A(n30773), .B(n31141), .Z(n30777) );
  XOR U249 ( .A(n29873), .B(n30241), .Z(n29877) );
  XOR U250 ( .A(n28949), .B(n29317), .Z(n28953) );
  XOR U251 ( .A(n28001), .B(n28369), .Z(n28005) );
  XOR U252 ( .A(n27029), .B(n27397), .Z(n27033) );
  XOR U253 ( .A(n26031), .B(n26399), .Z(n26035) );
  XOR U254 ( .A(n25009), .B(n25377), .Z(n25013) );
  XOR U255 ( .A(n23961), .B(n24329), .Z(n23965) );
  XOR U256 ( .A(n21799), .B(n22167), .Z(n21803) );
  XOR U257 ( .A(n19437), .B(n19931), .Z(n19441) );
  XOR U258 ( .A(n22892), .B(n23260), .Z(n22896) );
  XOR U259 ( .A(n20065), .B(n20493), .Z(n20069) );
  XOR U260 ( .A(n36043), .B(n36405), .Z(n36047) );
  XOR U261 ( .A(n35299), .B(n35661), .Z(n35303) );
  XOR U262 ( .A(n21194), .B(n21622), .Z(n21198) );
  XOR U263 ( .A(n20000), .B(n20506), .Z(n20004) );
  XOR U264 ( .A(n21219), .B(n21617), .Z(n21223) );
  XOR U265 ( .A(n20095), .B(n20487), .Z(n20099) );
  XOR U266 ( .A(n20050), .B(n20496), .Z(n20054) );
  XOR U267 ( .A(n20030), .B(n20500), .Z(n20034) );
  XOR U268 ( .A(n34928), .B(n35278), .Z(n34932) );
  XOR U269 ( .A(n34148), .B(n34498), .Z(n34152) );
  XOR U270 ( .A(n33344), .B(n33694), .Z(n33348) );
  XOR U271 ( .A(n32516), .B(n32866), .Z(n32520) );
  XOR U272 ( .A(n31664), .B(n32014), .Z(n31668) );
  XOR U273 ( .A(n30788), .B(n31138), .Z(n30792) );
  XOR U274 ( .A(n29888), .B(n30238), .Z(n29892) );
  XOR U275 ( .A(n28964), .B(n29314), .Z(n28968) );
  XOR U276 ( .A(n28016), .B(n28366), .Z(n28020) );
  XOR U277 ( .A(n27044), .B(n27394), .Z(n27048) );
  XOR U278 ( .A(n26046), .B(n26396), .Z(n26050) );
  XOR U279 ( .A(n25024), .B(n25374), .Z(n25028) );
  XOR U280 ( .A(n23976), .B(n24326), .Z(n23980) );
  XOR U281 ( .A(n22907), .B(n23257), .Z(n22911) );
  XOR U282 ( .A(n21249), .B(n21611), .Z(n21253) );
  XOR U283 ( .A(n18179), .B(n18747), .Z(n18183) );
  XOR U284 ( .A(n20125), .B(n20481), .Z(n20129) );
  XOR U285 ( .A(n36778), .B(n37122), .Z(n36782) );
  XOR U286 ( .A(n36058), .B(n36402), .Z(n36062) );
  XOR U287 ( .A(n19502), .B(n19918), .Z(n19506) );
  XOR U288 ( .A(n20707), .B(n21045), .Z(n20711) );
  XOR U289 ( .A(n35699), .B(n36031), .Z(n35703) );
  XOR U290 ( .A(n34943), .B(n35275), .Z(n34947) );
  XOR U291 ( .A(n34163), .B(n34495), .Z(n34167) );
  XOR U292 ( .A(n33359), .B(n33691), .Z(n33363) );
  XOR U293 ( .A(n32531), .B(n32863), .Z(n32535) );
  XOR U294 ( .A(n31679), .B(n32011), .Z(n31683) );
  XOR U295 ( .A(n30803), .B(n31135), .Z(n30807) );
  XOR U296 ( .A(n29903), .B(n30235), .Z(n29907) );
  XOR U297 ( .A(n28979), .B(n29311), .Z(n28983) );
  XOR U298 ( .A(n28031), .B(n28363), .Z(n28035) );
  XOR U299 ( .A(n27059), .B(n27391), .Z(n27063) );
  XOR U300 ( .A(n26061), .B(n26393), .Z(n26065) );
  XOR U301 ( .A(n25039), .B(n25371), .Z(n25043) );
  XOR U302 ( .A(n23991), .B(n24323), .Z(n23995) );
  XOR U303 ( .A(n22922), .B(n23254), .Z(n22926) );
  XOR U304 ( .A(n21829), .B(n22161), .Z(n21833) );
  XOR U305 ( .A(n19532), .B(n19912), .Z(n19536) );
  XOR U306 ( .A(n16370), .B(n16871), .Z(n16374) );
  XOR U307 ( .A(n38161), .B(n38487), .Z(n38165) );
  XOR U308 ( .A(n37489), .B(n37815), .Z(n37493) );
  XOR U309 ( .A(n19562), .B(n19906), .Z(n19566) );
  XOR U310 ( .A(n37154), .B(n37468), .Z(n37158) );
  XOR U311 ( .A(n36446), .B(n36760), .Z(n36450) );
  XOR U312 ( .A(n35714), .B(n36028), .Z(n35718) );
  XOR U313 ( .A(n34958), .B(n35272), .Z(n34962) );
  XOR U314 ( .A(n34178), .B(n34492), .Z(n34182) );
  XOR U315 ( .A(n33374), .B(n33688), .Z(n33378) );
  XOR U316 ( .A(n32546), .B(n32860), .Z(n32550) );
  XOR U317 ( .A(n31694), .B(n32008), .Z(n31698) );
  XOR U318 ( .A(n30818), .B(n31132), .Z(n30822) );
  XOR U319 ( .A(n29918), .B(n30232), .Z(n29922) );
  XOR U320 ( .A(n28994), .B(n29308), .Z(n28998) );
  XOR U321 ( .A(n28046), .B(n28360), .Z(n28050) );
  XOR U322 ( .A(n27074), .B(n27388), .Z(n27078) );
  XOR U323 ( .A(n26076), .B(n26390), .Z(n26080) );
  XOR U324 ( .A(n25054), .B(n25368), .Z(n25058) );
  XOR U325 ( .A(n24006), .B(n24320), .Z(n24010) );
  XOR U326 ( .A(n22937), .B(n23251), .Z(n22941) );
  XOR U327 ( .A(n21844), .B(n22158), .Z(n21848) );
  XOR U328 ( .A(n20727), .B(n21041), .Z(n20731) );
  XOR U329 ( .A(n19587), .B(n19901), .Z(n19591) );
  XOR U330 ( .A(n38824), .B(n39132), .Z(n38828) );
  XOR U331 ( .A(n38176), .B(n38484), .Z(n38180) );
  XNOR U332 ( .A(n20176), .B(n19600), .Z(n19602) );
  XOR U333 ( .A(n18329), .B(n18687), .Z(n18333) );
  XOR U334 ( .A(n37853), .B(n38149), .Z(n37857) );
  XOR U335 ( .A(n37169), .B(n37465), .Z(n37173) );
  XOR U336 ( .A(n36461), .B(n36757), .Z(n36465) );
  XOR U337 ( .A(n35729), .B(n36025), .Z(n35733) );
  XOR U338 ( .A(n34973), .B(n35269), .Z(n34977) );
  XOR U339 ( .A(n34193), .B(n34489), .Z(n34197) );
  XOR U340 ( .A(n33389), .B(n33685), .Z(n33393) );
  XOR U341 ( .A(n32561), .B(n32857), .Z(n32565) );
  XOR U342 ( .A(n31709), .B(n32005), .Z(n31713) );
  XOR U343 ( .A(n30833), .B(n31129), .Z(n30837) );
  XOR U344 ( .A(n29933), .B(n30229), .Z(n29937) );
  XOR U345 ( .A(n29009), .B(n29305), .Z(n29013) );
  XOR U346 ( .A(n28061), .B(n28357), .Z(n28065) );
  XOR U347 ( .A(n27089), .B(n27385), .Z(n27093) );
  XOR U348 ( .A(n26091), .B(n26387), .Z(n26095) );
  XOR U349 ( .A(n25069), .B(n25365), .Z(n25073) );
  XOR U350 ( .A(n24021), .B(n24317), .Z(n24025) );
  XOR U351 ( .A(n22952), .B(n23248), .Z(n22956) );
  XOR U352 ( .A(n21859), .B(n22155), .Z(n21863) );
  XOR U353 ( .A(n20742), .B(n21038), .Z(n20746) );
  XNOR U354 ( .A(n20181), .B(n19605), .Z(n19607) );
  XOR U355 ( .A(n11912), .B(n12487), .Z(n11916) );
  XOR U356 ( .A(n40063), .B(n40353), .Z(n40067) );
  XOR U357 ( .A(n39463), .B(n39753), .Z(n39467) );
  XOR U358 ( .A(n10587), .B(n11178), .Z(n10591) );
  XOR U359 ( .A(n18344), .B(n18681), .Z(n18348) );
  XOR U360 ( .A(n9213), .B(n9852), .Z(n9217) );
  XOR U361 ( .A(n39164), .B(n39442), .Z(n39168) );
  XOR U362 ( .A(n38528), .B(n38806), .Z(n38532) );
  XOR U363 ( .A(n37868), .B(n38146), .Z(n37872) );
  XOR U364 ( .A(n37184), .B(n37462), .Z(n37188) );
  XOR U365 ( .A(n36476), .B(n36754), .Z(n36480) );
  XOR U366 ( .A(n35744), .B(n36022), .Z(n35748) );
  XOR U367 ( .A(n34988), .B(n35266), .Z(n34992) );
  XOR U368 ( .A(n34208), .B(n34486), .Z(n34212) );
  XOR U369 ( .A(n33404), .B(n33682), .Z(n33408) );
  XOR U370 ( .A(n32576), .B(n32854), .Z(n32580) );
  XOR U371 ( .A(n31724), .B(n32002), .Z(n31728) );
  XOR U372 ( .A(n30848), .B(n31126), .Z(n30852) );
  XOR U373 ( .A(n29948), .B(n30226), .Z(n29952) );
  XOR U374 ( .A(n29024), .B(n29302), .Z(n29028) );
  XOR U375 ( .A(n28076), .B(n28354), .Z(n28080) );
  XOR U376 ( .A(n27104), .B(n27382), .Z(n27108) );
  XOR U377 ( .A(n26106), .B(n26384), .Z(n26110) );
  XOR U378 ( .A(n25084), .B(n25362), .Z(n25088) );
  XOR U379 ( .A(n24036), .B(n24314), .Z(n24040) );
  XOR U380 ( .A(n22967), .B(n23245), .Z(n22971) );
  XOR U381 ( .A(n21874), .B(n22152), .Z(n21878) );
  XOR U382 ( .A(n20757), .B(n21035), .Z(n20761) );
  XOR U383 ( .A(n19617), .B(n19895), .Z(n19621) );
  XOR U384 ( .A(n16550), .B(n16835), .Z(n16554) );
  XOR U385 ( .A(n40654), .B(n40926), .Z(n40658) );
  XOR U386 ( .A(n40078), .B(n40350), .Z(n40082) );
  XOR U387 ( .A(n8562), .B(n9171), .Z(n8566) );
  XOR U388 ( .A(n7152), .B(n7809), .Z(n7156) );
  XOR U389 ( .A(n9978), .B(n10503), .Z(n9982) );
  XOR U390 ( .A(n39791), .B(n40051), .Z(n39795) );
  XOR U391 ( .A(n39179), .B(n39439), .Z(n39183) );
  XOR U392 ( .A(n38543), .B(n38803), .Z(n38547) );
  XOR U393 ( .A(n37883), .B(n38143), .Z(n37887) );
  XOR U394 ( .A(n37199), .B(n37459), .Z(n37203) );
  XOR U395 ( .A(n36491), .B(n36751), .Z(n36495) );
  XOR U396 ( .A(n35759), .B(n36019), .Z(n35763) );
  XOR U397 ( .A(n35003), .B(n35263), .Z(n35007) );
  XOR U398 ( .A(n34223), .B(n34483), .Z(n34227) );
  XOR U399 ( .A(n33419), .B(n33679), .Z(n33423) );
  XOR U400 ( .A(n32591), .B(n32851), .Z(n32595) );
  XOR U401 ( .A(n31739), .B(n31999), .Z(n31743) );
  XOR U402 ( .A(n30863), .B(n31123), .Z(n30867) );
  XOR U403 ( .A(n29963), .B(n30223), .Z(n29967) );
  XOR U404 ( .A(n29039), .B(n29299), .Z(n29043) );
  XOR U405 ( .A(n28091), .B(n28351), .Z(n28095) );
  XOR U406 ( .A(n27119), .B(n27379), .Z(n27123) );
  XOR U407 ( .A(n26121), .B(n26381), .Z(n26125) );
  XOR U408 ( .A(n25099), .B(n25359), .Z(n25103) );
  XOR U409 ( .A(n24051), .B(n24311), .Z(n24055) );
  XOR U410 ( .A(n22982), .B(n23242), .Z(n22986) );
  XOR U411 ( .A(n21889), .B(n22149), .Z(n21893) );
  XOR U412 ( .A(n20772), .B(n21032), .Z(n20776) );
  XOR U413 ( .A(n19632), .B(n19892), .Z(n19636) );
  XOR U414 ( .A(n41749), .B(n42003), .Z(n41753) );
  XOR U415 ( .A(n41221), .B(n41475), .Z(n41225) );
  XOR U416 ( .A(n10008), .B(n10497), .Z(n10012) );
  XOR U417 ( .A(n16580), .B(n16829), .Z(n16584) );
  XOR U418 ( .A(n10038), .B(n10491), .Z(n10042) );
  XOR U419 ( .A(n40958), .B(n41200), .Z(n40962) );
  XOR U420 ( .A(n40394), .B(n40636), .Z(n40398) );
  XOR U421 ( .A(n39806), .B(n40048), .Z(n39810) );
  XOR U422 ( .A(n39194), .B(n39436), .Z(n39198) );
  XOR U423 ( .A(n38558), .B(n38800), .Z(n38562) );
  XOR U424 ( .A(n37898), .B(n38140), .Z(n37902) );
  XOR U425 ( .A(n37214), .B(n37456), .Z(n37218) );
  XOR U426 ( .A(n36506), .B(n36748), .Z(n36510) );
  XOR U427 ( .A(n35774), .B(n36016), .Z(n35778) );
  XOR U428 ( .A(n35018), .B(n35260), .Z(n35022) );
  XOR U429 ( .A(n34238), .B(n34480), .Z(n34242) );
  XOR U430 ( .A(n33434), .B(n33676), .Z(n33438) );
  XOR U431 ( .A(n32606), .B(n32848), .Z(n32610) );
  XOR U432 ( .A(n31754), .B(n31996), .Z(n31758) );
  XOR U433 ( .A(n30878), .B(n31120), .Z(n30882) );
  XOR U434 ( .A(n29978), .B(n30220), .Z(n29982) );
  XOR U435 ( .A(n29054), .B(n29296), .Z(n29058) );
  XOR U436 ( .A(n28106), .B(n28348), .Z(n28110) );
  XOR U437 ( .A(n27134), .B(n27376), .Z(n27138) );
  XOR U438 ( .A(n26136), .B(n26378), .Z(n26140) );
  XOR U439 ( .A(n25114), .B(n25356), .Z(n25118) );
  XOR U440 ( .A(n24066), .B(n24308), .Z(n24070) );
  XOR U441 ( .A(n22997), .B(n23239), .Z(n23001) );
  XOR U442 ( .A(n21904), .B(n22146), .Z(n21908) );
  XOR U443 ( .A(n20787), .B(n21029), .Z(n20791) );
  XOR U444 ( .A(n19647), .B(n19889), .Z(n19651) );
  XOR U445 ( .A(n15359), .B(n15602), .Z(n15363) );
  XOR U446 ( .A(n42268), .B(n42504), .Z(n42272) );
  XOR U447 ( .A(n41764), .B(n42000), .Z(n41768) );
  XOR U448 ( .A(n10068), .B(n10485), .Z(n10072) );
  XOR U449 ( .A(n3595), .B(n4282), .Z(n3599) );
  XOR U450 ( .A(n14747), .B(n14978), .Z(n14751) );
  XOR U451 ( .A(n10098), .B(n10479), .Z(n10102) );
  XOR U452 ( .A(n41513), .B(n41737), .Z(n41517) );
  XOR U453 ( .A(n40973), .B(n41197), .Z(n40977) );
  XOR U454 ( .A(n40409), .B(n40633), .Z(n40413) );
  XOR U455 ( .A(n39821), .B(n40045), .Z(n39825) );
  XOR U456 ( .A(n39209), .B(n39433), .Z(n39213) );
  XOR U457 ( .A(n38573), .B(n38797), .Z(n38577) );
  XOR U458 ( .A(n37913), .B(n38137), .Z(n37917) );
  XOR U459 ( .A(n37229), .B(n37453), .Z(n37233) );
  XOR U460 ( .A(n36521), .B(n36745), .Z(n36525) );
  XOR U461 ( .A(n35789), .B(n36013), .Z(n35793) );
  XOR U462 ( .A(n35033), .B(n35257), .Z(n35037) );
  XOR U463 ( .A(n34253), .B(n34477), .Z(n34257) );
  XOR U464 ( .A(n33449), .B(n33673), .Z(n33453) );
  XOR U465 ( .A(n32621), .B(n32845), .Z(n32625) );
  XOR U466 ( .A(n31769), .B(n31993), .Z(n31773) );
  XOR U467 ( .A(n30893), .B(n31117), .Z(n30897) );
  XOR U468 ( .A(n29993), .B(n30217), .Z(n29997) );
  XOR U469 ( .A(n29069), .B(n29293), .Z(n29073) );
  XOR U470 ( .A(n28121), .B(n28345), .Z(n28125) );
  XOR U471 ( .A(n27149), .B(n27373), .Z(n27153) );
  XOR U472 ( .A(n26151), .B(n26375), .Z(n26155) );
  XOR U473 ( .A(n25129), .B(n25353), .Z(n25133) );
  XOR U474 ( .A(n24081), .B(n24305), .Z(n24085) );
  XOR U475 ( .A(n23012), .B(n23236), .Z(n23016) );
  XOR U476 ( .A(n21919), .B(n22143), .Z(n21923) );
  XOR U477 ( .A(n20802), .B(n21026), .Z(n20806) );
  XOR U478 ( .A(n19662), .B(n19886), .Z(n19666) );
  XOR U479 ( .A(n43219), .B(n43437), .Z(n43223) );
  XOR U480 ( .A(n42763), .B(n42981), .Z(n42767) );
  XOR U481 ( .A(n14129), .B(n14348), .Z(n14133) );
  XOR U482 ( .A(n10128), .B(n10473), .Z(n10132) );
  XOR U483 ( .A(n12860), .B(n13073), .Z(n12864) );
  XOR U484 ( .A(n10158), .B(n10467), .Z(n10162) );
  XOR U485 ( .A(n42536), .B(n42742), .Z(n42540) );
  XOR U486 ( .A(n42044), .B(n42250), .Z(n42048) );
  XOR U487 ( .A(n41528), .B(n41734), .Z(n41532) );
  XOR U488 ( .A(n40988), .B(n41194), .Z(n40992) );
  XOR U489 ( .A(n40424), .B(n40630), .Z(n40428) );
  XOR U490 ( .A(n39836), .B(n40042), .Z(n39840) );
  XOR U491 ( .A(n39224), .B(n39430), .Z(n39228) );
  XOR U492 ( .A(n38588), .B(n38794), .Z(n38592) );
  XOR U493 ( .A(n37928), .B(n38134), .Z(n37932) );
  XOR U494 ( .A(n37244), .B(n37450), .Z(n37248) );
  XOR U495 ( .A(n36536), .B(n36742), .Z(n36540) );
  XOR U496 ( .A(n35804), .B(n36010), .Z(n35808) );
  XOR U497 ( .A(n35048), .B(n35254), .Z(n35052) );
  XOR U498 ( .A(n34268), .B(n34474), .Z(n34272) );
  XOR U499 ( .A(n33464), .B(n33670), .Z(n33468) );
  XOR U500 ( .A(n32636), .B(n32842), .Z(n32640) );
  XOR U501 ( .A(n31784), .B(n31990), .Z(n31788) );
  XOR U502 ( .A(n30908), .B(n31114), .Z(n30912) );
  XOR U503 ( .A(n30008), .B(n30214), .Z(n30012) );
  XOR U504 ( .A(n29084), .B(n29290), .Z(n29088) );
  XOR U505 ( .A(n28136), .B(n28342), .Z(n28140) );
  XOR U506 ( .A(n27164), .B(n27370), .Z(n27168) );
  XOR U507 ( .A(n26166), .B(n26372), .Z(n26170) );
  XOR U508 ( .A(n25144), .B(n25350), .Z(n25148) );
  XOR U509 ( .A(n24096), .B(n24302), .Z(n24100) );
  XOR U510 ( .A(n23027), .B(n23233), .Z(n23031) );
  XOR U511 ( .A(n21934), .B(n22140), .Z(n21938) );
  XOR U512 ( .A(n20817), .B(n21023), .Z(n20821) );
  XOR U513 ( .A(n19677), .B(n19883), .Z(n19681) );
  XOR U514 ( .A(n43666), .B(n43866), .Z(n43670) );
  XOR U515 ( .A(n43234), .B(n43434), .Z(n43238) );
  XOR U516 ( .A(n10188), .B(n10461), .Z(n10192) );
  XOR U517 ( .A(n10218), .B(n10455), .Z(n10222) );
  XOR U518 ( .A(n43019), .B(n43207), .Z(n43023) );
  XOR U519 ( .A(n42551), .B(n42739), .Z(n42555) );
  XOR U520 ( .A(n42059), .B(n42247), .Z(n42063) );
  XOR U521 ( .A(n41543), .B(n41731), .Z(n41547) );
  XOR U522 ( .A(n41003), .B(n41191), .Z(n41007) );
  XOR U523 ( .A(n40439), .B(n40627), .Z(n40443) );
  XOR U524 ( .A(n39851), .B(n40039), .Z(n39855) );
  XOR U525 ( .A(n39239), .B(n39427), .Z(n39243) );
  XOR U526 ( .A(n38603), .B(n38791), .Z(n38607) );
  XOR U527 ( .A(n37943), .B(n38131), .Z(n37947) );
  XOR U528 ( .A(n37259), .B(n37447), .Z(n37263) );
  XOR U529 ( .A(n36551), .B(n36739), .Z(n36555) );
  XOR U530 ( .A(n35819), .B(n36007), .Z(n35823) );
  XOR U531 ( .A(n35063), .B(n35251), .Z(n35067) );
  XOR U532 ( .A(n34283), .B(n34471), .Z(n34287) );
  XOR U533 ( .A(n33479), .B(n33667), .Z(n33483) );
  XOR U534 ( .A(n32651), .B(n32839), .Z(n32655) );
  XOR U535 ( .A(n31799), .B(n31987), .Z(n31803) );
  XOR U536 ( .A(n30923), .B(n31111), .Z(n30927) );
  XOR U537 ( .A(n30023), .B(n30211), .Z(n30027) );
  XOR U538 ( .A(n29099), .B(n29287), .Z(n29103) );
  XOR U539 ( .A(n28151), .B(n28339), .Z(n28155) );
  XOR U540 ( .A(n27179), .B(n27367), .Z(n27183) );
  XOR U541 ( .A(n26181), .B(n26369), .Z(n26185) );
  XOR U542 ( .A(n25159), .B(n25347), .Z(n25163) );
  XOR U543 ( .A(n24111), .B(n24299), .Z(n24115) );
  XOR U544 ( .A(n23042), .B(n23230), .Z(n23046) );
  XOR U545 ( .A(n21949), .B(n22137), .Z(n21953) );
  XOR U546 ( .A(n20832), .B(n21020), .Z(n20836) );
  XOR U547 ( .A(n19692), .B(n19880), .Z(n19696) );
  XOR U548 ( .A(n44473), .B(n44655), .Z(n44477) );
  XOR U549 ( .A(n44089), .B(n44271), .Z(n44093) );
  XOR U550 ( .A(n10248), .B(n10449), .Z(n10252) );
  XOR U551 ( .A(n10927), .B(n11110), .Z(n10931) );
  XOR U552 ( .A(n43898), .B(n44068), .Z(n43902) );
  XOR U553 ( .A(n43478), .B(n43648), .Z(n43482) );
  XOR U554 ( .A(n43034), .B(n43204), .Z(n43038) );
  XOR U555 ( .A(n42566), .B(n42736), .Z(n42570) );
  XOR U556 ( .A(n42074), .B(n42244), .Z(n42078) );
  XOR U557 ( .A(n41558), .B(n41728), .Z(n41562) );
  XOR U558 ( .A(n41018), .B(n41188), .Z(n41022) );
  XOR U559 ( .A(n40454), .B(n40624), .Z(n40458) );
  XOR U560 ( .A(n39866), .B(n40036), .Z(n39870) );
  XOR U561 ( .A(n39254), .B(n39424), .Z(n39258) );
  XOR U562 ( .A(n38618), .B(n38788), .Z(n38622) );
  XOR U563 ( .A(n37958), .B(n38128), .Z(n37962) );
  XOR U564 ( .A(n37274), .B(n37444), .Z(n37278) );
  XOR U565 ( .A(n36566), .B(n36736), .Z(n36570) );
  XOR U566 ( .A(n35834), .B(n36004), .Z(n35838) );
  XOR U567 ( .A(n35078), .B(n35248), .Z(n35082) );
  XOR U568 ( .A(n34298), .B(n34468), .Z(n34302) );
  XOR U569 ( .A(n33494), .B(n33664), .Z(n33498) );
  XOR U570 ( .A(n32666), .B(n32836), .Z(n32670) );
  XOR U571 ( .A(n31814), .B(n31984), .Z(n31818) );
  XOR U572 ( .A(n30938), .B(n31108), .Z(n30942) );
  XOR U573 ( .A(n30038), .B(n30208), .Z(n30042) );
  XOR U574 ( .A(n29114), .B(n29284), .Z(n29118) );
  XOR U575 ( .A(n28166), .B(n28336), .Z(n28170) );
  XOR U576 ( .A(n27194), .B(n27364), .Z(n27198) );
  XOR U577 ( .A(n26196), .B(n26366), .Z(n26200) );
  XOR U578 ( .A(n25174), .B(n25344), .Z(n25178) );
  XOR U579 ( .A(n24126), .B(n24296), .Z(n24130) );
  XOR U580 ( .A(n23057), .B(n23227), .Z(n23061) );
  XOR U581 ( .A(n21964), .B(n22134), .Z(n21968) );
  XOR U582 ( .A(n20847), .B(n21017), .Z(n20851) );
  XOR U583 ( .A(n19707), .B(n19877), .Z(n19711) );
  XOR U584 ( .A(n44848), .B(n45012), .Z(n44852) );
  XOR U585 ( .A(n44488), .B(n44652), .Z(n44492) );
  XOR U586 ( .A(n10278), .B(n10443), .Z(n10282) );
  XOR U587 ( .A(n11605), .B(n11764), .Z(n11609) );
  XOR U588 ( .A(n44309), .B(n44461), .Z(n44313) );
  XOR U589 ( .A(n43913), .B(n44065), .Z(n43917) );
  XOR U590 ( .A(n43493), .B(n43645), .Z(n43497) );
  XOR U591 ( .A(n43049), .B(n43201), .Z(n43053) );
  XOR U592 ( .A(n42581), .B(n42733), .Z(n42585) );
  XOR U593 ( .A(n42089), .B(n42241), .Z(n42093) );
  XOR U594 ( .A(n41573), .B(n41725), .Z(n41577) );
  XOR U595 ( .A(n41033), .B(n41185), .Z(n41037) );
  XOR U596 ( .A(n40469), .B(n40621), .Z(n40473) );
  XOR U597 ( .A(n39881), .B(n40033), .Z(n39885) );
  XOR U598 ( .A(n39269), .B(n39421), .Z(n39273) );
  XOR U599 ( .A(n38633), .B(n38785), .Z(n38637) );
  XOR U600 ( .A(n37973), .B(n38125), .Z(n37977) );
  XOR U601 ( .A(n37289), .B(n37441), .Z(n37293) );
  XOR U602 ( .A(n36581), .B(n36733), .Z(n36585) );
  XOR U603 ( .A(n35849), .B(n36001), .Z(n35853) );
  XOR U604 ( .A(n35093), .B(n35245), .Z(n35097) );
  XOR U605 ( .A(n34313), .B(n34465), .Z(n34317) );
  XOR U606 ( .A(n33509), .B(n33661), .Z(n33513) );
  XOR U607 ( .A(n32681), .B(n32833), .Z(n32685) );
  XOR U608 ( .A(n31829), .B(n31981), .Z(n31833) );
  XOR U609 ( .A(n30953), .B(n31105), .Z(n30957) );
  XOR U610 ( .A(n30053), .B(n30205), .Z(n30057) );
  XOR U611 ( .A(n29129), .B(n29281), .Z(n29133) );
  XOR U612 ( .A(n28181), .B(n28333), .Z(n28185) );
  XOR U613 ( .A(n27209), .B(n27361), .Z(n27213) );
  XOR U614 ( .A(n26211), .B(n26363), .Z(n26215) );
  XOR U615 ( .A(n25189), .B(n25341), .Z(n25193) );
  XOR U616 ( .A(n24141), .B(n24293), .Z(n24145) );
  XOR U617 ( .A(n23072), .B(n23224), .Z(n23076) );
  XOR U618 ( .A(n21979), .B(n22131), .Z(n21983) );
  XOR U619 ( .A(n20862), .B(n21014), .Z(n20866) );
  XOR U620 ( .A(n19722), .B(n19874), .Z(n19726) );
  XOR U621 ( .A(n45511), .B(n45657), .Z(n45515) );
  XOR U622 ( .A(n45199), .B(n45345), .Z(n45203) );
  XOR U623 ( .A(n8952), .B(n9093), .Z(n8956) );
  XOR U624 ( .A(n45044), .B(n45178), .Z(n45048) );
  XOR U625 ( .A(n44696), .B(n44830), .Z(n44700) );
  XOR U626 ( .A(n44324), .B(n44458), .Z(n44328) );
  XOR U627 ( .A(n43928), .B(n44062), .Z(n43932) );
  XOR U628 ( .A(n43508), .B(n43642), .Z(n43512) );
  XOR U629 ( .A(n43064), .B(n43198), .Z(n43068) );
  XOR U630 ( .A(n42596), .B(n42730), .Z(n42600) );
  XOR U631 ( .A(n42104), .B(n42238), .Z(n42108) );
  XOR U632 ( .A(n41588), .B(n41722), .Z(n41592) );
  XOR U633 ( .A(n41048), .B(n41182), .Z(n41052) );
  XOR U634 ( .A(n40484), .B(n40618), .Z(n40488) );
  XOR U635 ( .A(n39896), .B(n40030), .Z(n39900) );
  XOR U636 ( .A(n39284), .B(n39418), .Z(n39288) );
  XOR U637 ( .A(n38648), .B(n38782), .Z(n38652) );
  XOR U638 ( .A(n37988), .B(n38122), .Z(n37992) );
  XOR U639 ( .A(n37304), .B(n37438), .Z(n37308) );
  XOR U640 ( .A(n36596), .B(n36730), .Z(n36600) );
  XOR U641 ( .A(n35864), .B(n35998), .Z(n35868) );
  XOR U642 ( .A(n35108), .B(n35242), .Z(n35112) );
  XOR U643 ( .A(n34328), .B(n34462), .Z(n34332) );
  XOR U644 ( .A(n33524), .B(n33658), .Z(n33528) );
  XOR U645 ( .A(n32696), .B(n32830), .Z(n32700) );
  XOR U646 ( .A(n31844), .B(n31978), .Z(n31848) );
  XOR U647 ( .A(n30968), .B(n31102), .Z(n30972) );
  XOR U648 ( .A(n30068), .B(n30202), .Z(n30072) );
  XOR U649 ( .A(n29144), .B(n29278), .Z(n29148) );
  XOR U650 ( .A(n28196), .B(n28330), .Z(n28200) );
  XOR U651 ( .A(n27224), .B(n27358), .Z(n27228) );
  XOR U652 ( .A(n26226), .B(n26360), .Z(n26230) );
  XOR U653 ( .A(n25204), .B(n25338), .Z(n25208) );
  XOR U654 ( .A(n24156), .B(n24290), .Z(n24160) );
  XOR U655 ( .A(n23087), .B(n23221), .Z(n23091) );
  XOR U656 ( .A(n21994), .B(n22128), .Z(n21998) );
  XOR U657 ( .A(n20877), .B(n21011), .Z(n20881) );
  XOR U658 ( .A(n19737), .B(n19871), .Z(n19741) );
  XOR U659 ( .A(n45814), .B(n45942), .Z(n45818) );
  XOR U660 ( .A(n45526), .B(n45654), .Z(n45530) );
  XOR U661 ( .A(n8280), .B(n8409), .Z(n8284) );
  XOR U662 ( .A(n45383), .B(n45499), .Z(n45387) );
  XOR U663 ( .A(n45059), .B(n45175), .Z(n45063) );
  XOR U664 ( .A(n44711), .B(n44827), .Z(n44715) );
  XOR U665 ( .A(n44339), .B(n44455), .Z(n44343) );
  XOR U666 ( .A(n43943), .B(n44059), .Z(n43947) );
  XOR U667 ( .A(n43523), .B(n43639), .Z(n43527) );
  XOR U668 ( .A(n43079), .B(n43195), .Z(n43083) );
  XOR U669 ( .A(n42611), .B(n42727), .Z(n42615) );
  XOR U670 ( .A(n42119), .B(n42235), .Z(n42123) );
  XOR U671 ( .A(n41603), .B(n41719), .Z(n41607) );
  XOR U672 ( .A(n41063), .B(n41179), .Z(n41067) );
  XOR U673 ( .A(n40499), .B(n40615), .Z(n40503) );
  XOR U674 ( .A(n39911), .B(n40027), .Z(n39915) );
  XOR U675 ( .A(n39299), .B(n39415), .Z(n39303) );
  XOR U676 ( .A(n38663), .B(n38779), .Z(n38667) );
  XOR U677 ( .A(n38003), .B(n38119), .Z(n38007) );
  XOR U678 ( .A(n37319), .B(n37435), .Z(n37323) );
  XOR U679 ( .A(n36611), .B(n36727), .Z(n36615) );
  XOR U680 ( .A(n35879), .B(n35995), .Z(n35883) );
  XOR U681 ( .A(n35123), .B(n35239), .Z(n35127) );
  XOR U682 ( .A(n34343), .B(n34459), .Z(n34347) );
  XOR U683 ( .A(n33539), .B(n33655), .Z(n33543) );
  XOR U684 ( .A(n32711), .B(n32827), .Z(n32715) );
  XOR U685 ( .A(n31859), .B(n31975), .Z(n31863) );
  XOR U686 ( .A(n30983), .B(n31099), .Z(n30987) );
  XOR U687 ( .A(n30083), .B(n30199), .Z(n30087) );
  XOR U688 ( .A(n29159), .B(n29275), .Z(n29163) );
  XOR U689 ( .A(n28211), .B(n28327), .Z(n28215) );
  XOR U690 ( .A(n27239), .B(n27355), .Z(n27243) );
  XOR U691 ( .A(n26241), .B(n26357), .Z(n26245) );
  XOR U692 ( .A(n25219), .B(n25335), .Z(n25223) );
  XOR U693 ( .A(n24171), .B(n24287), .Z(n24175) );
  XOR U694 ( .A(n23102), .B(n23218), .Z(n23106) );
  XOR U695 ( .A(n22009), .B(n22125), .Z(n22013) );
  XOR U696 ( .A(n20892), .B(n21008), .Z(n20896) );
  XOR U697 ( .A(n19752), .B(n19868), .Z(n19756) );
  XOR U698 ( .A(n6203), .B(n6326), .Z(n6207) );
  XOR U699 ( .A(n46333), .B(n46443), .Z(n46337) );
  XOR U700 ( .A(n46093), .B(n46203), .Z(n46097) );
  XOR U701 ( .A(n6918), .B(n7023), .Z(n6922) );
  XOR U702 ( .A(n45974), .B(n46072), .Z(n45978) );
  XOR U703 ( .A(n45698), .B(n45796), .Z(n45702) );
  XOR U704 ( .A(n45398), .B(n45496), .Z(n45402) );
  XOR U705 ( .A(n45074), .B(n45172), .Z(n45078) );
  XOR U706 ( .A(n44726), .B(n44824), .Z(n44730) );
  XOR U707 ( .A(n44354), .B(n44452), .Z(n44358) );
  XOR U708 ( .A(n43958), .B(n44056), .Z(n43962) );
  XOR U709 ( .A(n43538), .B(n43636), .Z(n43542) );
  XOR U710 ( .A(n43094), .B(n43192), .Z(n43098) );
  XOR U711 ( .A(n42626), .B(n42724), .Z(n42630) );
  XOR U712 ( .A(n42134), .B(n42232), .Z(n42138) );
  XOR U713 ( .A(n41618), .B(n41716), .Z(n41622) );
  XOR U714 ( .A(n41078), .B(n41176), .Z(n41082) );
  XOR U715 ( .A(n40514), .B(n40612), .Z(n40518) );
  XOR U716 ( .A(n39926), .B(n40024), .Z(n39930) );
  XOR U717 ( .A(n39314), .B(n39412), .Z(n39318) );
  XOR U718 ( .A(n38678), .B(n38776), .Z(n38682) );
  XOR U719 ( .A(n38018), .B(n38116), .Z(n38022) );
  XOR U720 ( .A(n37334), .B(n37432), .Z(n37338) );
  XOR U721 ( .A(n36626), .B(n36724), .Z(n36630) );
  XOR U722 ( .A(n35894), .B(n35992), .Z(n35898) );
  XOR U723 ( .A(n35138), .B(n35236), .Z(n35142) );
  XOR U724 ( .A(n34358), .B(n34456), .Z(n34362) );
  XOR U725 ( .A(n33554), .B(n33652), .Z(n33558) );
  XOR U726 ( .A(n32726), .B(n32824), .Z(n32730) );
  XOR U727 ( .A(n31874), .B(n31972), .Z(n31878) );
  XOR U728 ( .A(n30998), .B(n31096), .Z(n31002) );
  XOR U729 ( .A(n30098), .B(n30196), .Z(n30102) );
  XOR U730 ( .A(n29174), .B(n29272), .Z(n29178) );
  XOR U731 ( .A(n28226), .B(n28324), .Z(n28230) );
  XOR U732 ( .A(n27254), .B(n27352), .Z(n27258) );
  XOR U733 ( .A(n26256), .B(n26354), .Z(n26260) );
  XOR U734 ( .A(n25234), .B(n25332), .Z(n25238) );
  XOR U735 ( .A(n24186), .B(n24284), .Z(n24190) );
  XOR U736 ( .A(n23117), .B(n23215), .Z(n23121) );
  XOR U737 ( .A(n22024), .B(n22122), .Z(n22028) );
  XOR U738 ( .A(n20907), .B(n21005), .Z(n20911) );
  XOR U739 ( .A(n19767), .B(n19865), .Z(n19771) );
  XOR U740 ( .A(n5515), .B(n5616), .Z(n5519) );
  XOR U741 ( .A(n46564), .B(n46656), .Z(n46568) );
  XOR U742 ( .A(n46348), .B(n46440), .Z(n46352) );
  XOR U743 ( .A(n46241), .B(n46321), .Z(n46245) );
  XOR U744 ( .A(n45989), .B(n46069), .Z(n45993) );
  XOR U745 ( .A(n45713), .B(n45793), .Z(n45717) );
  XOR U746 ( .A(n45413), .B(n45493), .Z(n45417) );
  XOR U747 ( .A(n45089), .B(n45169), .Z(n45093) );
  XOR U748 ( .A(n44741), .B(n44821), .Z(n44745) );
  XOR U749 ( .A(n44369), .B(n44449), .Z(n44373) );
  XOR U750 ( .A(n43973), .B(n44053), .Z(n43977) );
  XOR U751 ( .A(n43553), .B(n43633), .Z(n43557) );
  XOR U752 ( .A(n43109), .B(n43189), .Z(n43113) );
  XOR U753 ( .A(n42641), .B(n42721), .Z(n42645) );
  XOR U754 ( .A(n42149), .B(n42229), .Z(n42153) );
  XOR U755 ( .A(n41633), .B(n41713), .Z(n41637) );
  XOR U756 ( .A(n41093), .B(n41173), .Z(n41097) );
  XOR U757 ( .A(n40529), .B(n40609), .Z(n40533) );
  XOR U758 ( .A(n39941), .B(n40021), .Z(n39945) );
  XOR U759 ( .A(n39329), .B(n39409), .Z(n39333) );
  XOR U760 ( .A(n38693), .B(n38773), .Z(n38697) );
  XOR U761 ( .A(n38033), .B(n38113), .Z(n38037) );
  XOR U762 ( .A(n37349), .B(n37429), .Z(n37353) );
  XOR U763 ( .A(n36641), .B(n36721), .Z(n36645) );
  XOR U764 ( .A(n35909), .B(n35989), .Z(n35913) );
  XOR U765 ( .A(n35153), .B(n35233), .Z(n35157) );
  XOR U766 ( .A(n34373), .B(n34453), .Z(n34377) );
  XOR U767 ( .A(n33569), .B(n33649), .Z(n33573) );
  XOR U768 ( .A(n32741), .B(n32821), .Z(n32745) );
  XOR U769 ( .A(n31889), .B(n31969), .Z(n31893) );
  XOR U770 ( .A(n31013), .B(n31093), .Z(n31017) );
  XOR U771 ( .A(n30113), .B(n30193), .Z(n30117) );
  XOR U772 ( .A(n29189), .B(n29269), .Z(n29193) );
  XOR U773 ( .A(n28241), .B(n28321), .Z(n28245) );
  XOR U774 ( .A(n27269), .B(n27349), .Z(n27273) );
  XOR U775 ( .A(n26271), .B(n26351), .Z(n26275) );
  XOR U776 ( .A(n25249), .B(n25329), .Z(n25253) );
  XOR U777 ( .A(n24201), .B(n24281), .Z(n24205) );
  XOR U778 ( .A(n23132), .B(n23212), .Z(n23136) );
  XOR U779 ( .A(n22039), .B(n22119), .Z(n22043) );
  XOR U780 ( .A(n20922), .B(n21002), .Z(n20926) );
  XOR U781 ( .A(n19782), .B(n19862), .Z(n19786) );
  XOR U782 ( .A(n46939), .B(n47013), .Z(n46943) );
  XOR U783 ( .A(n46771), .B(n46845), .Z(n46775) );
  XOR U784 ( .A(n4105), .B(n4180), .Z(n4109) );
  XOR U785 ( .A(n46688), .B(n46750), .Z(n46692) );
  XOR U786 ( .A(n46484), .B(n46546), .Z(n46488) );
  XOR U787 ( .A(n46256), .B(n46318), .Z(n46260) );
  XOR U788 ( .A(n46004), .B(n46066), .Z(n46008) );
  XOR U789 ( .A(n45728), .B(n45790), .Z(n45732) );
  XOR U790 ( .A(n45428), .B(n45490), .Z(n45432) );
  XOR U791 ( .A(n45104), .B(n45166), .Z(n45108) );
  XOR U792 ( .A(n44756), .B(n44818), .Z(n44760) );
  XOR U793 ( .A(n44384), .B(n44446), .Z(n44388) );
  XOR U794 ( .A(n43988), .B(n44050), .Z(n43992) );
  XOR U795 ( .A(n43568), .B(n43630), .Z(n43572) );
  XOR U796 ( .A(n43124), .B(n43186), .Z(n43128) );
  XOR U797 ( .A(n42656), .B(n42718), .Z(n42660) );
  XOR U798 ( .A(n42164), .B(n42226), .Z(n42168) );
  XOR U799 ( .A(n41648), .B(n41710), .Z(n41652) );
  XOR U800 ( .A(n41108), .B(n41170), .Z(n41112) );
  XOR U801 ( .A(n40544), .B(n40606), .Z(n40548) );
  XOR U802 ( .A(n39956), .B(n40018), .Z(n39960) );
  XOR U803 ( .A(n39344), .B(n39406), .Z(n39348) );
  XOR U804 ( .A(n38708), .B(n38770), .Z(n38712) );
  XOR U805 ( .A(n38048), .B(n38110), .Z(n38052) );
  XOR U806 ( .A(n37364), .B(n37426), .Z(n37368) );
  XOR U807 ( .A(n36656), .B(n36718), .Z(n36660) );
  XOR U808 ( .A(n35924), .B(n35986), .Z(n35928) );
  XOR U809 ( .A(n35168), .B(n35230), .Z(n35172) );
  XOR U810 ( .A(n34388), .B(n34450), .Z(n34392) );
  XOR U811 ( .A(n33584), .B(n33646), .Z(n33588) );
  XOR U812 ( .A(n32756), .B(n32818), .Z(n32760) );
  XOR U813 ( .A(n31904), .B(n31966), .Z(n31908) );
  XOR U814 ( .A(n31028), .B(n31090), .Z(n31032) );
  XOR U815 ( .A(n30128), .B(n30190), .Z(n30132) );
  XOR U816 ( .A(n29204), .B(n29266), .Z(n29208) );
  XOR U817 ( .A(n28256), .B(n28318), .Z(n28260) );
  XOR U818 ( .A(n27284), .B(n27346), .Z(n27288) );
  XOR U819 ( .A(n26286), .B(n26348), .Z(n26290) );
  XOR U820 ( .A(n25264), .B(n25326), .Z(n25268) );
  XOR U821 ( .A(n24216), .B(n24278), .Z(n24220) );
  XOR U822 ( .A(n23147), .B(n23209), .Z(n23151) );
  XOR U823 ( .A(n22054), .B(n22116), .Z(n22058) );
  XOR U824 ( .A(n20937), .B(n20999), .Z(n20941) );
  XOR U825 ( .A(n19797), .B(n19859), .Z(n19801) );
  XOR U826 ( .A(n47098), .B(n47154), .Z(n47102) );
  XOR U827 ( .A(n46954), .B(n47010), .Z(n46958) );
  XOR U828 ( .A(n2666), .B(n2723), .Z(n2670) );
  XOR U829 ( .A(n46883), .B(n46927), .Z(n46887) );
  XOR U830 ( .A(n46703), .B(n46747), .Z(n46707) );
  XOR U831 ( .A(n46499), .B(n46543), .Z(n46503) );
  XOR U832 ( .A(n46271), .B(n46315), .Z(n46275) );
  XOR U833 ( .A(n46019), .B(n46063), .Z(n46023) );
  XOR U834 ( .A(n45743), .B(n45787), .Z(n45747) );
  XOR U835 ( .A(n45443), .B(n45487), .Z(n45447) );
  XOR U836 ( .A(n45119), .B(n45163), .Z(n45123) );
  XOR U837 ( .A(n44771), .B(n44815), .Z(n44775) );
  XOR U838 ( .A(n44399), .B(n44443), .Z(n44403) );
  XOR U839 ( .A(n44003), .B(n44047), .Z(n44007) );
  XOR U840 ( .A(n43583), .B(n43627), .Z(n43587) );
  XOR U841 ( .A(n43139), .B(n43183), .Z(n43143) );
  XOR U842 ( .A(n42671), .B(n42715), .Z(n42675) );
  XOR U843 ( .A(n42179), .B(n42223), .Z(n42183) );
  XOR U844 ( .A(n41663), .B(n41707), .Z(n41667) );
  XOR U845 ( .A(n41123), .B(n41167), .Z(n41127) );
  XOR U846 ( .A(n40559), .B(n40603), .Z(n40563) );
  XOR U847 ( .A(n39971), .B(n40015), .Z(n39975) );
  XOR U848 ( .A(n39359), .B(n39403), .Z(n39363) );
  XOR U849 ( .A(n38723), .B(n38767), .Z(n38727) );
  XOR U850 ( .A(n38063), .B(n38107), .Z(n38067) );
  XOR U851 ( .A(n37379), .B(n37423), .Z(n37383) );
  XOR U852 ( .A(n36671), .B(n36715), .Z(n36675) );
  XOR U853 ( .A(n35939), .B(n35983), .Z(n35943) );
  XOR U854 ( .A(n35183), .B(n35227), .Z(n35187) );
  XOR U855 ( .A(n34403), .B(n34447), .Z(n34407) );
  XOR U856 ( .A(n33599), .B(n33643), .Z(n33603) );
  XOR U857 ( .A(n32771), .B(n32815), .Z(n32775) );
  XOR U858 ( .A(n31919), .B(n31963), .Z(n31923) );
  XOR U859 ( .A(n31043), .B(n31087), .Z(n31047) );
  XOR U860 ( .A(n30143), .B(n30187), .Z(n30147) );
  XOR U861 ( .A(n29219), .B(n29263), .Z(n29223) );
  XOR U862 ( .A(n28271), .B(n28315), .Z(n28275) );
  XOR U863 ( .A(n27299), .B(n27343), .Z(n27303) );
  XOR U864 ( .A(n26301), .B(n26345), .Z(n26305) );
  XOR U865 ( .A(n25279), .B(n25323), .Z(n25283) );
  XOR U866 ( .A(n24231), .B(n24275), .Z(n24235) );
  XOR U867 ( .A(n23162), .B(n23206), .Z(n23166) );
  XOR U868 ( .A(n22069), .B(n22113), .Z(n22073) );
  XOR U869 ( .A(n20952), .B(n20996), .Z(n20956) );
  XOR U870 ( .A(n19812), .B(n19856), .Z(n19816) );
  XOR U871 ( .A(n47232), .B(n47270), .Z(n47236) );
  XOR U872 ( .A(n47377), .B(n47403), .Z(n47381) );
  XOR U873 ( .A(n47186), .B(n47211), .Z(n47190) );
  XOR U874 ( .A(n47054), .B(n47080), .Z(n47058) );
  XOR U875 ( .A(n46898), .B(n46924), .Z(n46902) );
  XOR U876 ( .A(n46718), .B(n46744), .Z(n46722) );
  XOR U877 ( .A(n46514), .B(n46540), .Z(n46518) );
  XOR U878 ( .A(n46286), .B(n46312), .Z(n46290) );
  XOR U879 ( .A(n46034), .B(n46060), .Z(n46038) );
  XOR U880 ( .A(n45758), .B(n45784), .Z(n45762) );
  XOR U881 ( .A(n45458), .B(n45484), .Z(n45462) );
  XOR U882 ( .A(n45134), .B(n45160), .Z(n45138) );
  XOR U883 ( .A(n44786), .B(n44812), .Z(n44790) );
  XOR U884 ( .A(n44414), .B(n44440), .Z(n44418) );
  XOR U885 ( .A(n44018), .B(n44044), .Z(n44022) );
  XOR U886 ( .A(n43598), .B(n43624), .Z(n43602) );
  XOR U887 ( .A(n43154), .B(n43180), .Z(n43158) );
  XOR U888 ( .A(n42686), .B(n42712), .Z(n42690) );
  XOR U889 ( .A(n42194), .B(n42220), .Z(n42198) );
  XOR U890 ( .A(n41678), .B(n41704), .Z(n41682) );
  XOR U891 ( .A(n41138), .B(n41164), .Z(n41142) );
  XOR U892 ( .A(n40574), .B(n40600), .Z(n40578) );
  XOR U893 ( .A(n39986), .B(n40012), .Z(n39990) );
  XOR U894 ( .A(n39374), .B(n39400), .Z(n39378) );
  XOR U895 ( .A(n38738), .B(n38764), .Z(n38742) );
  XOR U896 ( .A(n38078), .B(n38104), .Z(n38082) );
  XOR U897 ( .A(n37394), .B(n37420), .Z(n37398) );
  XOR U898 ( .A(n36686), .B(n36712), .Z(n36690) );
  XOR U899 ( .A(n35954), .B(n35980), .Z(n35958) );
  XOR U900 ( .A(n35198), .B(n35224), .Z(n35202) );
  XOR U901 ( .A(n34418), .B(n34444), .Z(n34422) );
  XOR U902 ( .A(n33614), .B(n33640), .Z(n33618) );
  XOR U903 ( .A(n32786), .B(n32812), .Z(n32790) );
  XOR U904 ( .A(n31934), .B(n31960), .Z(n31938) );
  XOR U905 ( .A(n31058), .B(n31084), .Z(n31062) );
  XOR U906 ( .A(n30158), .B(n30184), .Z(n30162) );
  XOR U907 ( .A(n29234), .B(n29260), .Z(n29238) );
  XOR U908 ( .A(n28286), .B(n28312), .Z(n28290) );
  XOR U909 ( .A(n27314), .B(n27340), .Z(n27318) );
  XOR U910 ( .A(n26316), .B(n26342), .Z(n26320) );
  XOR U911 ( .A(n25294), .B(n25320), .Z(n25298) );
  XOR U912 ( .A(n24246), .B(n24272), .Z(n24250) );
  XOR U913 ( .A(n23177), .B(n23203), .Z(n23181) );
  XOR U914 ( .A(n22084), .B(n22110), .Z(n22088) );
  XOR U915 ( .A(n20967), .B(n20993), .Z(n20971) );
  XOR U916 ( .A(n19827), .B(n19853), .Z(n19831) );
  XOR U917 ( .A(n28393), .B(n28863), .Z(n28397) );
  XOR U918 ( .A(n27433), .B(n27903), .Z(n27437) );
  XOR U919 ( .A(n26432), .B(n26922), .Z(n26436) );
  XNOR U920 ( .A(n26960), .B(n26460), .Z(n26462) );
  XOR U921 ( .A(n29344), .B(n29796), .Z(n29348) );
  XOR U922 ( .A(n28408), .B(n28860), .Z(n28412) );
  XOR U923 ( .A(n24888), .B(n25402), .Z(n24892) );
  XOR U924 ( .A(n26447), .B(n26919), .Z(n26451) );
  XOR U925 ( .A(n27941), .B(n28381), .Z(n27945) );
  XOR U926 ( .A(n26969), .B(n27409), .Z(n26973) );
  XOR U927 ( .A(n24918), .B(n25396), .Z(n24922) );
  XOR U928 ( .A(n25423), .B(n25912), .Z(n25427) );
  XOR U929 ( .A(n31159), .B(n31593), .Z(n31163) );
  XOR U930 ( .A(n30271), .B(n30705), .Z(n30275) );
  XOR U931 ( .A(n25966), .B(n26412), .Z(n25970) );
  XOR U932 ( .A(n24371), .B(n24880), .Z(n24375) );
  XOR U933 ( .A(n24421), .B(n24870), .Z(n24425) );
  XOR U934 ( .A(n29828), .B(n30250), .Z(n29832) );
  XOR U935 ( .A(n28904), .B(n29326), .Z(n28908) );
  XOR U936 ( .A(n27956), .B(n28378), .Z(n27960) );
  XOR U937 ( .A(n26984), .B(n27406), .Z(n26988) );
  XOR U938 ( .A(n25986), .B(n26408), .Z(n25990) );
  XOR U939 ( .A(n23866), .B(n24348), .Z(n23870) );
  XOR U940 ( .A(n23350), .B(n23814), .Z(n23354) );
  XOR U941 ( .A(n32038), .B(n32454), .Z(n32042) );
  XOR U942 ( .A(n31174), .B(n31590), .Z(n31178) );
  XOR U943 ( .A(n24406), .B(n24873), .Z(n24410) );
  XOR U944 ( .A(n23851), .B(n24351), .Z(n23855) );
  XOR U945 ( .A(n22762), .B(n23287), .Z(n22766) );
  XOR U946 ( .A(n21089), .B(n21643), .Z(n21093) );
  XOR U947 ( .A(n24436), .B(n24867), .Z(n24440) );
  XOR U948 ( .A(n30743), .B(n31147), .Z(n30747) );
  XOR U949 ( .A(n29843), .B(n30247), .Z(n29847) );
  XOR U950 ( .A(n28919), .B(n29323), .Z(n28923) );
  XOR U951 ( .A(n27971), .B(n28375), .Z(n27975) );
  XOR U952 ( .A(n26999), .B(n27403), .Z(n27003) );
  XOR U953 ( .A(n26001), .B(n26405), .Z(n26005) );
  XOR U954 ( .A(n24978), .B(n25383), .Z(n24982) );
  XOR U955 ( .A(n22792), .B(n23281), .Z(n22796) );
  XOR U956 ( .A(n33709), .B(n34107), .Z(n33713) );
  XOR U957 ( .A(n32893), .B(n33291), .Z(n32897) );
  XOR U958 ( .A(n23390), .B(n23806), .Z(n23394) );
  XNOR U959 ( .A(n23341), .B(n22800), .Z(n22802) );
  XOR U960 ( .A(n21684), .B(n22190), .Z(n21688) );
  XOR U961 ( .A(n20547), .B(n21078), .Z(n20551) );
  XOR U962 ( .A(n22223), .B(n22742), .Z(n22227) );
  XOR U963 ( .A(n22268), .B(n22733), .Z(n22272) );
  XOR U964 ( .A(n21734), .B(n22180), .Z(n21738) );
  XOR U965 ( .A(n20532), .B(n21081), .Z(n20536) );
  XOR U966 ( .A(n19372), .B(n19944), .Z(n19376) );
  XOR U967 ( .A(n23375), .B(n23809), .Z(n23379) );
  XOR U968 ( .A(n21149), .B(n21631), .Z(n21153) );
  XOR U969 ( .A(n22318), .B(n22723), .Z(n22322) );
  XOR U970 ( .A(n32486), .B(n32872), .Z(n32490) );
  XOR U971 ( .A(n31634), .B(n32020), .Z(n31638) );
  XOR U972 ( .A(n30758), .B(n31144), .Z(n30762) );
  XOR U973 ( .A(n29858), .B(n30244), .Z(n29862) );
  XOR U974 ( .A(n28934), .B(n29320), .Z(n28938) );
  XOR U975 ( .A(n27986), .B(n28372), .Z(n27990) );
  XOR U976 ( .A(n27014), .B(n27400), .Z(n27018) );
  XOR U977 ( .A(n26016), .B(n26402), .Z(n26020) );
  XOR U978 ( .A(n24994), .B(n25380), .Z(n24998) );
  XOR U979 ( .A(n23415), .B(n23801), .Z(n23419) );
  XOR U980 ( .A(n23941), .B(n24333), .Z(n23945) );
  XOR U981 ( .A(n34903), .B(n35283), .Z(n34907) );
  XOR U982 ( .A(n34123), .B(n34503), .Z(n34127) );
  XOR U983 ( .A(n22857), .B(n23268), .Z(n22861) );
  XOR U984 ( .A(n21134), .B(n21634), .Z(n21138) );
  XNOR U985 ( .A(n19981), .B(n19405), .Z(n19407) );
  XOR U986 ( .A(n18813), .B(n19361), .Z(n18817) );
  XOR U987 ( .A(n21794), .B(n22168), .Z(n21798) );
  XOR U988 ( .A(n21749), .B(n22177), .Z(n21753) );
  XOR U989 ( .A(n19387), .B(n19941), .Z(n19391) );
  XOR U990 ( .A(n21164), .B(n21628), .Z(n21168) );
  XOR U991 ( .A(n19432), .B(n19932), .Z(n19436) );
  XOR U992 ( .A(n21774), .B(n22172), .Z(n21778) );
  XOR U993 ( .A(n33734), .B(n34102), .Z(n33738) );
  XOR U994 ( .A(n32918), .B(n33286), .Z(n32922) );
  XOR U995 ( .A(n32078), .B(n32446), .Z(n32082) );
  XOR U996 ( .A(n31214), .B(n31582), .Z(n31218) );
  XOR U997 ( .A(n30326), .B(n30694), .Z(n30330) );
  XOR U998 ( .A(n29414), .B(n29782), .Z(n29418) );
  XOR U999 ( .A(n28478), .B(n28846), .Z(n28482) );
  XOR U1000 ( .A(n27518), .B(n27886), .Z(n27522) );
  XOR U1001 ( .A(n26532), .B(n26900), .Z(n26536) );
  XOR U1002 ( .A(n25523), .B(n25891), .Z(n25527) );
  XOR U1003 ( .A(n24486), .B(n24854), .Z(n24490) );
  XOR U1004 ( .A(n23430), .B(n23798), .Z(n23434) );
  XOR U1005 ( .A(n20617), .B(n21064), .Z(n20621) );
  XNOR U1006 ( .A(n23436), .B(n22895), .Z(n22897) );
  XOR U1007 ( .A(n35674), .B(n36036), .Z(n35678) );
  XOR U1008 ( .A(n34918), .B(n35280), .Z(n34922) );
  XOR U1009 ( .A(n19462), .B(n19926), .Z(n19466) );
  XOR U1010 ( .A(n19417), .B(n19935), .Z(n19421) );
  XOR U1011 ( .A(n20672), .B(n21053), .Z(n20676) );
  XOR U1012 ( .A(n16919), .B(n17486), .Z(n16923) );
  XOR U1013 ( .A(n19447), .B(n19929), .Z(n19451) );
  XOR U1014 ( .A(n17552), .B(n18077), .Z(n17556) );
  XOR U1015 ( .A(n21224), .B(n21616), .Z(n21228) );
  XOR U1016 ( .A(n18903), .B(n19343), .Z(n18907) );
  XOR U1017 ( .A(n34541), .B(n34891), .Z(n34545) );
  XOR U1018 ( .A(n33749), .B(n34099), .Z(n33753) );
  XOR U1019 ( .A(n32933), .B(n33283), .Z(n32937) );
  XOR U1020 ( .A(n32093), .B(n32443), .Z(n32097) );
  XOR U1021 ( .A(n31229), .B(n31579), .Z(n31233) );
  XOR U1022 ( .A(n30341), .B(n30691), .Z(n30345) );
  XOR U1023 ( .A(n29429), .B(n29779), .Z(n29433) );
  XOR U1024 ( .A(n28493), .B(n28843), .Z(n28497) );
  XOR U1025 ( .A(n27533), .B(n27883), .Z(n27537) );
  XOR U1026 ( .A(n26547), .B(n26897), .Z(n26551) );
  XOR U1027 ( .A(n25538), .B(n25888), .Z(n25542) );
  XOR U1028 ( .A(n24501), .B(n24851), .Z(n24505) );
  XOR U1029 ( .A(n23445), .B(n23795), .Z(n23449) );
  XOR U1030 ( .A(n22363), .B(n22713), .Z(n22367) );
  XOR U1031 ( .A(n20632), .B(n21061), .Z(n20636) );
  XOR U1032 ( .A(n16904), .B(n17489), .Z(n16908) );
  XOR U1033 ( .A(n19497), .B(n19919), .Z(n19501) );
  XNOR U1034 ( .A(n20698), .B(n20128), .Z(n20130) );
  XOR U1035 ( .A(n37129), .B(n37473), .Z(n37133) );
  XOR U1036 ( .A(n36421), .B(n36765), .Z(n36425) );
  XOR U1037 ( .A(n21254), .B(n21610), .Z(n21258) );
  XOR U1038 ( .A(n19477), .B(n19923), .Z(n19481) );
  XNOR U1039 ( .A(n20081), .B(n19505), .Z(n19507) );
  XOR U1040 ( .A(n19527), .B(n19913), .Z(n19531) );
  XOR U1041 ( .A(n17587), .B(n18070), .Z(n17591) );
  XOR U1042 ( .A(n16934), .B(n17483), .Z(n16938) );
  XOR U1043 ( .A(n15074), .B(n15659), .Z(n15078) );
  XOR U1044 ( .A(n17567), .B(n18074), .Z(n17571) );
  XOR U1045 ( .A(n15725), .B(n16268), .Z(n15729) );
  XOR U1046 ( .A(n20090), .B(n20488), .Z(n20094) );
  XOR U1047 ( .A(n36068), .B(n36400), .Z(n36072) );
  XOR U1048 ( .A(n35324), .B(n35656), .Z(n35328) );
  XOR U1049 ( .A(n34556), .B(n34888), .Z(n34560) );
  XOR U1050 ( .A(n33764), .B(n34096), .Z(n33768) );
  XOR U1051 ( .A(n32948), .B(n33280), .Z(n32952) );
  XOR U1052 ( .A(n32108), .B(n32440), .Z(n32112) );
  XOR U1053 ( .A(n31244), .B(n31576), .Z(n31248) );
  XOR U1054 ( .A(n30356), .B(n30688), .Z(n30360) );
  XOR U1055 ( .A(n29444), .B(n29776), .Z(n29448) );
  XOR U1056 ( .A(n28508), .B(n28840), .Z(n28512) );
  XOR U1057 ( .A(n27548), .B(n27880), .Z(n27552) );
  XOR U1058 ( .A(n26562), .B(n26894), .Z(n26566) );
  XOR U1059 ( .A(n25553), .B(n25885), .Z(n25557) );
  XOR U1060 ( .A(n24516), .B(n24848), .Z(n24520) );
  XOR U1061 ( .A(n23460), .B(n23792), .Z(n23464) );
  XOR U1062 ( .A(n22378), .B(n22710), .Z(n22382) );
  XOR U1063 ( .A(n21274), .B(n21606), .Z(n21278) );
  XNOR U1064 ( .A(n20111), .B(n19535), .Z(n19537) );
  XOR U1065 ( .A(n15059), .B(n15662), .Z(n15063) );
  XOR U1066 ( .A(n19557), .B(n19907), .Z(n19561) );
  XOR U1067 ( .A(n37828), .B(n38154), .Z(n37832) );
  XOR U1068 ( .A(n37144), .B(n37470), .Z(n37148) );
  XOR U1069 ( .A(n18993), .B(n19325), .Z(n18997) );
  XOR U1070 ( .A(n20120), .B(n20482), .Z(n20124) );
  XOR U1071 ( .A(n15755), .B(n16262), .Z(n15759) );
  XNOR U1072 ( .A(n20718), .B(n20148), .Z(n20150) );
  XNOR U1073 ( .A(n20141), .B(n19565), .Z(n19567) );
  XOR U1074 ( .A(n15089), .B(n15656), .Z(n15093) );
  XOR U1075 ( .A(n13175), .B(n13778), .Z(n13179) );
  XOR U1076 ( .A(n15740), .B(n16265), .Z(n15744) );
  XOR U1077 ( .A(n13844), .B(n14405), .Z(n13848) );
  XOR U1078 ( .A(n36803), .B(n37117), .Z(n36807) );
  XOR U1079 ( .A(n36083), .B(n36397), .Z(n36087) );
  XOR U1080 ( .A(n35339), .B(n35653), .Z(n35343) );
  XOR U1081 ( .A(n34571), .B(n34885), .Z(n34575) );
  XOR U1082 ( .A(n33779), .B(n34093), .Z(n33783) );
  XOR U1083 ( .A(n32963), .B(n33277), .Z(n32967) );
  XOR U1084 ( .A(n32123), .B(n32437), .Z(n32127) );
  XOR U1085 ( .A(n31259), .B(n31573), .Z(n31263) );
  XOR U1086 ( .A(n30371), .B(n30685), .Z(n30375) );
  XOR U1087 ( .A(n29459), .B(n29773), .Z(n29463) );
  XOR U1088 ( .A(n28523), .B(n28837), .Z(n28527) );
  XOR U1089 ( .A(n27563), .B(n27877), .Z(n27567) );
  XOR U1090 ( .A(n26577), .B(n26891), .Z(n26581) );
  XOR U1091 ( .A(n25568), .B(n25882), .Z(n25572) );
  XOR U1092 ( .A(n24531), .B(n24845), .Z(n24535) );
  XOR U1093 ( .A(n23475), .B(n23789), .Z(n23479) );
  XOR U1094 ( .A(n22393), .B(n22707), .Z(n22397) );
  XOR U1095 ( .A(n21289), .B(n21603), .Z(n21293) );
  XOR U1096 ( .A(n20160), .B(n20474), .Z(n20164) );
  XNOR U1097 ( .A(n20166), .B(n19590), .Z(n19592) );
  XOR U1098 ( .A(n13160), .B(n13781), .Z(n13164) );
  XOR U1099 ( .A(n39139), .B(n39447), .Z(n39143) );
  XOR U1100 ( .A(n38503), .B(n38811), .Z(n38507) );
  XOR U1101 ( .A(n13874), .B(n14399), .Z(n13878) );
  XOR U1102 ( .A(n13190), .B(n13775), .Z(n13194) );
  XOR U1103 ( .A(n11220), .B(n11841), .Z(n11224) );
  XOR U1104 ( .A(n13859), .B(n14402), .Z(n13863) );
  XOR U1105 ( .A(n11907), .B(n12488), .Z(n11911) );
  XOR U1106 ( .A(n38186), .B(n38482), .Z(n38190) );
  XOR U1107 ( .A(n37514), .B(n37810), .Z(n37518) );
  XOR U1108 ( .A(n36818), .B(n37114), .Z(n36822) );
  XOR U1109 ( .A(n36098), .B(n36394), .Z(n36102) );
  XOR U1110 ( .A(n35354), .B(n35650), .Z(n35358) );
  XOR U1111 ( .A(n34586), .B(n34882), .Z(n34590) );
  XOR U1112 ( .A(n33794), .B(n34090), .Z(n33798) );
  XOR U1113 ( .A(n32978), .B(n33274), .Z(n32982) );
  XOR U1114 ( .A(n32138), .B(n32434), .Z(n32142) );
  XOR U1115 ( .A(n31274), .B(n31570), .Z(n31278) );
  XOR U1116 ( .A(n30386), .B(n30682), .Z(n30390) );
  XOR U1117 ( .A(n29474), .B(n29770), .Z(n29478) );
  XOR U1118 ( .A(n28538), .B(n28834), .Z(n28542) );
  XOR U1119 ( .A(n27578), .B(n27874), .Z(n27582) );
  XOR U1120 ( .A(n26592), .B(n26888), .Z(n26596) );
  XOR U1121 ( .A(n25583), .B(n25879), .Z(n25587) );
  XOR U1122 ( .A(n24546), .B(n24842), .Z(n24550) );
  XOR U1123 ( .A(n23490), .B(n23786), .Z(n23494) );
  XOR U1124 ( .A(n22408), .B(n22704), .Z(n22412) );
  XOR U1125 ( .A(n21304), .B(n21600), .Z(n21308) );
  XOR U1126 ( .A(n20175), .B(n20471), .Z(n20179) );
  XOR U1127 ( .A(n19023), .B(n19319), .Z(n19027) );
  XOR U1128 ( .A(n11205), .B(n11844), .Z(n11209) );
  XOR U1129 ( .A(n39766), .B(n40056), .Z(n39770) );
  XOR U1130 ( .A(n39154), .B(n39444), .Z(n39158) );
  XOR U1131 ( .A(n13245), .B(n13764), .Z(n13249) );
  XOR U1132 ( .A(n12620), .B(n13121), .Z(n12624) );
  XOR U1133 ( .A(n11280), .B(n11829), .Z(n11284) );
  XOR U1134 ( .A(n11235), .B(n11838), .Z(n11239) );
  XOR U1135 ( .A(n10592), .B(n11177), .Z(n10596) );
  XOR U1136 ( .A(n38849), .B(n39127), .Z(n38853) );
  XOR U1137 ( .A(n38201), .B(n38479), .Z(n38205) );
  XOR U1138 ( .A(n37529), .B(n37807), .Z(n37533) );
  XOR U1139 ( .A(n36833), .B(n37111), .Z(n36837) );
  XOR U1140 ( .A(n36113), .B(n36391), .Z(n36117) );
  XOR U1141 ( .A(n35369), .B(n35647), .Z(n35373) );
  XOR U1142 ( .A(n34601), .B(n34879), .Z(n34605) );
  XOR U1143 ( .A(n33809), .B(n34087), .Z(n33813) );
  XOR U1144 ( .A(n32993), .B(n33271), .Z(n32997) );
  XOR U1145 ( .A(n32153), .B(n32431), .Z(n32157) );
  XOR U1146 ( .A(n31289), .B(n31567), .Z(n31293) );
  XOR U1147 ( .A(n30401), .B(n30679), .Z(n30405) );
  XOR U1148 ( .A(n29489), .B(n29767), .Z(n29493) );
  XOR U1149 ( .A(n28553), .B(n28831), .Z(n28557) );
  XOR U1150 ( .A(n27593), .B(n27871), .Z(n27597) );
  XOR U1151 ( .A(n26607), .B(n26885), .Z(n26611) );
  XOR U1152 ( .A(n25598), .B(n25876), .Z(n25602) );
  XOR U1153 ( .A(n24561), .B(n24839), .Z(n24565) );
  XOR U1154 ( .A(n23505), .B(n23783), .Z(n23509) );
  XOR U1155 ( .A(n22423), .B(n22701), .Z(n22427) );
  XOR U1156 ( .A(n21319), .B(n21597), .Z(n21323) );
  XOR U1157 ( .A(n20190), .B(n20468), .Z(n20194) );
  XOR U1158 ( .A(n19038), .B(n19316), .Z(n19042) );
  XOR U1159 ( .A(n12650), .B(n13115), .Z(n12654) );
  XOR U1160 ( .A(n8532), .B(n9177), .Z(n8536) );
  XOR U1161 ( .A(n9198), .B(n9855), .Z(n9202) );
  XOR U1162 ( .A(n9243), .B(n9846), .Z(n9247) );
  XOR U1163 ( .A(n40933), .B(n41205), .Z(n40937) );
  XOR U1164 ( .A(n40369), .B(n40641), .Z(n40373) );
  XOR U1165 ( .A(n17762), .B(n18035), .Z(n17766) );
  XOR U1166 ( .A(n11977), .B(n12474), .Z(n11981) );
  XOR U1167 ( .A(n12680), .B(n13109), .Z(n12684) );
  XOR U1168 ( .A(n9273), .B(n9840), .Z(n9277) );
  XOR U1169 ( .A(n9228), .B(n9849), .Z(n9232) );
  XOR U1170 ( .A(n40088), .B(n40348), .Z(n40092) );
  XOR U1171 ( .A(n39488), .B(n39748), .Z(n39492) );
  XOR U1172 ( .A(n38864), .B(n39124), .Z(n38868) );
  XOR U1173 ( .A(n38216), .B(n38476), .Z(n38220) );
  XOR U1174 ( .A(n37544), .B(n37804), .Z(n37548) );
  XOR U1175 ( .A(n36848), .B(n37108), .Z(n36852) );
  XOR U1176 ( .A(n36128), .B(n36388), .Z(n36132) );
  XOR U1177 ( .A(n35384), .B(n35644), .Z(n35388) );
  XOR U1178 ( .A(n34616), .B(n34876), .Z(n34620) );
  XOR U1179 ( .A(n33824), .B(n34084), .Z(n33828) );
  XOR U1180 ( .A(n33008), .B(n33268), .Z(n33012) );
  XOR U1181 ( .A(n32168), .B(n32428), .Z(n32172) );
  XOR U1182 ( .A(n31304), .B(n31564), .Z(n31308) );
  XOR U1183 ( .A(n30416), .B(n30676), .Z(n30420) );
  XOR U1184 ( .A(n29504), .B(n29764), .Z(n29508) );
  XOR U1185 ( .A(n28568), .B(n28828), .Z(n28572) );
  XOR U1186 ( .A(n27608), .B(n27868), .Z(n27612) );
  XOR U1187 ( .A(n26622), .B(n26882), .Z(n26626) );
  XOR U1188 ( .A(n25613), .B(n25873), .Z(n25617) );
  XOR U1189 ( .A(n24576), .B(n24836), .Z(n24580) );
  XOR U1190 ( .A(n23520), .B(n23780), .Z(n23524) );
  XOR U1191 ( .A(n22438), .B(n22698), .Z(n22442) );
  XOR U1192 ( .A(n21334), .B(n21594), .Z(n21338) );
  XOR U1193 ( .A(n20205), .B(n20465), .Z(n20209) );
  XOR U1194 ( .A(n19053), .B(n19313), .Z(n19057) );
  XOR U1195 ( .A(n16565), .B(n16832), .Z(n16569) );
  XOR U1196 ( .A(n12710), .B(n13103), .Z(n12714) );
  XOR U1197 ( .A(n12007), .B(n12468), .Z(n12011) );
  XOR U1198 ( .A(n10632), .B(n11169), .Z(n10636) );
  XOR U1199 ( .A(n7137), .B(n7812), .Z(n7141) );
  XOR U1200 ( .A(n7182), .B(n7803), .Z(n7186) );
  XOR U1201 ( .A(n9303), .B(n9834), .Z(n9307) );
  XOR U1202 ( .A(n41488), .B(n41742), .Z(n41492) );
  XOR U1203 ( .A(n40948), .B(n41202), .Z(n40952) );
  XOR U1204 ( .A(n7162), .B(n7807), .Z(n7166) );
  XOR U1205 ( .A(n8577), .B(n9168), .Z(n8581) );
  XOR U1206 ( .A(n10662), .B(n11163), .Z(n10666) );
  XOR U1207 ( .A(n12037), .B(n12462), .Z(n12041) );
  XOR U1208 ( .A(n12740), .B(n13097), .Z(n12744) );
  XOR U1209 ( .A(n17184), .B(n17433), .Z(n17188) );
  XOR U1210 ( .A(n15970), .B(n16219), .Z(n15974) );
  XOR U1211 ( .A(n9333), .B(n9828), .Z(n9337) );
  XOR U1212 ( .A(n7212), .B(n7797), .Z(n7216) );
  XOR U1213 ( .A(n40679), .B(n40921), .Z(n40683) );
  XOR U1214 ( .A(n40103), .B(n40345), .Z(n40107) );
  XOR U1215 ( .A(n39503), .B(n39745), .Z(n39507) );
  XOR U1216 ( .A(n38879), .B(n39121), .Z(n38883) );
  XOR U1217 ( .A(n38231), .B(n38473), .Z(n38235) );
  XOR U1218 ( .A(n37559), .B(n37801), .Z(n37563) );
  XOR U1219 ( .A(n36863), .B(n37105), .Z(n36867) );
  XOR U1220 ( .A(n36143), .B(n36385), .Z(n36147) );
  XOR U1221 ( .A(n35399), .B(n35641), .Z(n35403) );
  XOR U1222 ( .A(n34631), .B(n34873), .Z(n34635) );
  XOR U1223 ( .A(n33839), .B(n34081), .Z(n33843) );
  XOR U1224 ( .A(n33023), .B(n33265), .Z(n33027) );
  XOR U1225 ( .A(n32183), .B(n32425), .Z(n32187) );
  XOR U1226 ( .A(n31319), .B(n31561), .Z(n31323) );
  XOR U1227 ( .A(n30431), .B(n30673), .Z(n30435) );
  XOR U1228 ( .A(n29519), .B(n29761), .Z(n29523) );
  XOR U1229 ( .A(n28583), .B(n28825), .Z(n28587) );
  XOR U1230 ( .A(n27623), .B(n27865), .Z(n27627) );
  XOR U1231 ( .A(n26637), .B(n26879), .Z(n26641) );
  XOR U1232 ( .A(n25628), .B(n25870), .Z(n25632) );
  XOR U1233 ( .A(n24591), .B(n24833), .Z(n24595) );
  XOR U1234 ( .A(n23535), .B(n23777), .Z(n23539) );
  XOR U1235 ( .A(n22453), .B(n22695), .Z(n22457) );
  XOR U1236 ( .A(n21349), .B(n21591), .Z(n21353) );
  XOR U1237 ( .A(n20220), .B(n20462), .Z(n20224) );
  XOR U1238 ( .A(n19068), .B(n19310), .Z(n19072) );
  XOR U1239 ( .A(n12770), .B(n13091), .Z(n12774) );
  XOR U1240 ( .A(n12067), .B(n12456), .Z(n12071) );
  XOR U1241 ( .A(n10692), .B(n11157), .Z(n10696) );
  XOR U1242 ( .A(n8607), .B(n9162), .Z(n8611) );
  XOR U1243 ( .A(n5040), .B(n5711), .Z(n5044) );
  XOR U1244 ( .A(n5020), .B(n5715), .Z(n5024) );
  XOR U1245 ( .A(n5065), .B(n5706), .Z(n5069) );
  XOR U1246 ( .A(n7242), .B(n7791), .Z(n7246) );
  XOR U1247 ( .A(n9363), .B(n9822), .Z(n9367) );
  XOR U1248 ( .A(n42511), .B(n42747), .Z(n42515) );
  XOR U1249 ( .A(n42019), .B(n42255), .Z(n42023) );
  XOR U1250 ( .A(n6498), .B(n7107), .Z(n6502) );
  XOR U1251 ( .A(n8637), .B(n9156), .Z(n8641) );
  XOR U1252 ( .A(n10722), .B(n11151), .Z(n10726) );
  XOR U1253 ( .A(n12097), .B(n12450), .Z(n12101) );
  XOR U1254 ( .A(n12800), .B(n13085), .Z(n12804) );
  XOR U1255 ( .A(n9393), .B(n9816), .Z(n9397) );
  XOR U1256 ( .A(n7272), .B(n7785), .Z(n7276) );
  XOR U1257 ( .A(n5095), .B(n5700), .Z(n5099) );
  XOR U1258 ( .A(n2866), .B(n3559), .Z(n2870) );
  XOR U1259 ( .A(n15369), .B(n15600), .Z(n15373) );
  XOR U1260 ( .A(n41774), .B(n41998), .Z(n41778) );
  XOR U1261 ( .A(n41246), .B(n41470), .Z(n41250) );
  XOR U1262 ( .A(n40694), .B(n40918), .Z(n40698) );
  XOR U1263 ( .A(n40118), .B(n40342), .Z(n40122) );
  XOR U1264 ( .A(n39518), .B(n39742), .Z(n39522) );
  XOR U1265 ( .A(n38894), .B(n39118), .Z(n38898) );
  XOR U1266 ( .A(n38246), .B(n38470), .Z(n38250) );
  XOR U1267 ( .A(n37574), .B(n37798), .Z(n37578) );
  XOR U1268 ( .A(n36878), .B(n37102), .Z(n36882) );
  XOR U1269 ( .A(n36158), .B(n36382), .Z(n36162) );
  XOR U1270 ( .A(n35414), .B(n35638), .Z(n35418) );
  XOR U1271 ( .A(n34646), .B(n34870), .Z(n34650) );
  XOR U1272 ( .A(n33854), .B(n34078), .Z(n33858) );
  XOR U1273 ( .A(n33038), .B(n33262), .Z(n33042) );
  XOR U1274 ( .A(n32198), .B(n32422), .Z(n32202) );
  XOR U1275 ( .A(n31334), .B(n31558), .Z(n31338) );
  XOR U1276 ( .A(n30446), .B(n30670), .Z(n30450) );
  XOR U1277 ( .A(n29534), .B(n29758), .Z(n29538) );
  XOR U1278 ( .A(n28598), .B(n28822), .Z(n28602) );
  XOR U1279 ( .A(n27638), .B(n27862), .Z(n27642) );
  XOR U1280 ( .A(n26652), .B(n26876), .Z(n26656) );
  XOR U1281 ( .A(n25643), .B(n25867), .Z(n25647) );
  XOR U1282 ( .A(n24606), .B(n24830), .Z(n24610) );
  XOR U1283 ( .A(n23550), .B(n23774), .Z(n23554) );
  XOR U1284 ( .A(n22468), .B(n22692), .Z(n22472) );
  XOR U1285 ( .A(n21364), .B(n21588), .Z(n21368) );
  XOR U1286 ( .A(n20235), .B(n20459), .Z(n20239) );
  XOR U1287 ( .A(n19083), .B(n19307), .Z(n19087) );
  XOR U1288 ( .A(n12830), .B(n13079), .Z(n12834) );
  XOR U1289 ( .A(n12127), .B(n12444), .Z(n12131) );
  XOR U1290 ( .A(n10752), .B(n11145), .Z(n10756) );
  XOR U1291 ( .A(n8667), .B(n9150), .Z(n8671) );
  XOR U1292 ( .A(n6528), .B(n7101), .Z(n6532) );
  XOR U1293 ( .A(n2851), .B(n3562), .Z(n2855) );
  XOR U1294 ( .A(n2896), .B(n3553), .Z(n2900) );
  XOR U1295 ( .A(n5125), .B(n5694), .Z(n5129) );
  XOR U1296 ( .A(n7302), .B(n7779), .Z(n7306) );
  XOR U1297 ( .A(n9423), .B(n9810), .Z(n9427) );
  XOR U1298 ( .A(n42994), .B(n43212), .Z(n42998) );
  XOR U1299 ( .A(n42526), .B(n42744), .Z(n42530) );
  XOR U1300 ( .A(n4363), .B(n4990), .Z(n4367) );
  XOR U1301 ( .A(n6558), .B(n7095), .Z(n6562) );
  XOR U1302 ( .A(n8697), .B(n9144), .Z(n8701) );
  XOR U1303 ( .A(n10782), .B(n11139), .Z(n10786) );
  XOR U1304 ( .A(n12157), .B(n12438), .Z(n12161) );
  XOR U1305 ( .A(n14762), .B(n14975), .Z(n14766) );
  XOR U1306 ( .A(n9453), .B(n9804), .Z(n9457) );
  XOR U1307 ( .A(n7332), .B(n7773), .Z(n7336) );
  XOR U1308 ( .A(n5155), .B(n5688), .Z(n5159) );
  XOR U1309 ( .A(n2926), .B(n3547), .Z(n2930) );
  XOR U1310 ( .A(n42293), .B(n42499), .Z(n42297) );
  XOR U1311 ( .A(n41789), .B(n41995), .Z(n41793) );
  XOR U1312 ( .A(n41261), .B(n41467), .Z(n41265) );
  XOR U1313 ( .A(n40709), .B(n40915), .Z(n40713) );
  XOR U1314 ( .A(n40133), .B(n40339), .Z(n40137) );
  XOR U1315 ( .A(n39533), .B(n39739), .Z(n39537) );
  XOR U1316 ( .A(n38909), .B(n39115), .Z(n38913) );
  XOR U1317 ( .A(n38261), .B(n38467), .Z(n38265) );
  XOR U1318 ( .A(n37589), .B(n37795), .Z(n37593) );
  XOR U1319 ( .A(n36893), .B(n37099), .Z(n36897) );
  XOR U1320 ( .A(n36173), .B(n36379), .Z(n36177) );
  XOR U1321 ( .A(n35429), .B(n35635), .Z(n35433) );
  XOR U1322 ( .A(n34661), .B(n34867), .Z(n34665) );
  XOR U1323 ( .A(n33869), .B(n34075), .Z(n33873) );
  XOR U1324 ( .A(n33053), .B(n33259), .Z(n33057) );
  XOR U1325 ( .A(n32213), .B(n32419), .Z(n32217) );
  XOR U1326 ( .A(n31349), .B(n31555), .Z(n31353) );
  XOR U1327 ( .A(n30461), .B(n30667), .Z(n30465) );
  XOR U1328 ( .A(n29549), .B(n29755), .Z(n29553) );
  XOR U1329 ( .A(n28613), .B(n28819), .Z(n28617) );
  XOR U1330 ( .A(n27653), .B(n27859), .Z(n27657) );
  XOR U1331 ( .A(n26667), .B(n26873), .Z(n26671) );
  XOR U1332 ( .A(n25658), .B(n25864), .Z(n25662) );
  XOR U1333 ( .A(n24621), .B(n24827), .Z(n24625) );
  XOR U1334 ( .A(n23565), .B(n23771), .Z(n23569) );
  XOR U1335 ( .A(n22483), .B(n22689), .Z(n22487) );
  XOR U1336 ( .A(n21379), .B(n21585), .Z(n21383) );
  XOR U1337 ( .A(n20250), .B(n20456), .Z(n20254) );
  XOR U1338 ( .A(n19098), .B(n19304), .Z(n19102) );
  XOR U1339 ( .A(n13505), .B(n13712), .Z(n13509) );
  XOR U1340 ( .A(n12187), .B(n12432), .Z(n12191) );
  XOR U1341 ( .A(n10812), .B(n11133), .Z(n10816) );
  XOR U1342 ( .A(n8727), .B(n9138), .Z(n8731) );
  XOR U1343 ( .A(n6588), .B(n7089), .Z(n6592) );
  XOR U1344 ( .A(n4393), .B(n4984), .Z(n4397) );
  XOR U1345 ( .A(n2956), .B(n3541), .Z(n2960) );
  XOR U1346 ( .A(n5185), .B(n5682), .Z(n5189) );
  XOR U1347 ( .A(n7362), .B(n7767), .Z(n7366) );
  XOR U1348 ( .A(n9483), .B(n9798), .Z(n9487) );
  XOR U1349 ( .A(n43873), .B(n44073), .Z(n43877) );
  XOR U1350 ( .A(n43453), .B(n43653), .Z(n43457) );
  XOR U1351 ( .A(n12870), .B(n13071), .Z(n12874) );
  XOR U1352 ( .A(n4423), .B(n4978), .Z(n4427) );
  XOR U1353 ( .A(n6618), .B(n7083), .Z(n6622) );
  XOR U1354 ( .A(n8757), .B(n9132), .Z(n8761) );
  XOR U1355 ( .A(n10842), .B(n11127), .Z(n10846) );
  XOR U1356 ( .A(n9513), .B(n9792), .Z(n9517) );
  XOR U1357 ( .A(n7392), .B(n7761), .Z(n7396) );
  XOR U1358 ( .A(n5215), .B(n5676), .Z(n5219) );
  XOR U1359 ( .A(n2986), .B(n3535), .Z(n2990) );
  XOR U1360 ( .A(n43244), .B(n43432), .Z(n43248) );
  XOR U1361 ( .A(n42788), .B(n42976), .Z(n42792) );
  XOR U1362 ( .A(n42308), .B(n42496), .Z(n42312) );
  XOR U1363 ( .A(n41804), .B(n41992), .Z(n41808) );
  XOR U1364 ( .A(n41276), .B(n41464), .Z(n41280) );
  XOR U1365 ( .A(n40724), .B(n40912), .Z(n40728) );
  XOR U1366 ( .A(n40148), .B(n40336), .Z(n40152) );
  XOR U1367 ( .A(n39548), .B(n39736), .Z(n39552) );
  XOR U1368 ( .A(n38924), .B(n39112), .Z(n38928) );
  XOR U1369 ( .A(n38276), .B(n38464), .Z(n38280) );
  XOR U1370 ( .A(n37604), .B(n37792), .Z(n37608) );
  XOR U1371 ( .A(n36908), .B(n37096), .Z(n36912) );
  XOR U1372 ( .A(n36188), .B(n36376), .Z(n36192) );
  XOR U1373 ( .A(n35444), .B(n35632), .Z(n35448) );
  XOR U1374 ( .A(n34676), .B(n34864), .Z(n34680) );
  XOR U1375 ( .A(n33884), .B(n34072), .Z(n33888) );
  XOR U1376 ( .A(n33068), .B(n33256), .Z(n33072) );
  XOR U1377 ( .A(n32228), .B(n32416), .Z(n32232) );
  XOR U1378 ( .A(n31364), .B(n31552), .Z(n31368) );
  XOR U1379 ( .A(n30476), .B(n30664), .Z(n30480) );
  XOR U1380 ( .A(n29564), .B(n29752), .Z(n29568) );
  XOR U1381 ( .A(n28628), .B(n28816), .Z(n28632) );
  XOR U1382 ( .A(n27668), .B(n27856), .Z(n27672) );
  XOR U1383 ( .A(n26682), .B(n26870), .Z(n26686) );
  XOR U1384 ( .A(n25673), .B(n25861), .Z(n25677) );
  XOR U1385 ( .A(n24636), .B(n24824), .Z(n24640) );
  XOR U1386 ( .A(n23580), .B(n23768), .Z(n23584) );
  XOR U1387 ( .A(n22498), .B(n22686), .Z(n22502) );
  XOR U1388 ( .A(n21394), .B(n21582), .Z(n21398) );
  XOR U1389 ( .A(n20265), .B(n20453), .Z(n20269) );
  XOR U1390 ( .A(n19113), .B(n19301), .Z(n19117) );
  XOR U1391 ( .A(n11580), .B(n11769), .Z(n11584) );
  XOR U1392 ( .A(n10872), .B(n11121), .Z(n10876) );
  XOR U1393 ( .A(n8787), .B(n9126), .Z(n8791) );
  XOR U1394 ( .A(n6648), .B(n7077), .Z(n6652) );
  XOR U1395 ( .A(n4453), .B(n4972), .Z(n4457) );
  XOR U1396 ( .A(n3016), .B(n3529), .Z(n3020) );
  XOR U1397 ( .A(n5245), .B(n5670), .Z(n5249) );
  XOR U1398 ( .A(n7422), .B(n7755), .Z(n7426) );
  XOR U1399 ( .A(n12227), .B(n12424), .Z(n12231) );
  XOR U1400 ( .A(n9543), .B(n9786), .Z(n9547) );
  XOR U1401 ( .A(n44284), .B(n44466), .Z(n44288) );
  XOR U1402 ( .A(n43888), .B(n44070), .Z(n43892) );
  XOR U1403 ( .A(n4483), .B(n4966), .Z(n4487) );
  XOR U1404 ( .A(n6678), .B(n7071), .Z(n6682) );
  XOR U1405 ( .A(n8817), .B(n9120), .Z(n8821) );
  XOR U1406 ( .A(n10902), .B(n11115), .Z(n10906) );
  XOR U1407 ( .A(n9573), .B(n9780), .Z(n9577) );
  XOR U1408 ( .A(n7452), .B(n7749), .Z(n7456) );
  XOR U1409 ( .A(n5275), .B(n5664), .Z(n5279) );
  XOR U1410 ( .A(n3046), .B(n3523), .Z(n3050) );
  XOR U1411 ( .A(n43691), .B(n43861), .Z(n43695) );
  XOR U1412 ( .A(n43259), .B(n43429), .Z(n43263) );
  XOR U1413 ( .A(n42803), .B(n42973), .Z(n42807) );
  XOR U1414 ( .A(n42323), .B(n42493), .Z(n42327) );
  XOR U1415 ( .A(n41819), .B(n41989), .Z(n41823) );
  XOR U1416 ( .A(n41291), .B(n41461), .Z(n41295) );
  XOR U1417 ( .A(n40739), .B(n40909), .Z(n40743) );
  XOR U1418 ( .A(n40163), .B(n40333), .Z(n40167) );
  XOR U1419 ( .A(n39563), .B(n39733), .Z(n39567) );
  XOR U1420 ( .A(n38939), .B(n39109), .Z(n38943) );
  XOR U1421 ( .A(n38291), .B(n38461), .Z(n38295) );
  XOR U1422 ( .A(n37619), .B(n37789), .Z(n37623) );
  XOR U1423 ( .A(n36923), .B(n37093), .Z(n36927) );
  XOR U1424 ( .A(n36203), .B(n36373), .Z(n36207) );
  XOR U1425 ( .A(n35459), .B(n35629), .Z(n35463) );
  XOR U1426 ( .A(n34691), .B(n34861), .Z(n34695) );
  XOR U1427 ( .A(n33899), .B(n34069), .Z(n33903) );
  XOR U1428 ( .A(n33083), .B(n33253), .Z(n33087) );
  XOR U1429 ( .A(n32243), .B(n32413), .Z(n32247) );
  XOR U1430 ( .A(n31379), .B(n31549), .Z(n31383) );
  XOR U1431 ( .A(n30491), .B(n30661), .Z(n30495) );
  XOR U1432 ( .A(n29579), .B(n29749), .Z(n29583) );
  XOR U1433 ( .A(n28643), .B(n28813), .Z(n28647) );
  XOR U1434 ( .A(n27683), .B(n27853), .Z(n27687) );
  XOR U1435 ( .A(n26697), .B(n26867), .Z(n26701) );
  XOR U1436 ( .A(n25688), .B(n25858), .Z(n25692) );
  XOR U1437 ( .A(n24651), .B(n24821), .Z(n24655) );
  XOR U1438 ( .A(n23595), .B(n23765), .Z(n23599) );
  XOR U1439 ( .A(n22513), .B(n22683), .Z(n22517) );
  XOR U1440 ( .A(n21409), .B(n21579), .Z(n21413) );
  XOR U1441 ( .A(n20280), .B(n20450), .Z(n20284) );
  XOR U1442 ( .A(n19128), .B(n19298), .Z(n19132) );
  XOR U1443 ( .A(n10932), .B(n11109), .Z(n10936) );
  XOR U1444 ( .A(n8847), .B(n9114), .Z(n8851) );
  XOR U1445 ( .A(n6708), .B(n7065), .Z(n6712) );
  XOR U1446 ( .A(n4513), .B(n4960), .Z(n4517) );
  XOR U1447 ( .A(n3076), .B(n3517), .Z(n3080) );
  XOR U1448 ( .A(n5305), .B(n5658), .Z(n5309) );
  XOR U1449 ( .A(n7482), .B(n7743), .Z(n7486) );
  XOR U1450 ( .A(n45019), .B(n45183), .Z(n45023) );
  XOR U1451 ( .A(n44671), .B(n44835), .Z(n44675) );
  XOR U1452 ( .A(n4543), .B(n4954), .Z(n4547) );
  XOR U1453 ( .A(n6738), .B(n7059), .Z(n6742) );
  XOR U1454 ( .A(n8877), .B(n9108), .Z(n8881) );
  XOR U1455 ( .A(n14179), .B(n14338), .Z(n14183) );
  XOR U1456 ( .A(n10947), .B(n11106), .Z(n10951) );
  XOR U1457 ( .A(n7512), .B(n7737), .Z(n7516) );
  XOR U1458 ( .A(n5335), .B(n5652), .Z(n5339) );
  XOR U1459 ( .A(n3106), .B(n3511), .Z(n3110) );
  XOR U1460 ( .A(n44498), .B(n44650), .Z(n44502) );
  XOR U1461 ( .A(n44114), .B(n44266), .Z(n44118) );
  XOR U1462 ( .A(n43706), .B(n43858), .Z(n43710) );
  XOR U1463 ( .A(n43274), .B(n43426), .Z(n43278) );
  XOR U1464 ( .A(n42818), .B(n42970), .Z(n42822) );
  XOR U1465 ( .A(n42338), .B(n42490), .Z(n42342) );
  XOR U1466 ( .A(n41834), .B(n41986), .Z(n41838) );
  XOR U1467 ( .A(n41306), .B(n41458), .Z(n41310) );
  XOR U1468 ( .A(n40754), .B(n40906), .Z(n40758) );
  XOR U1469 ( .A(n40178), .B(n40330), .Z(n40182) );
  XOR U1470 ( .A(n39578), .B(n39730), .Z(n39582) );
  XOR U1471 ( .A(n38954), .B(n39106), .Z(n38958) );
  XOR U1472 ( .A(n38306), .B(n38458), .Z(n38310) );
  XOR U1473 ( .A(n37634), .B(n37786), .Z(n37638) );
  XOR U1474 ( .A(n36938), .B(n37090), .Z(n36942) );
  XOR U1475 ( .A(n36218), .B(n36370), .Z(n36222) );
  XOR U1476 ( .A(n35474), .B(n35626), .Z(n35478) );
  XOR U1477 ( .A(n34706), .B(n34858), .Z(n34710) );
  XOR U1478 ( .A(n33914), .B(n34066), .Z(n33918) );
  XOR U1479 ( .A(n33098), .B(n33250), .Z(n33102) );
  XOR U1480 ( .A(n32258), .B(n32410), .Z(n32262) );
  XOR U1481 ( .A(n31394), .B(n31546), .Z(n31398) );
  XOR U1482 ( .A(n30506), .B(n30658), .Z(n30510) );
  XOR U1483 ( .A(n29594), .B(n29746), .Z(n29598) );
  XOR U1484 ( .A(n28658), .B(n28810), .Z(n28662) );
  XOR U1485 ( .A(n27698), .B(n27850), .Z(n27702) );
  XOR U1486 ( .A(n26712), .B(n26864), .Z(n26716) );
  XOR U1487 ( .A(n25703), .B(n25855), .Z(n25707) );
  XOR U1488 ( .A(n24666), .B(n24818), .Z(n24670) );
  XOR U1489 ( .A(n23610), .B(n23762), .Z(n23614) );
  XOR U1490 ( .A(n22528), .B(n22680), .Z(n22532) );
  XOR U1491 ( .A(n21424), .B(n21576), .Z(n21428) );
  XOR U1492 ( .A(n20295), .B(n20447), .Z(n20299) );
  XOR U1493 ( .A(n19143), .B(n19295), .Z(n19147) );
  XOR U1494 ( .A(n8907), .B(n9102), .Z(n8911) );
  XOR U1495 ( .A(n6768), .B(n7053), .Z(n6772) );
  XOR U1496 ( .A(n4573), .B(n4948), .Z(n4577) );
  XOR U1497 ( .A(n3136), .B(n3505), .Z(n3140) );
  XOR U1498 ( .A(n5365), .B(n5646), .Z(n5369) );
  XOR U1499 ( .A(n7542), .B(n7731), .Z(n7546) );
  XOR U1500 ( .A(n45358), .B(n45504), .Z(n45362) );
  XOR U1501 ( .A(n45034), .B(n45180), .Z(n45038) );
  XOR U1502 ( .A(n4603), .B(n4942), .Z(n4607) );
  XOR U1503 ( .A(n6798), .B(n7047), .Z(n6802) );
  XOR U1504 ( .A(n8937), .B(n9096), .Z(n8941) );
  XOR U1505 ( .A(n15444), .B(n15585), .Z(n15448) );
  XOR U1506 ( .A(n11620), .B(n11761), .Z(n11624) );
  XOR U1507 ( .A(n7572), .B(n7725), .Z(n7576) );
  XOR U1508 ( .A(n5395), .B(n5640), .Z(n5399) );
  XOR U1509 ( .A(n3166), .B(n3499), .Z(n3170) );
  XOR U1510 ( .A(n44873), .B(n45007), .Z(n44877) );
  XOR U1511 ( .A(n44513), .B(n44647), .Z(n44517) );
  XOR U1512 ( .A(n44129), .B(n44263), .Z(n44133) );
  XOR U1513 ( .A(n43721), .B(n43855), .Z(n43725) );
  XOR U1514 ( .A(n43289), .B(n43423), .Z(n43293) );
  XOR U1515 ( .A(n42833), .B(n42967), .Z(n42837) );
  XOR U1516 ( .A(n42353), .B(n42487), .Z(n42357) );
  XOR U1517 ( .A(n41849), .B(n41983), .Z(n41853) );
  XOR U1518 ( .A(n41321), .B(n41455), .Z(n41325) );
  XOR U1519 ( .A(n40769), .B(n40903), .Z(n40773) );
  XOR U1520 ( .A(n40193), .B(n40327), .Z(n40197) );
  XOR U1521 ( .A(n39593), .B(n39727), .Z(n39597) );
  XOR U1522 ( .A(n38969), .B(n39103), .Z(n38973) );
  XOR U1523 ( .A(n38321), .B(n38455), .Z(n38325) );
  XOR U1524 ( .A(n37649), .B(n37783), .Z(n37653) );
  XOR U1525 ( .A(n36953), .B(n37087), .Z(n36957) );
  XOR U1526 ( .A(n36233), .B(n36367), .Z(n36237) );
  XOR U1527 ( .A(n35489), .B(n35623), .Z(n35493) );
  XOR U1528 ( .A(n34721), .B(n34855), .Z(n34725) );
  XOR U1529 ( .A(n33929), .B(n34063), .Z(n33933) );
  XOR U1530 ( .A(n33113), .B(n33247), .Z(n33117) );
  XOR U1531 ( .A(n32273), .B(n32407), .Z(n32277) );
  XOR U1532 ( .A(n31409), .B(n31543), .Z(n31413) );
  XOR U1533 ( .A(n30521), .B(n30655), .Z(n30525) );
  XOR U1534 ( .A(n29609), .B(n29743), .Z(n29613) );
  XOR U1535 ( .A(n28673), .B(n28807), .Z(n28677) );
  XOR U1536 ( .A(n27713), .B(n27847), .Z(n27717) );
  XOR U1537 ( .A(n26727), .B(n26861), .Z(n26731) );
  XOR U1538 ( .A(n25718), .B(n25852), .Z(n25722) );
  XOR U1539 ( .A(n24681), .B(n24815), .Z(n24685) );
  XOR U1540 ( .A(n23625), .B(n23759), .Z(n23629) );
  XOR U1541 ( .A(n22543), .B(n22677), .Z(n22547) );
  XOR U1542 ( .A(n21439), .B(n21573), .Z(n21443) );
  XOR U1543 ( .A(n20310), .B(n20444), .Z(n20314) );
  XOR U1544 ( .A(n19158), .B(n19292), .Z(n19162) );
  XOR U1545 ( .A(n16675), .B(n16810), .Z(n16679) );
  XOR U1546 ( .A(n9633), .B(n9768), .Z(n9637) );
  XOR U1547 ( .A(n6828), .B(n7041), .Z(n6832) );
  XOR U1548 ( .A(n4633), .B(n4936), .Z(n4637) );
  XOR U1549 ( .A(n3196), .B(n3493), .Z(n3200) );
  XOR U1550 ( .A(n5425), .B(n5634), .Z(n5429) );
  XOR U1551 ( .A(n45949), .B(n46077), .Z(n45953) );
  XOR U1552 ( .A(n45673), .B(n45801), .Z(n45677) );
  XOR U1553 ( .A(n4663), .B(n4930), .Z(n4667) );
  XOR U1554 ( .A(n6858), .B(n7035), .Z(n6862) );
  XOR U1555 ( .A(n8285), .B(n8408), .Z(n8289) );
  XOR U1556 ( .A(n5455), .B(n5628), .Z(n5459) );
  XOR U1557 ( .A(n3226), .B(n3487), .Z(n3230) );
  XOR U1558 ( .A(n45536), .B(n45652), .Z(n45540) );
  XOR U1559 ( .A(n45224), .B(n45340), .Z(n45228) );
  XOR U1560 ( .A(n44888), .B(n45004), .Z(n44892) );
  XOR U1561 ( .A(n44528), .B(n44644), .Z(n44532) );
  XOR U1562 ( .A(n44144), .B(n44260), .Z(n44148) );
  XOR U1563 ( .A(n43736), .B(n43852), .Z(n43740) );
  XOR U1564 ( .A(n43304), .B(n43420), .Z(n43308) );
  XOR U1565 ( .A(n42848), .B(n42964), .Z(n42852) );
  XOR U1566 ( .A(n42368), .B(n42484), .Z(n42372) );
  XOR U1567 ( .A(n41864), .B(n41980), .Z(n41868) );
  XOR U1568 ( .A(n41336), .B(n41452), .Z(n41340) );
  XOR U1569 ( .A(n40784), .B(n40900), .Z(n40788) );
  XOR U1570 ( .A(n40208), .B(n40324), .Z(n40212) );
  XOR U1571 ( .A(n39608), .B(n39724), .Z(n39612) );
  XOR U1572 ( .A(n38984), .B(n39100), .Z(n38988) );
  XOR U1573 ( .A(n38336), .B(n38452), .Z(n38340) );
  XOR U1574 ( .A(n37664), .B(n37780), .Z(n37668) );
  XOR U1575 ( .A(n36968), .B(n37084), .Z(n36972) );
  XOR U1576 ( .A(n36248), .B(n36364), .Z(n36252) );
  XOR U1577 ( .A(n35504), .B(n35620), .Z(n35508) );
  XOR U1578 ( .A(n34736), .B(n34852), .Z(n34740) );
  XOR U1579 ( .A(n33944), .B(n34060), .Z(n33948) );
  XOR U1580 ( .A(n33128), .B(n33244), .Z(n33132) );
  XOR U1581 ( .A(n32288), .B(n32404), .Z(n32292) );
  XOR U1582 ( .A(n31424), .B(n31540), .Z(n31428) );
  XOR U1583 ( .A(n30536), .B(n30652), .Z(n30540) );
  XOR U1584 ( .A(n29624), .B(n29740), .Z(n29628) );
  XOR U1585 ( .A(n28688), .B(n28804), .Z(n28692) );
  XOR U1586 ( .A(n27728), .B(n27844), .Z(n27732) );
  XOR U1587 ( .A(n26742), .B(n26858), .Z(n26746) );
  XOR U1588 ( .A(n25733), .B(n25849), .Z(n25737) );
  XOR U1589 ( .A(n24696), .B(n24812), .Z(n24700) );
  XOR U1590 ( .A(n23640), .B(n23756), .Z(n23644) );
  XOR U1591 ( .A(n22558), .B(n22674), .Z(n22562) );
  XOR U1592 ( .A(n21454), .B(n21570), .Z(n21458) );
  XOR U1593 ( .A(n20325), .B(n20441), .Z(n20329) );
  XOR U1594 ( .A(n19173), .B(n19289), .Z(n19177) );
  XOR U1595 ( .A(n11640), .B(n11757), .Z(n11644) );
  XOR U1596 ( .A(n6888), .B(n7029), .Z(n6892) );
  XOR U1597 ( .A(n4693), .B(n4924), .Z(n4697) );
  XOR U1598 ( .A(n3256), .B(n3481), .Z(n3260) );
  XOR U1599 ( .A(n5485), .B(n5622), .Z(n5489) );
  XOR U1600 ( .A(n46216), .B(n46326), .Z(n46220) );
  XOR U1601 ( .A(n45964), .B(n46074), .Z(n45968) );
  XOR U1602 ( .A(n14847), .B(n14958), .Z(n14851) );
  XOR U1603 ( .A(n4723), .B(n4918), .Z(n4727) );
  XOR U1604 ( .A(n13590), .B(n13695), .Z(n13594) );
  XOR U1605 ( .A(n3286), .B(n3475), .Z(n3290) );
  XOR U1606 ( .A(n45839), .B(n45937), .Z(n45843) );
  XOR U1607 ( .A(n45551), .B(n45649), .Z(n45555) );
  XOR U1608 ( .A(n45239), .B(n45337), .Z(n45243) );
  XOR U1609 ( .A(n44903), .B(n45001), .Z(n44907) );
  XOR U1610 ( .A(n44543), .B(n44641), .Z(n44547) );
  XOR U1611 ( .A(n44159), .B(n44257), .Z(n44163) );
  XOR U1612 ( .A(n43751), .B(n43849), .Z(n43755) );
  XOR U1613 ( .A(n43319), .B(n43417), .Z(n43323) );
  XOR U1614 ( .A(n42863), .B(n42961), .Z(n42867) );
  XOR U1615 ( .A(n42383), .B(n42481), .Z(n42387) );
  XOR U1616 ( .A(n41879), .B(n41977), .Z(n41883) );
  XOR U1617 ( .A(n41351), .B(n41449), .Z(n41355) );
  XOR U1618 ( .A(n40799), .B(n40897), .Z(n40803) );
  XOR U1619 ( .A(n40223), .B(n40321), .Z(n40227) );
  XOR U1620 ( .A(n39623), .B(n39721), .Z(n39627) );
  XOR U1621 ( .A(n38999), .B(n39097), .Z(n39003) );
  XOR U1622 ( .A(n38351), .B(n38449), .Z(n38355) );
  XOR U1623 ( .A(n37679), .B(n37777), .Z(n37683) );
  XOR U1624 ( .A(n36983), .B(n37081), .Z(n36987) );
  XOR U1625 ( .A(n36263), .B(n36361), .Z(n36267) );
  XOR U1626 ( .A(n35519), .B(n35617), .Z(n35523) );
  XOR U1627 ( .A(n34751), .B(n34849), .Z(n34755) );
  XOR U1628 ( .A(n33959), .B(n34057), .Z(n33963) );
  XOR U1629 ( .A(n33143), .B(n33241), .Z(n33147) );
  XOR U1630 ( .A(n32303), .B(n32401), .Z(n32307) );
  XOR U1631 ( .A(n31439), .B(n31537), .Z(n31443) );
  XOR U1632 ( .A(n30551), .B(n30649), .Z(n30555) );
  XOR U1633 ( .A(n29639), .B(n29737), .Z(n29643) );
  XOR U1634 ( .A(n28703), .B(n28801), .Z(n28707) );
  XOR U1635 ( .A(n27743), .B(n27841), .Z(n27747) );
  XOR U1636 ( .A(n26757), .B(n26855), .Z(n26761) );
  XOR U1637 ( .A(n25748), .B(n25846), .Z(n25752) );
  XOR U1638 ( .A(n24711), .B(n24809), .Z(n24715) );
  XOR U1639 ( .A(n23655), .B(n23753), .Z(n23659) );
  XOR U1640 ( .A(n22573), .B(n22671), .Z(n22577) );
  XOR U1641 ( .A(n21469), .B(n21567), .Z(n21473) );
  XOR U1642 ( .A(n20340), .B(n20438), .Z(n20344) );
  XOR U1643 ( .A(n19188), .B(n19286), .Z(n19192) );
  XOR U1644 ( .A(n4753), .B(n4912), .Z(n4757) );
  XOR U1645 ( .A(n3316), .B(n3469), .Z(n3320) );
  XOR U1646 ( .A(n46663), .B(n46755), .Z(n46667) );
  XOR U1647 ( .A(n46459), .B(n46551), .Z(n46463) );
  XOR U1648 ( .A(n16710), .B(n16803), .Z(n16714) );
  XOR U1649 ( .A(n6928), .B(n7021), .Z(n6932) );
  XOR U1650 ( .A(n5520), .B(n5615), .Z(n5524) );
  XOR U1651 ( .A(n4783), .B(n4906), .Z(n4787) );
  XOR U1652 ( .A(n3346), .B(n3463), .Z(n3350) );
  XOR U1653 ( .A(n46358), .B(n46438), .Z(n46362) );
  XOR U1654 ( .A(n46118), .B(n46198), .Z(n46122) );
  XOR U1655 ( .A(n45854), .B(n45934), .Z(n45858) );
  XOR U1656 ( .A(n45566), .B(n45646), .Z(n45570) );
  XOR U1657 ( .A(n45254), .B(n45334), .Z(n45258) );
  XOR U1658 ( .A(n44918), .B(n44998), .Z(n44922) );
  XOR U1659 ( .A(n44558), .B(n44638), .Z(n44562) );
  XOR U1660 ( .A(n44174), .B(n44254), .Z(n44178) );
  XOR U1661 ( .A(n43766), .B(n43846), .Z(n43770) );
  XOR U1662 ( .A(n43334), .B(n43414), .Z(n43338) );
  XOR U1663 ( .A(n42878), .B(n42958), .Z(n42882) );
  XOR U1664 ( .A(n42398), .B(n42478), .Z(n42402) );
  XOR U1665 ( .A(n41894), .B(n41974), .Z(n41898) );
  XOR U1666 ( .A(n41366), .B(n41446), .Z(n41370) );
  XOR U1667 ( .A(n40814), .B(n40894), .Z(n40818) );
  XOR U1668 ( .A(n40238), .B(n40318), .Z(n40242) );
  XOR U1669 ( .A(n39638), .B(n39718), .Z(n39642) );
  XOR U1670 ( .A(n39014), .B(n39094), .Z(n39018) );
  XOR U1671 ( .A(n38366), .B(n38446), .Z(n38370) );
  XOR U1672 ( .A(n37694), .B(n37774), .Z(n37698) );
  XOR U1673 ( .A(n36998), .B(n37078), .Z(n37002) );
  XOR U1674 ( .A(n36278), .B(n36358), .Z(n36282) );
  XOR U1675 ( .A(n35534), .B(n35614), .Z(n35538) );
  XOR U1676 ( .A(n34766), .B(n34846), .Z(n34770) );
  XOR U1677 ( .A(n33974), .B(n34054), .Z(n33978) );
  XOR U1678 ( .A(n33158), .B(n33238), .Z(n33162) );
  XOR U1679 ( .A(n32318), .B(n32398), .Z(n32322) );
  XOR U1680 ( .A(n31454), .B(n31534), .Z(n31458) );
  XOR U1681 ( .A(n30566), .B(n30646), .Z(n30570) );
  XOR U1682 ( .A(n29654), .B(n29734), .Z(n29658) );
  XOR U1683 ( .A(n28718), .B(n28798), .Z(n28722) );
  XOR U1684 ( .A(n27758), .B(n27838), .Z(n27762) );
  XOR U1685 ( .A(n26772), .B(n26852), .Z(n26776) );
  XOR U1686 ( .A(n25763), .B(n25843), .Z(n25767) );
  XOR U1687 ( .A(n24726), .B(n24806), .Z(n24730) );
  XOR U1688 ( .A(n23670), .B(n23750), .Z(n23674) );
  XOR U1689 ( .A(n22588), .B(n22668), .Z(n22592) );
  XOR U1690 ( .A(n21484), .B(n21564), .Z(n21488) );
  XOR U1691 ( .A(n20355), .B(n20435), .Z(n20359) );
  XOR U1692 ( .A(n19203), .B(n19283), .Z(n19207) );
  XOR U1693 ( .A(n4813), .B(n4900), .Z(n4817) );
  XOR U1694 ( .A(n3376), .B(n3457), .Z(n3380) );
  XOR U1695 ( .A(n46858), .B(n46932), .Z(n46862) );
  XOR U1696 ( .A(n46678), .B(n46752), .Z(n46682) );
  XOR U1697 ( .A(n5540), .B(n5611), .Z(n5544) );
  XOR U1698 ( .A(n46589), .B(n46651), .Z(n46593) );
  XOR U1699 ( .A(n46373), .B(n46435), .Z(n46377) );
  XOR U1700 ( .A(n46133), .B(n46195), .Z(n46137) );
  XOR U1701 ( .A(n45869), .B(n45931), .Z(n45873) );
  XOR U1702 ( .A(n45581), .B(n45643), .Z(n45585) );
  XOR U1703 ( .A(n45269), .B(n45331), .Z(n45273) );
  XOR U1704 ( .A(n44933), .B(n44995), .Z(n44937) );
  XOR U1705 ( .A(n44573), .B(n44635), .Z(n44577) );
  XOR U1706 ( .A(n44189), .B(n44251), .Z(n44193) );
  XOR U1707 ( .A(n43781), .B(n43843), .Z(n43785) );
  XOR U1708 ( .A(n43349), .B(n43411), .Z(n43353) );
  XOR U1709 ( .A(n42893), .B(n42955), .Z(n42897) );
  XOR U1710 ( .A(n42413), .B(n42475), .Z(n42417) );
  XOR U1711 ( .A(n41909), .B(n41971), .Z(n41913) );
  XOR U1712 ( .A(n41381), .B(n41443), .Z(n41385) );
  XOR U1713 ( .A(n40829), .B(n40891), .Z(n40833) );
  XOR U1714 ( .A(n40253), .B(n40315), .Z(n40257) );
  XOR U1715 ( .A(n39653), .B(n39715), .Z(n39657) );
  XOR U1716 ( .A(n39029), .B(n39091), .Z(n39033) );
  XOR U1717 ( .A(n38381), .B(n38443), .Z(n38385) );
  XOR U1718 ( .A(n37709), .B(n37771), .Z(n37713) );
  XOR U1719 ( .A(n37013), .B(n37075), .Z(n37017) );
  XOR U1720 ( .A(n36293), .B(n36355), .Z(n36297) );
  XOR U1721 ( .A(n35549), .B(n35611), .Z(n35553) );
  XOR U1722 ( .A(n34781), .B(n34843), .Z(n34785) );
  XOR U1723 ( .A(n33989), .B(n34051), .Z(n33993) );
  XOR U1724 ( .A(n33173), .B(n33235), .Z(n33177) );
  XOR U1725 ( .A(n32333), .B(n32395), .Z(n32337) );
  XOR U1726 ( .A(n31469), .B(n31531), .Z(n31473) );
  XOR U1727 ( .A(n30581), .B(n30643), .Z(n30585) );
  XOR U1728 ( .A(n29669), .B(n29731), .Z(n29673) );
  XOR U1729 ( .A(n28733), .B(n28795), .Z(n28737) );
  XOR U1730 ( .A(n27773), .B(n27835), .Z(n27777) );
  XOR U1731 ( .A(n26787), .B(n26849), .Z(n26791) );
  XOR U1732 ( .A(n25778), .B(n25840), .Z(n25782) );
  XOR U1733 ( .A(n24741), .B(n24803), .Z(n24745) );
  XOR U1734 ( .A(n23685), .B(n23747), .Z(n23689) );
  XOR U1735 ( .A(n22603), .B(n22665), .Z(n22607) );
  XOR U1736 ( .A(n21499), .B(n21561), .Z(n21503) );
  XOR U1737 ( .A(n20370), .B(n20432), .Z(n20374) );
  XOR U1738 ( .A(n19218), .B(n19280), .Z(n19222) );
  XOR U1739 ( .A(n15509), .B(n15572), .Z(n15513) );
  XOR U1740 ( .A(n4115), .B(n4178), .Z(n4119) );
  XOR U1741 ( .A(n47029), .B(n47085), .Z(n47033) );
  XOR U1742 ( .A(n3396), .B(n3453), .Z(n3400) );
  XOR U1743 ( .A(n47278), .B(n47322), .Z(n47282) );
  XOR U1744 ( .A(n46964), .B(n47008), .Z(n46968) );
  XOR U1745 ( .A(n46796), .B(n46840), .Z(n46800) );
  XOR U1746 ( .A(n46604), .B(n46648), .Z(n46608) );
  XOR U1747 ( .A(n46388), .B(n46432), .Z(n46392) );
  XOR U1748 ( .A(n46148), .B(n46192), .Z(n46152) );
  XOR U1749 ( .A(n45884), .B(n45928), .Z(n45888) );
  XOR U1750 ( .A(n45596), .B(n45640), .Z(n45600) );
  XOR U1751 ( .A(n45284), .B(n45328), .Z(n45288) );
  XOR U1752 ( .A(n44948), .B(n44992), .Z(n44952) );
  XOR U1753 ( .A(n44588), .B(n44632), .Z(n44592) );
  XOR U1754 ( .A(n44204), .B(n44248), .Z(n44208) );
  XOR U1755 ( .A(n43796), .B(n43840), .Z(n43800) );
  XOR U1756 ( .A(n43364), .B(n43408), .Z(n43368) );
  XOR U1757 ( .A(n42908), .B(n42952), .Z(n42912) );
  XOR U1758 ( .A(n42428), .B(n42472), .Z(n42432) );
  XOR U1759 ( .A(n41924), .B(n41968), .Z(n41928) );
  XOR U1760 ( .A(n41396), .B(n41440), .Z(n41400) );
  XOR U1761 ( .A(n40844), .B(n40888), .Z(n40848) );
  XOR U1762 ( .A(n40268), .B(n40312), .Z(n40272) );
  XOR U1763 ( .A(n39668), .B(n39712), .Z(n39672) );
  XOR U1764 ( .A(n39044), .B(n39088), .Z(n39048) );
  XOR U1765 ( .A(n38396), .B(n38440), .Z(n38400) );
  XOR U1766 ( .A(n37724), .B(n37768), .Z(n37728) );
  XOR U1767 ( .A(n37028), .B(n37072), .Z(n37032) );
  XOR U1768 ( .A(n36308), .B(n36352), .Z(n36312) );
  XOR U1769 ( .A(n35564), .B(n35608), .Z(n35568) );
  XOR U1770 ( .A(n34796), .B(n34840), .Z(n34800) );
  XOR U1771 ( .A(n34004), .B(n34048), .Z(n34008) );
  XOR U1772 ( .A(n33188), .B(n33232), .Z(n33192) );
  XOR U1773 ( .A(n32348), .B(n32392), .Z(n32352) );
  XOR U1774 ( .A(n31484), .B(n31528), .Z(n31488) );
  XOR U1775 ( .A(n30596), .B(n30640), .Z(n30600) );
  XOR U1776 ( .A(n29684), .B(n29728), .Z(n29688) );
  XOR U1777 ( .A(n28748), .B(n28792), .Z(n28752) );
  XOR U1778 ( .A(n27788), .B(n27832), .Z(n27792) );
  XOR U1779 ( .A(n26802), .B(n26846), .Z(n26806) );
  XOR U1780 ( .A(n25793), .B(n25837), .Z(n25797) );
  XOR U1781 ( .A(n24756), .B(n24800), .Z(n24760) );
  XOR U1782 ( .A(n23700), .B(n23744), .Z(n23704) );
  XOR U1783 ( .A(n22618), .B(n22662), .Z(n22622) );
  XOR U1784 ( .A(n21514), .B(n21558), .Z(n21518) );
  XOR U1785 ( .A(n20385), .B(n20429), .Z(n20389) );
  XOR U1786 ( .A(n19233), .B(n19277), .Z(n19237) );
  XOR U1787 ( .A(n16750), .B(n16795), .Z(n16754) );
  XOR U1788 ( .A(n47176), .B(n47213), .Z(n47180) );
  XNOR U1789 ( .A(n47182), .B(n47116), .Z(n47118) );
  XOR U1790 ( .A(n47410), .B(n47436), .Z(n47414) );
  XOR U1791 ( .A(n47338), .B(n47364), .Z(n47342) );
  XOR U1792 ( .A(n46979), .B(n47005), .Z(n46983) );
  XOR U1793 ( .A(n46811), .B(n46837), .Z(n46815) );
  XOR U1794 ( .A(n46619), .B(n46645), .Z(n46623) );
  XOR U1795 ( .A(n46403), .B(n46429), .Z(n46407) );
  XOR U1796 ( .A(n46163), .B(n46189), .Z(n46167) );
  XOR U1797 ( .A(n45899), .B(n45925), .Z(n45903) );
  XOR U1798 ( .A(n45611), .B(n45637), .Z(n45615) );
  XOR U1799 ( .A(n45299), .B(n45325), .Z(n45303) );
  XOR U1800 ( .A(n44963), .B(n44989), .Z(n44967) );
  XOR U1801 ( .A(n44603), .B(n44629), .Z(n44607) );
  XOR U1802 ( .A(n44219), .B(n44245), .Z(n44223) );
  XOR U1803 ( .A(n43811), .B(n43837), .Z(n43815) );
  XOR U1804 ( .A(n43379), .B(n43405), .Z(n43383) );
  XOR U1805 ( .A(n42923), .B(n42949), .Z(n42927) );
  XOR U1806 ( .A(n42443), .B(n42469), .Z(n42447) );
  XOR U1807 ( .A(n41939), .B(n41965), .Z(n41943) );
  XOR U1808 ( .A(n41411), .B(n41437), .Z(n41415) );
  XOR U1809 ( .A(n40859), .B(n40885), .Z(n40863) );
  XOR U1810 ( .A(n40283), .B(n40309), .Z(n40287) );
  XOR U1811 ( .A(n39683), .B(n39709), .Z(n39687) );
  XOR U1812 ( .A(n39059), .B(n39085), .Z(n39063) );
  XOR U1813 ( .A(n38411), .B(n38437), .Z(n38415) );
  XOR U1814 ( .A(n37739), .B(n37765), .Z(n37743) );
  XOR U1815 ( .A(n37043), .B(n37069), .Z(n37047) );
  XOR U1816 ( .A(n36323), .B(n36349), .Z(n36327) );
  XOR U1817 ( .A(n35579), .B(n35605), .Z(n35583) );
  XOR U1818 ( .A(n34811), .B(n34837), .Z(n34815) );
  XOR U1819 ( .A(n34019), .B(n34045), .Z(n34023) );
  XOR U1820 ( .A(n33203), .B(n33229), .Z(n33207) );
  XOR U1821 ( .A(n32363), .B(n32389), .Z(n32367) );
  XOR U1822 ( .A(n31499), .B(n31525), .Z(n31503) );
  XOR U1823 ( .A(n30611), .B(n30637), .Z(n30615) );
  XOR U1824 ( .A(n29699), .B(n29725), .Z(n29703) );
  XOR U1825 ( .A(n28763), .B(n28789), .Z(n28767) );
  XOR U1826 ( .A(n27803), .B(n27829), .Z(n27807) );
  XOR U1827 ( .A(n26817), .B(n26843), .Z(n26821) );
  XOR U1828 ( .A(n25808), .B(n25834), .Z(n25812) );
  XOR U1829 ( .A(n24771), .B(n24797), .Z(n24775) );
  XOR U1830 ( .A(n23715), .B(n23741), .Z(n23719) );
  XOR U1831 ( .A(n22633), .B(n22659), .Z(n22637) );
  XOR U1832 ( .A(n21529), .B(n21555), .Z(n21533) );
  XOR U1833 ( .A(n20400), .B(n20426), .Z(n20404) );
  XOR U1834 ( .A(n19248), .B(n19274), .Z(n19252) );
  XOR U1835 ( .A(n47298), .B(n47318), .Z(n47302) );
  XOR U1836 ( .A(n47191), .B(n47210), .Z(n47195) );
  XOR U1837 ( .A(n27911), .B(n28387), .Z(n27915) );
  XNOR U1838 ( .A(n27917), .B(n27431), .Z(n27433) );
  XNOR U1839 ( .A(n27922), .B(n27436), .Z(n27438) );
  XOR U1840 ( .A(n26427), .B(n26923), .Z(n26431) );
  XOR U1841 ( .A(n28874), .B(n29332), .Z(n28878) );
  XOR U1842 ( .A(n27931), .B(n28383), .Z(n27935) );
  XOR U1843 ( .A(n27448), .B(n27900), .Z(n27452) );
  XOR U1844 ( .A(n26442), .B(n26920), .Z(n26446) );
  XOR U1845 ( .A(n25413), .B(n25914), .Z(n25417) );
  XOR U1846 ( .A(n25956), .B(n26414), .Z(n25960) );
  XNOR U1847 ( .A(n24889), .B(n24364), .Z(n24366) );
  XOR U1848 ( .A(n30266), .B(n30706), .Z(n30270) );
  XOR U1849 ( .A(n29354), .B(n29794), .Z(n29358) );
  XOR U1850 ( .A(n25463), .B(n25904), .Z(n25467) );
  XNOR U1851 ( .A(n29824), .B(n29362), .Z(n29364) );
  XOR U1852 ( .A(n28423), .B(n28857), .Z(n28427) );
  XOR U1853 ( .A(n27463), .B(n27897), .Z(n27467) );
  XNOR U1854 ( .A(n26980), .B(n26480), .Z(n26482) );
  XNOR U1855 ( .A(n26473), .B(n25969), .Z(n25971) );
  XOR U1856 ( .A(n25428), .B(n25911), .Z(n25432) );
  XOR U1857 ( .A(n24396), .B(n24875), .Z(n24400) );
  XOR U1858 ( .A(n24376), .B(n24879), .Z(n24380) );
  XOR U1859 ( .A(n24953), .B(n25389), .Z(n24957) );
  XOR U1860 ( .A(n31604), .B(n32026), .Z(n31608) );
  XOR U1861 ( .A(n30728), .B(n31150), .Z(n30732) );
  XOR U1862 ( .A(n25478), .B(n25900), .Z(n25482) );
  XOR U1863 ( .A(n23325), .B(n23819), .Z(n23329) );
  XOR U1864 ( .A(n23305), .B(n23823), .Z(n23309) );
  XOR U1865 ( .A(n23891), .B(n24343), .Z(n23895) );
  XOR U1866 ( .A(n30286), .B(n30702), .Z(n30290) );
  XOR U1867 ( .A(n29374), .B(n29790), .Z(n29378) );
  XOR U1868 ( .A(n28438), .B(n28854), .Z(n28442) );
  XOR U1869 ( .A(n27478), .B(n27894), .Z(n27482) );
  XOR U1870 ( .A(n26492), .B(n26908), .Z(n26496) );
  XNOR U1871 ( .A(n24934), .B(n24409), .Z(n24411) );
  XOR U1872 ( .A(n22208), .B(n22745), .Z(n22212) );
  XOR U1873 ( .A(n24968), .B(n25385), .Z(n24972) );
  XOR U1874 ( .A(n32888), .B(n33292), .Z(n32892) );
  XOR U1875 ( .A(n32048), .B(n32452), .Z(n32052) );
  XOR U1876 ( .A(n21679), .B(n22191), .Z(n21683) );
  XOR U1877 ( .A(n22772), .B(n23285), .Z(n22776) );
  XOR U1878 ( .A(n23906), .B(n24340), .Z(n23910) );
  XOR U1879 ( .A(n22817), .B(n23276), .Z(n22821) );
  XOR U1880 ( .A(n21704), .B(n22186), .Z(n21708) );
  XNOR U1881 ( .A(n32482), .B(n32056), .Z(n32058) );
  XOR U1882 ( .A(n31189), .B(n31587), .Z(n31193) );
  XOR U1883 ( .A(n30301), .B(n30699), .Z(n30305) );
  XOR U1884 ( .A(n29389), .B(n29787), .Z(n29393) );
  XOR U1885 ( .A(n28453), .B(n28851), .Z(n28457) );
  XOR U1886 ( .A(n27493), .B(n27891), .Z(n27497) );
  XOR U1887 ( .A(n26507), .B(n26905), .Z(n26511) );
  XOR U1888 ( .A(n25498), .B(n25896), .Z(n25502) );
  XOR U1889 ( .A(n23931), .B(n24335), .Z(n23935) );
  XOR U1890 ( .A(n22842), .B(n23271), .Z(n22846) );
  XOR U1891 ( .A(n23345), .B(n23815), .Z(n23349) );
  XOR U1892 ( .A(n21664), .B(n22194), .Z(n21668) );
  XOR U1893 ( .A(n20527), .B(n21082), .Z(n20531) );
  XOR U1894 ( .A(n22248), .B(n22737), .Z(n22252) );
  XOR U1895 ( .A(n34118), .B(n34504), .Z(n34122) );
  XOR U1896 ( .A(n33314), .B(n33700), .Z(n33318) );
  XNOR U1897 ( .A(n25000), .B(n24474), .Z(n24476) );
  XOR U1898 ( .A(n20557), .B(n21076), .Z(n20561) );
  XOR U1899 ( .A(n21719), .B(n22183), .Z(n21723) );
  XNOR U1900 ( .A(n23421), .B(n22880), .Z(n22882) );
  XOR U1901 ( .A(n22323), .B(n22722), .Z(n22327) );
  XOR U1902 ( .A(n32908), .B(n33288), .Z(n32912) );
  XOR U1903 ( .A(n32068), .B(n32448), .Z(n32072) );
  XOR U1904 ( .A(n31204), .B(n31584), .Z(n31208) );
  XOR U1905 ( .A(n30316), .B(n30696), .Z(n30320) );
  XOR U1906 ( .A(n29404), .B(n29784), .Z(n29408) );
  XOR U1907 ( .A(n28468), .B(n28848), .Z(n28472) );
  XOR U1908 ( .A(n27508), .B(n27888), .Z(n27512) );
  XOR U1909 ( .A(n26522), .B(n26902), .Z(n26526) );
  XOR U1910 ( .A(n25513), .B(n25893), .Z(n25517) );
  XOR U1911 ( .A(n23951), .B(n24331), .Z(n23955) );
  XNOR U1912 ( .A(n23401), .B(n22860), .Z(n22862) );
  XOR U1913 ( .A(n22303), .B(n22726), .Z(n22307) );
  XOR U1914 ( .A(n20542), .B(n21079), .Z(n20546) );
  XOR U1915 ( .A(n19382), .B(n19942), .Z(n19386) );
  XOR U1916 ( .A(n22283), .B(n22730), .Z(n22287) );
  XOR U1917 ( .A(n20587), .B(n21070), .Z(n20591) );
  XNOR U1918 ( .A(n23426), .B(n22885), .Z(n22887) );
  XOR U1919 ( .A(n21184), .B(n21624), .Z(n21188) );
  XNOR U1920 ( .A(n19966), .B(n19390), .Z(n19392) );
  XOR U1921 ( .A(n18843), .B(n19355), .Z(n18847) );
  XOR U1922 ( .A(n35294), .B(n35662), .Z(n35298) );
  XOR U1923 ( .A(n34526), .B(n34894), .Z(n34530) );
  XNOR U1924 ( .A(n23967), .B(n23433), .Z(n23435) );
  XOR U1925 ( .A(n20572), .B(n21073), .Z(n20576) );
  XOR U1926 ( .A(n18119), .B(n18771), .Z(n18123) );
  XOR U1927 ( .A(n19412), .B(n19936), .Z(n19416) );
  XOR U1928 ( .A(n21214), .B(n21618), .Z(n21218) );
  XNOR U1929 ( .A(n34924), .B(n34534), .Z(n34536) );
  XOR U1930 ( .A(n33739), .B(n34101), .Z(n33743) );
  XOR U1931 ( .A(n32923), .B(n33285), .Z(n32927) );
  XOR U1932 ( .A(n32083), .B(n32445), .Z(n32087) );
  XOR U1933 ( .A(n31219), .B(n31581), .Z(n31223) );
  XOR U1934 ( .A(n30331), .B(n30693), .Z(n30335) );
  XOR U1935 ( .A(n29419), .B(n29781), .Z(n29423) );
  XOR U1936 ( .A(n28483), .B(n28845), .Z(n28487) );
  XOR U1937 ( .A(n27523), .B(n27885), .Z(n27527) );
  XOR U1938 ( .A(n26537), .B(n26899), .Z(n26541) );
  XOR U1939 ( .A(n25528), .B(n25890), .Z(n25532) );
  XOR U1940 ( .A(n24491), .B(n24853), .Z(n24495) );
  XNOR U1941 ( .A(n22903), .B(n22356), .Z(n22358) );
  XOR U1942 ( .A(n21759), .B(n22175), .Z(n21763) );
  XNOR U1943 ( .A(n20041), .B(n19465), .Z(n19467) );
  XOR U1944 ( .A(n18873), .B(n19349), .Z(n18877) );
  XNOR U1945 ( .A(n19996), .B(n19420), .Z(n19422) );
  XOR U1946 ( .A(n20602), .B(n21067), .Z(n20606) );
  XOR U1947 ( .A(n19442), .B(n19930), .Z(n19446) );
  XOR U1948 ( .A(n22343), .B(n22718), .Z(n22347) );
  XNOR U1949 ( .A(n21780), .B(n21222), .Z(n21224) );
  XOR U1950 ( .A(n20070), .B(n20492), .Z(n20074) );
  XOR U1951 ( .A(n21244), .B(n21612), .Z(n21248) );
  XOR U1952 ( .A(n20627), .B(n21062), .Z(n20631) );
  XOR U1953 ( .A(n17507), .B(n18086), .Z(n17511) );
  XNOR U1954 ( .A(n20026), .B(n19450), .Z(n19452) );
  XOR U1955 ( .A(n36416), .B(n36766), .Z(n36420) );
  XOR U1956 ( .A(n35684), .B(n36034), .Z(n35688) );
  XNOR U1957 ( .A(n22369), .B(n21817), .Z(n21819) );
  XNOR U1958 ( .A(n21810), .B(n21252), .Z(n21254) );
  XOR U1959 ( .A(n20100), .B(n20486), .Z(n20104) );
  XOR U1960 ( .A(n16310), .B(n16883), .Z(n16314) );
  XOR U1961 ( .A(n16949), .B(n17480), .Z(n16953) );
  XNOR U1962 ( .A(n36064), .B(n35692), .Z(n35694) );
  XOR U1963 ( .A(n34933), .B(n35277), .Z(n34937) );
  XOR U1964 ( .A(n34153), .B(n34497), .Z(n34157) );
  XOR U1965 ( .A(n33349), .B(n33693), .Z(n33353) );
  XOR U1966 ( .A(n32521), .B(n32865), .Z(n32525) );
  XOR U1967 ( .A(n31669), .B(n32013), .Z(n31673) );
  XOR U1968 ( .A(n30793), .B(n31137), .Z(n30797) );
  XOR U1969 ( .A(n29893), .B(n30237), .Z(n29897) );
  XOR U1970 ( .A(n28969), .B(n29313), .Z(n28973) );
  XOR U1971 ( .A(n28021), .B(n28365), .Z(n28025) );
  XOR U1972 ( .A(n27049), .B(n27393), .Z(n27053) );
  XOR U1973 ( .A(n26051), .B(n26395), .Z(n26055) );
  XOR U1974 ( .A(n25029), .B(n25373), .Z(n25033) );
  XOR U1975 ( .A(n23981), .B(n24325), .Z(n23985) );
  XOR U1976 ( .A(n22912), .B(n23256), .Z(n22916) );
  XOR U1977 ( .A(n18933), .B(n19337), .Z(n18937) );
  XOR U1978 ( .A(n18888), .B(n19346), .Z(n18892) );
  XOR U1979 ( .A(n17537), .B(n18080), .Z(n17541) );
  XOR U1980 ( .A(n20662), .B(n21055), .Z(n20666) );
  XOR U1981 ( .A(n20130), .B(n20480), .Z(n20134) );
  XOR U1982 ( .A(n19482), .B(n19922), .Z(n19486) );
  XOR U1983 ( .A(n16979), .B(n17474), .Z(n16983) );
  XOR U1984 ( .A(n15680), .B(n16277), .Z(n15684) );
  XOR U1985 ( .A(n19507), .B(n19917), .Z(n19511) );
  XOR U1986 ( .A(n18963), .B(n19331), .Z(n18967) );
  XOR U1987 ( .A(n37484), .B(n37816), .Z(n37488) );
  XOR U1988 ( .A(n36788), .B(n37120), .Z(n36792) );
  XOR U1989 ( .A(n20712), .B(n21044), .Z(n20716) );
  XOR U1990 ( .A(n20692), .B(n21049), .Z(n20696) );
  XOR U1991 ( .A(n14447), .B(n15038), .Z(n14451) );
  XOR U1992 ( .A(n16964), .B(n17477), .Z(n16968) );
  XOR U1993 ( .A(n15104), .B(n15653), .Z(n15108) );
  XOR U1994 ( .A(n18219), .B(n18731), .Z(n18223) );
  XOR U1995 ( .A(n17009), .B(n17468), .Z(n17013) );
  XOR U1996 ( .A(n36436), .B(n36762), .Z(n36440) );
  XOR U1997 ( .A(n35704), .B(n36030), .Z(n35708) );
  XOR U1998 ( .A(n34948), .B(n35274), .Z(n34952) );
  XOR U1999 ( .A(n34168), .B(n34494), .Z(n34172) );
  XOR U2000 ( .A(n33364), .B(n33690), .Z(n33368) );
  XOR U2001 ( .A(n32536), .B(n32862), .Z(n32540) );
  XOR U2002 ( .A(n31684), .B(n32010), .Z(n31688) );
  XOR U2003 ( .A(n30808), .B(n31134), .Z(n30812) );
  XOR U2004 ( .A(n29908), .B(n30234), .Z(n29912) );
  XOR U2005 ( .A(n28984), .B(n29310), .Z(n28988) );
  XOR U2006 ( .A(n28036), .B(n28362), .Z(n28040) );
  XOR U2007 ( .A(n27064), .B(n27390), .Z(n27068) );
  XOR U2008 ( .A(n26066), .B(n26392), .Z(n26070) );
  XOR U2009 ( .A(n25044), .B(n25370), .Z(n25048) );
  XOR U2010 ( .A(n23996), .B(n24322), .Z(n24000) );
  XOR U2011 ( .A(n22927), .B(n23253), .Z(n22931) );
  XOR U2012 ( .A(n21834), .B(n22160), .Z(n21838) );
  XOR U2013 ( .A(n19537), .B(n19911), .Z(n19541) );
  XOR U2014 ( .A(n15710), .B(n16271), .Z(n15714) );
  XOR U2015 ( .A(n18998), .B(n19324), .Z(n19002) );
  XOR U2016 ( .A(n18249), .B(n18719), .Z(n18253) );
  XOR U2017 ( .A(n17039), .B(n17462), .Z(n17043) );
  XOR U2018 ( .A(n17602), .B(n18067), .Z(n17606) );
  XOR U2019 ( .A(n16380), .B(n16869), .Z(n16384) );
  XOR U2020 ( .A(n15134), .B(n15647), .Z(n15138) );
  XOR U2021 ( .A(n13799), .B(n14414), .Z(n13803) );
  XOR U2022 ( .A(n20150), .B(n20476), .Z(n20154) );
  XOR U2023 ( .A(n19567), .B(n19905), .Z(n19571) );
  XOR U2024 ( .A(n38498), .B(n38812), .Z(n38502) );
  XOR U2025 ( .A(n37838), .B(n38152), .Z(n37842) );
  XOR U2026 ( .A(n12530), .B(n13139), .Z(n12534) );
  XOR U2027 ( .A(n15119), .B(n15650), .Z(n15123) );
  XOR U2028 ( .A(n13205), .B(n13772), .Z(n13209) );
  XOR U2029 ( .A(n17632), .B(n18061), .Z(n17636) );
  XOR U2030 ( .A(n16410), .B(n16863), .Z(n16414) );
  XOR U2031 ( .A(n15164), .B(n15641), .Z(n15168) );
  XOR U2032 ( .A(n18279), .B(n18707), .Z(n18283) );
  XOR U2033 ( .A(n17069), .B(n17456), .Z(n17073) );
  XNOR U2034 ( .A(n38182), .B(n37846), .Z(n37848) );
  XOR U2035 ( .A(n37159), .B(n37467), .Z(n37163) );
  XOR U2036 ( .A(n36451), .B(n36759), .Z(n36455) );
  XOR U2037 ( .A(n35719), .B(n36027), .Z(n35723) );
  XOR U2038 ( .A(n34963), .B(n35271), .Z(n34967) );
  XOR U2039 ( .A(n34183), .B(n34491), .Z(n34187) );
  XOR U2040 ( .A(n33379), .B(n33687), .Z(n33383) );
  XOR U2041 ( .A(n32551), .B(n32859), .Z(n32555) );
  XOR U2042 ( .A(n31699), .B(n32007), .Z(n31703) );
  XOR U2043 ( .A(n30823), .B(n31131), .Z(n30827) );
  XOR U2044 ( .A(n29923), .B(n30231), .Z(n29927) );
  XOR U2045 ( .A(n28999), .B(n29307), .Z(n29003) );
  XOR U2046 ( .A(n28051), .B(n28359), .Z(n28055) );
  XOR U2047 ( .A(n27079), .B(n27387), .Z(n27083) );
  XOR U2048 ( .A(n26081), .B(n26389), .Z(n26085) );
  XOR U2049 ( .A(n25059), .B(n25367), .Z(n25063) );
  XOR U2050 ( .A(n24011), .B(n24319), .Z(n24015) );
  XOR U2051 ( .A(n22942), .B(n23250), .Z(n22946) );
  XOR U2052 ( .A(n21849), .B(n22157), .Z(n21853) );
  XOR U2053 ( .A(n20732), .B(n21040), .Z(n20736) );
  XNOR U2054 ( .A(n20171), .B(n19595), .Z(n19597) );
  XOR U2055 ( .A(n13829), .B(n14408), .Z(n13833) );
  XOR U2056 ( .A(n18309), .B(n18695), .Z(n18313) );
  XOR U2057 ( .A(n17099), .B(n17450), .Z(n17103) );
  XOR U2058 ( .A(n17662), .B(n18055), .Z(n17666) );
  XOR U2059 ( .A(n16440), .B(n16857), .Z(n16444) );
  XOR U2060 ( .A(n15194), .B(n15635), .Z(n15198) );
  XOR U2061 ( .A(n15775), .B(n16258), .Z(n15779) );
  XOR U2062 ( .A(n14517), .B(n15024), .Z(n14521) );
  XOR U2063 ( .A(n13235), .B(n13766), .Z(n13239) );
  XOR U2064 ( .A(n11862), .B(n12497), .Z(n11866) );
  XOR U2065 ( .A(n39458), .B(n39754), .Z(n39462) );
  XOR U2066 ( .A(n38834), .B(n39130), .Z(n38838) );
  XOR U2067 ( .A(n18334), .B(n18685), .Z(n18338) );
  XOR U2068 ( .A(n10557), .B(n11184), .Z(n10561) );
  XOR U2069 ( .A(n13220), .B(n13769), .Z(n13224) );
  XOR U2070 ( .A(n11250), .B(n11835), .Z(n11254) );
  XOR U2071 ( .A(n15805), .B(n16252), .Z(n15809) );
  XOR U2072 ( .A(n14547), .B(n15018), .Z(n14551) );
  XOR U2073 ( .A(n13265), .B(n13760), .Z(n13269) );
  XOR U2074 ( .A(n17692), .B(n18049), .Z(n17696) );
  XOR U2075 ( .A(n16470), .B(n16851), .Z(n16474) );
  XOR U2076 ( .A(n15224), .B(n15629), .Z(n15228) );
  XOR U2077 ( .A(n17129), .B(n17444), .Z(n17133) );
  XOR U2078 ( .A(n38518), .B(n38808), .Z(n38522) );
  XOR U2079 ( .A(n37858), .B(n38148), .Z(n37862) );
  XOR U2080 ( .A(n37174), .B(n37464), .Z(n37178) );
  XOR U2081 ( .A(n36466), .B(n36756), .Z(n36470) );
  XOR U2082 ( .A(n35734), .B(n36024), .Z(n35738) );
  XOR U2083 ( .A(n34978), .B(n35268), .Z(n34982) );
  XOR U2084 ( .A(n34198), .B(n34488), .Z(n34202) );
  XOR U2085 ( .A(n33394), .B(n33684), .Z(n33398) );
  XOR U2086 ( .A(n32566), .B(n32856), .Z(n32570) );
  XOR U2087 ( .A(n31714), .B(n32004), .Z(n31718) );
  XOR U2088 ( .A(n30838), .B(n31128), .Z(n30842) );
  XOR U2089 ( .A(n29938), .B(n30228), .Z(n29942) );
  XOR U2090 ( .A(n29014), .B(n29304), .Z(n29018) );
  XOR U2091 ( .A(n28066), .B(n28356), .Z(n28070) );
  XOR U2092 ( .A(n27094), .B(n27384), .Z(n27098) );
  XOR U2093 ( .A(n26096), .B(n26386), .Z(n26100) );
  XOR U2094 ( .A(n25074), .B(n25364), .Z(n25078) );
  XOR U2095 ( .A(n24026), .B(n24316), .Z(n24030) );
  XOR U2096 ( .A(n22957), .B(n23247), .Z(n22961) );
  XOR U2097 ( .A(n21864), .B(n22154), .Z(n21868) );
  XOR U2098 ( .A(n20747), .B(n21037), .Z(n20751) );
  XOR U2099 ( .A(n19607), .B(n19897), .Z(n19611) );
  XOR U2100 ( .A(n11892), .B(n12491), .Z(n11896) );
  XOR U2101 ( .A(n17722), .B(n18043), .Z(n17726) );
  XOR U2102 ( .A(n16500), .B(n16845), .Z(n16504) );
  XOR U2103 ( .A(n15254), .B(n15623), .Z(n15258) );
  XOR U2104 ( .A(n15835), .B(n16246), .Z(n15839) );
  XOR U2105 ( .A(n14577), .B(n15012), .Z(n14581) );
  XOR U2106 ( .A(n13295), .B(n13754), .Z(n13299) );
  XOR U2107 ( .A(n13894), .B(n14395), .Z(n13898) );
  XOR U2108 ( .A(n12600), .B(n13125), .Z(n12604) );
  XOR U2109 ( .A(n9873), .B(n10524), .Z(n9877) );
  XOR U2110 ( .A(n17747), .B(n18038), .Z(n17751) );
  XOR U2111 ( .A(n40364), .B(n40642), .Z(n40368) );
  XOR U2112 ( .A(n39776), .B(n40054), .Z(n39780) );
  XOR U2113 ( .A(n17159), .B(n17438), .Z(n17163) );
  XOR U2114 ( .A(n11285), .B(n11828), .Z(n11289) );
  XOR U2115 ( .A(n11927), .B(n12484), .Z(n11931) );
  XOR U2116 ( .A(n10597), .B(n11176), .Z(n10601) );
  XOR U2117 ( .A(n13924), .B(n14389), .Z(n13928) );
  XOR U2118 ( .A(n12630), .B(n13119), .Z(n12634) );
  XOR U2119 ( .A(n11310), .B(n11823), .Z(n11314) );
  XOR U2120 ( .A(n15865), .B(n16240), .Z(n15869) );
  XOR U2121 ( .A(n14607), .B(n15006), .Z(n14611) );
  XOR U2122 ( .A(n13325), .B(n13748), .Z(n13329) );
  XOR U2123 ( .A(n16530), .B(n16839), .Z(n16534) );
  XOR U2124 ( .A(n15284), .B(n15617), .Z(n15288) );
  XNOR U2125 ( .A(n40084), .B(n39784), .Z(n39786) );
  XOR U2126 ( .A(n39169), .B(n39441), .Z(n39173) );
  XOR U2127 ( .A(n38533), .B(n38805), .Z(n38537) );
  XOR U2128 ( .A(n37873), .B(n38145), .Z(n37877) );
  XOR U2129 ( .A(n37189), .B(n37461), .Z(n37193) );
  XOR U2130 ( .A(n36481), .B(n36753), .Z(n36485) );
  XOR U2131 ( .A(n35749), .B(n36021), .Z(n35753) );
  XOR U2132 ( .A(n34993), .B(n35265), .Z(n34997) );
  XOR U2133 ( .A(n34213), .B(n34485), .Z(n34217) );
  XOR U2134 ( .A(n33409), .B(n33681), .Z(n33413) );
  XOR U2135 ( .A(n32581), .B(n32853), .Z(n32585) );
  XOR U2136 ( .A(n31729), .B(n32001), .Z(n31733) );
  XOR U2137 ( .A(n30853), .B(n31125), .Z(n30857) );
  XOR U2138 ( .A(n29953), .B(n30225), .Z(n29957) );
  XOR U2139 ( .A(n29029), .B(n29301), .Z(n29033) );
  XOR U2140 ( .A(n28081), .B(n28353), .Z(n28085) );
  XOR U2141 ( .A(n27109), .B(n27381), .Z(n27113) );
  XOR U2142 ( .A(n26111), .B(n26383), .Z(n26115) );
  XOR U2143 ( .A(n25089), .B(n25361), .Z(n25093) );
  XOR U2144 ( .A(n24041), .B(n24313), .Z(n24045) );
  XOR U2145 ( .A(n22972), .B(n23244), .Z(n22976) );
  XOR U2146 ( .A(n21879), .B(n22151), .Z(n21883) );
  XOR U2147 ( .A(n20762), .B(n21034), .Z(n20766) );
  XOR U2148 ( .A(n19622), .B(n19894), .Z(n19626) );
  XOR U2149 ( .A(n9903), .B(n10518), .Z(n9907) );
  XOR U2150 ( .A(n8537), .B(n9176), .Z(n8541) );
  XOR U2151 ( .A(n9248), .B(n9845), .Z(n9252) );
  XOR U2152 ( .A(n15314), .B(n15611), .Z(n15318) );
  XOR U2153 ( .A(n15895), .B(n16234), .Z(n15899) );
  XOR U2154 ( .A(n14637), .B(n15000), .Z(n14641) );
  XOR U2155 ( .A(n13355), .B(n13742), .Z(n13359) );
  XOR U2156 ( .A(n13954), .B(n14383), .Z(n13958) );
  XOR U2157 ( .A(n12660), .B(n13113), .Z(n12664) );
  XOR U2158 ( .A(n11340), .B(n11817), .Z(n11344) );
  XOR U2159 ( .A(n11957), .B(n12478), .Z(n11961) );
  XOR U2160 ( .A(n7830), .B(n8499), .Z(n7834) );
  XOR U2161 ( .A(n41216), .B(n41476), .Z(n41220) );
  XOR U2162 ( .A(n40664), .B(n40924), .Z(n40668) );
  XOR U2163 ( .A(n18364), .B(n18673), .Z(n18368) );
  XOR U2164 ( .A(n17174), .B(n17435), .Z(n17178) );
  XOR U2165 ( .A(n9958), .B(n10507), .Z(n9962) );
  XOR U2166 ( .A(n8592), .B(n9165), .Z(n8596) );
  XOR U2167 ( .A(n6453), .B(n7116), .Z(n6457) );
  XOR U2168 ( .A(n9938), .B(n10511), .Z(n9942) );
  XOR U2169 ( .A(n11987), .B(n12472), .Z(n11991) );
  XOR U2170 ( .A(n13984), .B(n14377), .Z(n13988) );
  XOR U2171 ( .A(n12690), .B(n13107), .Z(n12694) );
  XOR U2172 ( .A(n11370), .B(n11811), .Z(n11374) );
  XOR U2173 ( .A(n15925), .B(n16228), .Z(n15929) );
  XOR U2174 ( .A(n14667), .B(n14994), .Z(n14671) );
  XOR U2175 ( .A(n13385), .B(n13736), .Z(n13389) );
  XOR U2176 ( .A(n15344), .B(n15605), .Z(n15348) );
  XOR U2177 ( .A(n40384), .B(n40638), .Z(n40388) );
  XOR U2178 ( .A(n39796), .B(n40050), .Z(n39800) );
  XOR U2179 ( .A(n39184), .B(n39438), .Z(n39188) );
  XOR U2180 ( .A(n38548), .B(n38802), .Z(n38552) );
  XOR U2181 ( .A(n37888), .B(n38142), .Z(n37892) );
  XOR U2182 ( .A(n37204), .B(n37458), .Z(n37208) );
  XOR U2183 ( .A(n36496), .B(n36750), .Z(n36500) );
  XOR U2184 ( .A(n35764), .B(n36018), .Z(n35768) );
  XOR U2185 ( .A(n35008), .B(n35262), .Z(n35012) );
  XOR U2186 ( .A(n34228), .B(n34482), .Z(n34232) );
  XOR U2187 ( .A(n33424), .B(n33678), .Z(n33428) );
  XOR U2188 ( .A(n32596), .B(n32850), .Z(n32600) );
  XOR U2189 ( .A(n31744), .B(n31998), .Z(n31748) );
  XOR U2190 ( .A(n30868), .B(n31122), .Z(n30872) );
  XOR U2191 ( .A(n29968), .B(n30222), .Z(n29972) );
  XOR U2192 ( .A(n29044), .B(n29298), .Z(n29048) );
  XOR U2193 ( .A(n28096), .B(n28350), .Z(n28100) );
  XOR U2194 ( .A(n27124), .B(n27378), .Z(n27128) );
  XOR U2195 ( .A(n26126), .B(n26380), .Z(n26130) );
  XOR U2196 ( .A(n25104), .B(n25358), .Z(n25108) );
  XOR U2197 ( .A(n24056), .B(n24310), .Z(n24060) );
  XOR U2198 ( .A(n22987), .B(n23241), .Z(n22991) );
  XOR U2199 ( .A(n21894), .B(n22148), .Z(n21898) );
  XOR U2200 ( .A(n20777), .B(n21031), .Z(n20781) );
  XOR U2201 ( .A(n19637), .B(n19891), .Z(n19641) );
  XOR U2202 ( .A(n8552), .B(n9173), .Z(n8556) );
  XOR U2203 ( .A(n7885), .B(n8488), .Z(n7889) );
  XOR U2204 ( .A(n6483), .B(n7110), .Z(n6487) );
  XOR U2205 ( .A(n9988), .B(n10501), .Z(n9992) );
  XOR U2206 ( .A(n8622), .B(n9159), .Z(n8626) );
  XOR U2207 ( .A(n15955), .B(n16222), .Z(n15959) );
  XOR U2208 ( .A(n14697), .B(n14988), .Z(n14701) );
  XOR U2209 ( .A(n13415), .B(n13730), .Z(n13419) );
  XOR U2210 ( .A(n14014), .B(n14371), .Z(n14018) );
  XOR U2211 ( .A(n12720), .B(n13101), .Z(n12724) );
  XOR U2212 ( .A(n11400), .B(n11805), .Z(n11404) );
  XOR U2213 ( .A(n12017), .B(n12466), .Z(n12021) );
  XOR U2214 ( .A(n7167), .B(n7806), .Z(n7171) );
  XOR U2215 ( .A(n5733), .B(n6420), .Z(n5737) );
  XOR U2216 ( .A(n42014), .B(n42256), .Z(n42018) );
  XOR U2217 ( .A(n41498), .B(n41740), .Z(n41502) );
  XOR U2218 ( .A(n17787), .B(n18030), .Z(n17791) );
  XOR U2219 ( .A(n16585), .B(n16828), .Z(n16589) );
  XOR U2220 ( .A(n10018), .B(n10495), .Z(n10022) );
  XOR U2221 ( .A(n8652), .B(n9153), .Z(n8656) );
  XOR U2222 ( .A(n7915), .B(n8482), .Z(n7919) );
  XOR U2223 ( .A(n6513), .B(n7104), .Z(n6517) );
  XOR U2224 ( .A(n4318), .B(n4999), .Z(n4322) );
  XOR U2225 ( .A(n12047), .B(n12460), .Z(n12051) );
  XOR U2226 ( .A(n14044), .B(n14365), .Z(n14048) );
  XOR U2227 ( .A(n12750), .B(n13095), .Z(n12754) );
  XOR U2228 ( .A(n11430), .B(n11799), .Z(n11434) );
  XOR U2229 ( .A(n14727), .B(n14982), .Z(n14731) );
  XOR U2230 ( .A(n13445), .B(n13724), .Z(n13449) );
  XNOR U2231 ( .A(n41770), .B(n41506), .Z(n41508) );
  XOR U2232 ( .A(n40963), .B(n41199), .Z(n40967) );
  XOR U2233 ( .A(n40399), .B(n40635), .Z(n40403) );
  XOR U2234 ( .A(n39811), .B(n40047), .Z(n39815) );
  XOR U2235 ( .A(n39199), .B(n39435), .Z(n39203) );
  XOR U2236 ( .A(n38563), .B(n38799), .Z(n38567) );
  XOR U2237 ( .A(n37903), .B(n38139), .Z(n37907) );
  XOR U2238 ( .A(n37219), .B(n37455), .Z(n37223) );
  XOR U2239 ( .A(n36511), .B(n36747), .Z(n36515) );
  XOR U2240 ( .A(n35779), .B(n36015), .Z(n35783) );
  XOR U2241 ( .A(n35023), .B(n35259), .Z(n35027) );
  XOR U2242 ( .A(n34243), .B(n34479), .Z(n34247) );
  XOR U2243 ( .A(n33439), .B(n33675), .Z(n33443) );
  XOR U2244 ( .A(n32611), .B(n32847), .Z(n32615) );
  XOR U2245 ( .A(n31759), .B(n31995), .Z(n31763) );
  XOR U2246 ( .A(n30883), .B(n31119), .Z(n30887) );
  XOR U2247 ( .A(n29983), .B(n30219), .Z(n29987) );
  XOR U2248 ( .A(n29059), .B(n29295), .Z(n29063) );
  XOR U2249 ( .A(n28111), .B(n28347), .Z(n28115) );
  XOR U2250 ( .A(n27139), .B(n27375), .Z(n27143) );
  XOR U2251 ( .A(n26141), .B(n26377), .Z(n26145) );
  XOR U2252 ( .A(n25119), .B(n25355), .Z(n25123) );
  XOR U2253 ( .A(n24071), .B(n24307), .Z(n24075) );
  XOR U2254 ( .A(n23002), .B(n23238), .Z(n23006) );
  XOR U2255 ( .A(n21909), .B(n22145), .Z(n21913) );
  XOR U2256 ( .A(n20792), .B(n21028), .Z(n20796) );
  XOR U2257 ( .A(n19652), .B(n19888), .Z(n19656) );
  XOR U2258 ( .A(n5788), .B(n6409), .Z(n5792) );
  XOR U2259 ( .A(n4348), .B(n4993), .Z(n4352) );
  XOR U2260 ( .A(n7945), .B(n8476), .Z(n7949) );
  XOR U2261 ( .A(n6543), .B(n7098), .Z(n6547) );
  XOR U2262 ( .A(n10048), .B(n10489), .Z(n10052) );
  XOR U2263 ( .A(n8682), .B(n9147), .Z(n8686) );
  XOR U2264 ( .A(n13475), .B(n13718), .Z(n13479) );
  XOR U2265 ( .A(n14074), .B(n14359), .Z(n14078) );
  XOR U2266 ( .A(n12780), .B(n13089), .Z(n12784) );
  XOR U2267 ( .A(n11460), .B(n11793), .Z(n11464) );
  XOR U2268 ( .A(n12077), .B(n12454), .Z(n12081) );
  XOR U2269 ( .A(n5768), .B(n6413), .Z(n5772) );
  XOR U2270 ( .A(n3580), .B(n4285), .Z(n3584) );
  XOR U2271 ( .A(n42758), .B(n42982), .Z(n42762) );
  XOR U2272 ( .A(n42278), .B(n42502), .Z(n42282) );
  XOR U2273 ( .A(n18394), .B(n18661), .Z(n18398) );
  XOR U2274 ( .A(n17204), .B(n17429), .Z(n17208) );
  XOR U2275 ( .A(n15990), .B(n16215), .Z(n15994) );
  XOR U2276 ( .A(n10078), .B(n10483), .Z(n10082) );
  XOR U2277 ( .A(n8712), .B(n9141), .Z(n8716) );
  XOR U2278 ( .A(n7975), .B(n8470), .Z(n7979) );
  XOR U2279 ( .A(n6573), .B(n7092), .Z(n6577) );
  XOR U2280 ( .A(n5818), .B(n6403), .Z(n5822) );
  XOR U2281 ( .A(n4378), .B(n4987), .Z(n4382) );
  XOR U2282 ( .A(n4333), .B(n4996), .Z(n4337) );
  XOR U2283 ( .A(n2871), .B(n3558), .Z(n2875) );
  XOR U2284 ( .A(n2111), .B(n2834), .Z(n2115) );
  XOR U2285 ( .A(n12107), .B(n12448), .Z(n12111) );
  XOR U2286 ( .A(n14104), .B(n14353), .Z(n14108) );
  XOR U2287 ( .A(n12810), .B(n13083), .Z(n12814) );
  XOR U2288 ( .A(n11490), .B(n11787), .Z(n11494) );
  XOR U2289 ( .A(n42034), .B(n42252), .Z(n42038) );
  XOR U2290 ( .A(n41518), .B(n41736), .Z(n41522) );
  XOR U2291 ( .A(n40978), .B(n41196), .Z(n40982) );
  XOR U2292 ( .A(n40414), .B(n40632), .Z(n40418) );
  XOR U2293 ( .A(n39826), .B(n40044), .Z(n39830) );
  XOR U2294 ( .A(n39214), .B(n39432), .Z(n39218) );
  XOR U2295 ( .A(n38578), .B(n38796), .Z(n38582) );
  XOR U2296 ( .A(n37918), .B(n38136), .Z(n37922) );
  XOR U2297 ( .A(n37234), .B(n37452), .Z(n37238) );
  XOR U2298 ( .A(n36526), .B(n36744), .Z(n36530) );
  XOR U2299 ( .A(n35794), .B(n36012), .Z(n35798) );
  XOR U2300 ( .A(n35038), .B(n35256), .Z(n35042) );
  XOR U2301 ( .A(n34258), .B(n34476), .Z(n34262) );
  XOR U2302 ( .A(n33454), .B(n33672), .Z(n33458) );
  XOR U2303 ( .A(n32626), .B(n32844), .Z(n32630) );
  XOR U2304 ( .A(n31774), .B(n31992), .Z(n31778) );
  XOR U2305 ( .A(n30898), .B(n31116), .Z(n30902) );
  XOR U2306 ( .A(n29998), .B(n30216), .Z(n30002) );
  XOR U2307 ( .A(n29074), .B(n29292), .Z(n29078) );
  XOR U2308 ( .A(n28126), .B(n28344), .Z(n28130) );
  XOR U2309 ( .A(n27154), .B(n27372), .Z(n27158) );
  XOR U2310 ( .A(n26156), .B(n26374), .Z(n26160) );
  XOR U2311 ( .A(n25134), .B(n25352), .Z(n25138) );
  XOR U2312 ( .A(n24086), .B(n24304), .Z(n24090) );
  XOR U2313 ( .A(n23017), .B(n23235), .Z(n23021) );
  XOR U2314 ( .A(n21924), .B(n22142), .Z(n21928) );
  XOR U2315 ( .A(n20807), .B(n21025), .Z(n20811) );
  XOR U2316 ( .A(n19667), .B(n19885), .Z(n19671) );
  XOR U2317 ( .A(n3635), .B(n4274), .Z(n3639) );
  XOR U2318 ( .A(n2161), .B(n2824), .Z(n2165) );
  XOR U2319 ( .A(n5848), .B(n6397), .Z(n5852) );
  XOR U2320 ( .A(n4408), .B(n4981), .Z(n4412) );
  XOR U2321 ( .A(n8005), .B(n8464), .Z(n8009) );
  XOR U2322 ( .A(n6603), .B(n7086), .Z(n6607) );
  XOR U2323 ( .A(n10108), .B(n10477), .Z(n10112) );
  XOR U2324 ( .A(n8742), .B(n9135), .Z(n8746) );
  XOR U2325 ( .A(n12840), .B(n13077), .Z(n12844) );
  XOR U2326 ( .A(n11520), .B(n11781), .Z(n11524) );
  XOR U2327 ( .A(n12137), .B(n12442), .Z(n12141) );
  XOR U2328 ( .A(n43448), .B(n43654), .Z(n43452) );
  XOR U2329 ( .A(n43004), .B(n43210), .Z(n43008) );
  XOR U2330 ( .A(n17817), .B(n18024), .Z(n17821) );
  XOR U2331 ( .A(n16615), .B(n16822), .Z(n16619) );
  XOR U2332 ( .A(n15389), .B(n15596), .Z(n15393) );
  XOR U2333 ( .A(n12865), .B(n13072), .Z(n12869) );
  XOR U2334 ( .A(n14139), .B(n14346), .Z(n14143) );
  XOR U2335 ( .A(n10138), .B(n10471), .Z(n10142) );
  XOR U2336 ( .A(n8772), .B(n9129), .Z(n8776) );
  XOR U2337 ( .A(n8035), .B(n8458), .Z(n8039) );
  XOR U2338 ( .A(n6633), .B(n7080), .Z(n6637) );
  XOR U2339 ( .A(n5878), .B(n6391), .Z(n5882) );
  XOR U2340 ( .A(n4438), .B(n4975), .Z(n4442) );
  XOR U2341 ( .A(n3665), .B(n4268), .Z(n3669) );
  XOR U2342 ( .A(n2191), .B(n2818), .Z(n2195) );
  XOR U2343 ( .A(n2146), .B(n2827), .Z(n2150) );
  XOR U2344 ( .A(n12167), .B(n12436), .Z(n12171) );
  XOR U2345 ( .A(n11550), .B(n11775), .Z(n11554) );
  XNOR U2346 ( .A(n43240), .B(n43012), .Z(n43014) );
  XOR U2347 ( .A(n42541), .B(n42741), .Z(n42545) );
  XOR U2348 ( .A(n42049), .B(n42249), .Z(n42053) );
  XOR U2349 ( .A(n41533), .B(n41733), .Z(n41537) );
  XOR U2350 ( .A(n40993), .B(n41193), .Z(n40997) );
  XOR U2351 ( .A(n40429), .B(n40629), .Z(n40433) );
  XOR U2352 ( .A(n39841), .B(n40041), .Z(n39845) );
  XOR U2353 ( .A(n39229), .B(n39429), .Z(n39233) );
  XOR U2354 ( .A(n38593), .B(n38793), .Z(n38597) );
  XOR U2355 ( .A(n37933), .B(n38133), .Z(n37937) );
  XOR U2356 ( .A(n37249), .B(n37449), .Z(n37253) );
  XOR U2357 ( .A(n36541), .B(n36741), .Z(n36545) );
  XOR U2358 ( .A(n35809), .B(n36009), .Z(n35813) );
  XOR U2359 ( .A(n35053), .B(n35253), .Z(n35057) );
  XOR U2360 ( .A(n34273), .B(n34473), .Z(n34277) );
  XOR U2361 ( .A(n33469), .B(n33669), .Z(n33473) );
  XOR U2362 ( .A(n32641), .B(n32841), .Z(n32645) );
  XOR U2363 ( .A(n31789), .B(n31989), .Z(n31793) );
  XOR U2364 ( .A(n30913), .B(n31113), .Z(n30917) );
  XOR U2365 ( .A(n30013), .B(n30213), .Z(n30017) );
  XOR U2366 ( .A(n29089), .B(n29289), .Z(n29093) );
  XOR U2367 ( .A(n28141), .B(n28341), .Z(n28145) );
  XOR U2368 ( .A(n27169), .B(n27369), .Z(n27173) );
  XOR U2369 ( .A(n26171), .B(n26371), .Z(n26175) );
  XOR U2370 ( .A(n25149), .B(n25349), .Z(n25153) );
  XOR U2371 ( .A(n24101), .B(n24301), .Z(n24105) );
  XOR U2372 ( .A(n23032), .B(n23232), .Z(n23036) );
  XOR U2373 ( .A(n21939), .B(n22139), .Z(n21943) );
  XOR U2374 ( .A(n20822), .B(n21022), .Z(n20826) );
  XOR U2375 ( .A(n19682), .B(n19882), .Z(n19686) );
  XOR U2376 ( .A(n2176), .B(n2821), .Z(n2180) );
  XOR U2377 ( .A(n3695), .B(n4262), .Z(n3699) );
  XOR U2378 ( .A(n2221), .B(n2812), .Z(n2225) );
  XOR U2379 ( .A(n5908), .B(n6385), .Z(n5912) );
  XOR U2380 ( .A(n4468), .B(n4969), .Z(n4472) );
  XOR U2381 ( .A(n8065), .B(n8452), .Z(n8069) );
  XOR U2382 ( .A(n6663), .B(n7074), .Z(n6667) );
  XOR U2383 ( .A(n10168), .B(n10465), .Z(n10172) );
  XOR U2384 ( .A(n8802), .B(n9123), .Z(n8806) );
  XOR U2385 ( .A(n12197), .B(n12430), .Z(n12201) );
  XOR U2386 ( .A(n44084), .B(n44272), .Z(n44088) );
  XOR U2387 ( .A(n43676), .B(n43864), .Z(n43680) );
  XOR U2388 ( .A(n18424), .B(n18649), .Z(n18428) );
  XOR U2389 ( .A(n17234), .B(n17423), .Z(n17238) );
  XOR U2390 ( .A(n16020), .B(n16209), .Z(n16024) );
  XOR U2391 ( .A(n14782), .B(n14971), .Z(n14786) );
  XOR U2392 ( .A(n13520), .B(n13709), .Z(n13524) );
  XOR U2393 ( .A(n10198), .B(n10459), .Z(n10202) );
  XOR U2394 ( .A(n8832), .B(n9117), .Z(n8836) );
  XOR U2395 ( .A(n8095), .B(n8446), .Z(n8099) );
  XOR U2396 ( .A(n6693), .B(n7068), .Z(n6697) );
  XOR U2397 ( .A(n5938), .B(n6379), .Z(n5942) );
  XOR U2398 ( .A(n4498), .B(n4963), .Z(n4502) );
  XOR U2399 ( .A(n3725), .B(n4256), .Z(n3729) );
  XOR U2400 ( .A(n2251), .B(n2806), .Z(n2255) );
  XOR U2401 ( .A(n2206), .B(n2815), .Z(n2210) );
  XOR U2402 ( .A(n43468), .B(n43650), .Z(n43472) );
  XOR U2403 ( .A(n43024), .B(n43206), .Z(n43028) );
  XOR U2404 ( .A(n42556), .B(n42738), .Z(n42560) );
  XOR U2405 ( .A(n42064), .B(n42246), .Z(n42068) );
  XOR U2406 ( .A(n41548), .B(n41730), .Z(n41552) );
  XOR U2407 ( .A(n41008), .B(n41190), .Z(n41012) );
  XOR U2408 ( .A(n40444), .B(n40626), .Z(n40448) );
  XOR U2409 ( .A(n39856), .B(n40038), .Z(n39860) );
  XOR U2410 ( .A(n39244), .B(n39426), .Z(n39248) );
  XOR U2411 ( .A(n38608), .B(n38790), .Z(n38612) );
  XOR U2412 ( .A(n37948), .B(n38130), .Z(n37952) );
  XOR U2413 ( .A(n37264), .B(n37446), .Z(n37268) );
  XOR U2414 ( .A(n36556), .B(n36738), .Z(n36560) );
  XOR U2415 ( .A(n35824), .B(n36006), .Z(n35828) );
  XOR U2416 ( .A(n35068), .B(n35250), .Z(n35072) );
  XOR U2417 ( .A(n34288), .B(n34470), .Z(n34292) );
  XOR U2418 ( .A(n33484), .B(n33666), .Z(n33488) );
  XOR U2419 ( .A(n32656), .B(n32838), .Z(n32660) );
  XOR U2420 ( .A(n31804), .B(n31986), .Z(n31808) );
  XOR U2421 ( .A(n30928), .B(n31110), .Z(n30932) );
  XOR U2422 ( .A(n30028), .B(n30210), .Z(n30032) );
  XOR U2423 ( .A(n29104), .B(n29286), .Z(n29108) );
  XOR U2424 ( .A(n28156), .B(n28338), .Z(n28160) );
  XOR U2425 ( .A(n27184), .B(n27366), .Z(n27188) );
  XOR U2426 ( .A(n26186), .B(n26368), .Z(n26190) );
  XOR U2427 ( .A(n25164), .B(n25346), .Z(n25168) );
  XOR U2428 ( .A(n24116), .B(n24298), .Z(n24120) );
  XOR U2429 ( .A(n23047), .B(n23229), .Z(n23051) );
  XOR U2430 ( .A(n21954), .B(n22136), .Z(n21958) );
  XOR U2431 ( .A(n20837), .B(n21019), .Z(n20841) );
  XOR U2432 ( .A(n19697), .B(n19879), .Z(n19701) );
  XOR U2433 ( .A(n12237), .B(n12422), .Z(n12241) );
  XOR U2434 ( .A(n2236), .B(n2809), .Z(n2240) );
  XOR U2435 ( .A(n3755), .B(n4250), .Z(n3759) );
  XOR U2436 ( .A(n2281), .B(n2800), .Z(n2285) );
  XOR U2437 ( .A(n5968), .B(n6373), .Z(n5972) );
  XOR U2438 ( .A(n4528), .B(n4957), .Z(n4532) );
  XOR U2439 ( .A(n8125), .B(n8440), .Z(n8129) );
  XOR U2440 ( .A(n6723), .B(n7062), .Z(n6727) );
  XOR U2441 ( .A(n10228), .B(n10453), .Z(n10232) );
  XOR U2442 ( .A(n8862), .B(n9111), .Z(n8866) );
  XOR U2443 ( .A(n44666), .B(n44836), .Z(n44670) );
  XOR U2444 ( .A(n44294), .B(n44464), .Z(n44298) );
  XOR U2445 ( .A(n17847), .B(n18018), .Z(n17851) );
  XOR U2446 ( .A(n16645), .B(n16816), .Z(n16649) );
  XOR U2447 ( .A(n15419), .B(n15590), .Z(n15423) );
  XOR U2448 ( .A(n14169), .B(n14340), .Z(n14173) );
  XOR U2449 ( .A(n10258), .B(n10447), .Z(n10262) );
  XOR U2450 ( .A(n8892), .B(n9105), .Z(n8896) );
  XOR U2451 ( .A(n8155), .B(n8434), .Z(n8159) );
  XOR U2452 ( .A(n6753), .B(n7056), .Z(n6757) );
  XOR U2453 ( .A(n5998), .B(n6367), .Z(n6002) );
  XOR U2454 ( .A(n4558), .B(n4951), .Z(n4562) );
  XOR U2455 ( .A(n3785), .B(n4244), .Z(n3789) );
  XOR U2456 ( .A(n2311), .B(n2794), .Z(n2315) );
  XOR U2457 ( .A(n2266), .B(n2803), .Z(n2270) );
  XNOR U2458 ( .A(n44494), .B(n44302), .Z(n44304) );
  XOR U2459 ( .A(n43903), .B(n44067), .Z(n43907) );
  XOR U2460 ( .A(n43483), .B(n43647), .Z(n43487) );
  XOR U2461 ( .A(n43039), .B(n43203), .Z(n43043) );
  XOR U2462 ( .A(n42571), .B(n42735), .Z(n42575) );
  XOR U2463 ( .A(n42079), .B(n42243), .Z(n42083) );
  XOR U2464 ( .A(n41563), .B(n41727), .Z(n41567) );
  XOR U2465 ( .A(n41023), .B(n41187), .Z(n41027) );
  XOR U2466 ( .A(n40459), .B(n40623), .Z(n40463) );
  XOR U2467 ( .A(n39871), .B(n40035), .Z(n39875) );
  XOR U2468 ( .A(n39259), .B(n39423), .Z(n39263) );
  XOR U2469 ( .A(n38623), .B(n38787), .Z(n38627) );
  XOR U2470 ( .A(n37963), .B(n38127), .Z(n37967) );
  XOR U2471 ( .A(n37279), .B(n37443), .Z(n37283) );
  XOR U2472 ( .A(n36571), .B(n36735), .Z(n36575) );
  XOR U2473 ( .A(n35839), .B(n36003), .Z(n35843) );
  XOR U2474 ( .A(n35083), .B(n35247), .Z(n35087) );
  XOR U2475 ( .A(n34303), .B(n34467), .Z(n34307) );
  XOR U2476 ( .A(n33499), .B(n33663), .Z(n33503) );
  XOR U2477 ( .A(n32671), .B(n32835), .Z(n32675) );
  XOR U2478 ( .A(n31819), .B(n31983), .Z(n31823) );
  XOR U2479 ( .A(n30943), .B(n31107), .Z(n30947) );
  XOR U2480 ( .A(n30043), .B(n30207), .Z(n30047) );
  XOR U2481 ( .A(n29119), .B(n29283), .Z(n29123) );
  XOR U2482 ( .A(n28171), .B(n28335), .Z(n28175) );
  XOR U2483 ( .A(n27199), .B(n27363), .Z(n27203) );
  XOR U2484 ( .A(n26201), .B(n26365), .Z(n26205) );
  XOR U2485 ( .A(n25179), .B(n25343), .Z(n25183) );
  XOR U2486 ( .A(n24131), .B(n24295), .Z(n24135) );
  XOR U2487 ( .A(n23062), .B(n23226), .Z(n23066) );
  XOR U2488 ( .A(n21969), .B(n22133), .Z(n21973) );
  XOR U2489 ( .A(n20852), .B(n21016), .Z(n20856) );
  XOR U2490 ( .A(n19712), .B(n19876), .Z(n19716) );
  XOR U2491 ( .A(n12900), .B(n13065), .Z(n12904) );
  XOR U2492 ( .A(n11600), .B(n11765), .Z(n11604) );
  XOR U2493 ( .A(n2296), .B(n2797), .Z(n2300) );
  XOR U2494 ( .A(n3815), .B(n4238), .Z(n3819) );
  XOR U2495 ( .A(n2341), .B(n2788), .Z(n2345) );
  XOR U2496 ( .A(n6028), .B(n6361), .Z(n6032) );
  XOR U2497 ( .A(n4588), .B(n4945), .Z(n4592) );
  XOR U2498 ( .A(n8185), .B(n8428), .Z(n8189) );
  XOR U2499 ( .A(n6783), .B(n7050), .Z(n6787) );
  XOR U2500 ( .A(n8922), .B(n9099), .Z(n8926) );
  XOR U2501 ( .A(n10283), .B(n10442), .Z(n10287) );
  XOR U2502 ( .A(n45194), .B(n45346), .Z(n45198) );
  XOR U2503 ( .A(n44858), .B(n45010), .Z(n44862) );
  XOR U2504 ( .A(n18454), .B(n18637), .Z(n18458) );
  XOR U2505 ( .A(n17264), .B(n17417), .Z(n17268) );
  XOR U2506 ( .A(n16050), .B(n16203), .Z(n16054) );
  XOR U2507 ( .A(n8215), .B(n8422), .Z(n8219) );
  XOR U2508 ( .A(n6813), .B(n7044), .Z(n6817) );
  XOR U2509 ( .A(n6058), .B(n6355), .Z(n6062) );
  XOR U2510 ( .A(n4618), .B(n4939), .Z(n4622) );
  XOR U2511 ( .A(n3845), .B(n4232), .Z(n3849) );
  XOR U2512 ( .A(n2371), .B(n2782), .Z(n2375) );
  XOR U2513 ( .A(n2326), .B(n2791), .Z(n2330) );
  XOR U2514 ( .A(n9618), .B(n9771), .Z(n9622) );
  XOR U2515 ( .A(n44686), .B(n44832), .Z(n44690) );
  XOR U2516 ( .A(n44314), .B(n44460), .Z(n44318) );
  XOR U2517 ( .A(n43918), .B(n44064), .Z(n43922) );
  XOR U2518 ( .A(n43498), .B(n43644), .Z(n43502) );
  XOR U2519 ( .A(n43054), .B(n43200), .Z(n43058) );
  XOR U2520 ( .A(n42586), .B(n42732), .Z(n42590) );
  XOR U2521 ( .A(n42094), .B(n42240), .Z(n42098) );
  XOR U2522 ( .A(n41578), .B(n41724), .Z(n41582) );
  XOR U2523 ( .A(n41038), .B(n41184), .Z(n41042) );
  XOR U2524 ( .A(n40474), .B(n40620), .Z(n40478) );
  XOR U2525 ( .A(n39886), .B(n40032), .Z(n39890) );
  XOR U2526 ( .A(n39274), .B(n39420), .Z(n39278) );
  XOR U2527 ( .A(n38638), .B(n38784), .Z(n38642) );
  XOR U2528 ( .A(n37978), .B(n38124), .Z(n37982) );
  XOR U2529 ( .A(n37294), .B(n37440), .Z(n37298) );
  XOR U2530 ( .A(n36586), .B(n36732), .Z(n36590) );
  XOR U2531 ( .A(n35854), .B(n36000), .Z(n35858) );
  XOR U2532 ( .A(n35098), .B(n35244), .Z(n35102) );
  XOR U2533 ( .A(n34318), .B(n34464), .Z(n34322) );
  XOR U2534 ( .A(n33514), .B(n33660), .Z(n33518) );
  XOR U2535 ( .A(n32686), .B(n32832), .Z(n32690) );
  XOR U2536 ( .A(n31834), .B(n31980), .Z(n31838) );
  XOR U2537 ( .A(n30958), .B(n31104), .Z(n30962) );
  XOR U2538 ( .A(n30058), .B(n30204), .Z(n30062) );
  XOR U2539 ( .A(n29134), .B(n29280), .Z(n29138) );
  XOR U2540 ( .A(n28186), .B(n28332), .Z(n28190) );
  XOR U2541 ( .A(n27214), .B(n27360), .Z(n27218) );
  XOR U2542 ( .A(n26216), .B(n26362), .Z(n26220) );
  XOR U2543 ( .A(n25194), .B(n25340), .Z(n25198) );
  XOR U2544 ( .A(n24146), .B(n24292), .Z(n24150) );
  XOR U2545 ( .A(n23077), .B(n23223), .Z(n23081) );
  XOR U2546 ( .A(n21984), .B(n22130), .Z(n21988) );
  XOR U2547 ( .A(n20867), .B(n21013), .Z(n20871) );
  XOR U2548 ( .A(n19727), .B(n19873), .Z(n19731) );
  XOR U2549 ( .A(n14189), .B(n14336), .Z(n14193) );
  XOR U2550 ( .A(n12915), .B(n13062), .Z(n12919) );
  XOR U2551 ( .A(n2356), .B(n2785), .Z(n2360) );
  XOR U2552 ( .A(n3875), .B(n4226), .Z(n3879) );
  XOR U2553 ( .A(n2401), .B(n2776), .Z(n2405) );
  XOR U2554 ( .A(n6088), .B(n6349), .Z(n6092) );
  XOR U2555 ( .A(n4648), .B(n4933), .Z(n4652) );
  XOR U2556 ( .A(n8245), .B(n8416), .Z(n8249) );
  XOR U2557 ( .A(n6843), .B(n7038), .Z(n6847) );
  XOR U2558 ( .A(n45668), .B(n45802), .Z(n45672) );
  XOR U2559 ( .A(n45368), .B(n45502), .Z(n45372) );
  XOR U2560 ( .A(n17877), .B(n18012), .Z(n17881) );
  XOR U2561 ( .A(n10303), .B(n10438), .Z(n10307) );
  XOR U2562 ( .A(n8275), .B(n8410), .Z(n8279) );
  XOR U2563 ( .A(n6873), .B(n7032), .Z(n6877) );
  XOR U2564 ( .A(n6118), .B(n6343), .Z(n6122) );
  XOR U2565 ( .A(n4678), .B(n4927), .Z(n4682) );
  XOR U2566 ( .A(n3905), .B(n4220), .Z(n3909) );
  XOR U2567 ( .A(n2431), .B(n2770), .Z(n2435) );
  XOR U2568 ( .A(n2386), .B(n2779), .Z(n2390) );
  XNOR U2569 ( .A(n45532), .B(n45376), .Z(n45378) );
  XOR U2570 ( .A(n45049), .B(n45177), .Z(n45053) );
  XOR U2571 ( .A(n44701), .B(n44829), .Z(n44705) );
  XOR U2572 ( .A(n44329), .B(n44457), .Z(n44333) );
  XOR U2573 ( .A(n43933), .B(n44061), .Z(n43937) );
  XOR U2574 ( .A(n43513), .B(n43641), .Z(n43517) );
  XOR U2575 ( .A(n43069), .B(n43197), .Z(n43073) );
  XOR U2576 ( .A(n42601), .B(n42729), .Z(n42605) );
  XOR U2577 ( .A(n42109), .B(n42237), .Z(n42113) );
  XOR U2578 ( .A(n41593), .B(n41721), .Z(n41597) );
  XOR U2579 ( .A(n41053), .B(n41181), .Z(n41057) );
  XOR U2580 ( .A(n40489), .B(n40617), .Z(n40493) );
  XOR U2581 ( .A(n39901), .B(n40029), .Z(n39905) );
  XOR U2582 ( .A(n39289), .B(n39417), .Z(n39293) );
  XOR U2583 ( .A(n38653), .B(n38781), .Z(n38657) );
  XOR U2584 ( .A(n37993), .B(n38121), .Z(n37997) );
  XOR U2585 ( .A(n37309), .B(n37437), .Z(n37313) );
  XOR U2586 ( .A(n36601), .B(n36729), .Z(n36605) );
  XOR U2587 ( .A(n35869), .B(n35997), .Z(n35873) );
  XOR U2588 ( .A(n35113), .B(n35241), .Z(n35117) );
  XOR U2589 ( .A(n34333), .B(n34461), .Z(n34337) );
  XOR U2590 ( .A(n33529), .B(n33657), .Z(n33533) );
  XOR U2591 ( .A(n32701), .B(n32829), .Z(n32705) );
  XOR U2592 ( .A(n31849), .B(n31977), .Z(n31853) );
  XOR U2593 ( .A(n30973), .B(n31101), .Z(n30977) );
  XOR U2594 ( .A(n30073), .B(n30201), .Z(n30077) );
  XOR U2595 ( .A(n29149), .B(n29277), .Z(n29153) );
  XOR U2596 ( .A(n28201), .B(n28329), .Z(n28205) );
  XOR U2597 ( .A(n27229), .B(n27357), .Z(n27233) );
  XOR U2598 ( .A(n26231), .B(n26359), .Z(n26235) );
  XOR U2599 ( .A(n25209), .B(n25337), .Z(n25213) );
  XOR U2600 ( .A(n24161), .B(n24289), .Z(n24165) );
  XOR U2601 ( .A(n23092), .B(n23220), .Z(n23096) );
  XOR U2602 ( .A(n21999), .B(n22127), .Z(n22003) );
  XOR U2603 ( .A(n20882), .B(n21010), .Z(n20886) );
  XOR U2604 ( .A(n19742), .B(n19870), .Z(n19746) );
  XOR U2605 ( .A(n15454), .B(n15583), .Z(n15458) );
  XOR U2606 ( .A(n14204), .B(n14333), .Z(n14208) );
  XOR U2607 ( .A(n12930), .B(n13059), .Z(n12934) );
  XOR U2608 ( .A(n9638), .B(n9767), .Z(n9642) );
  XOR U2609 ( .A(n2416), .B(n2773), .Z(n2420) );
  XOR U2610 ( .A(n3935), .B(n4214), .Z(n3939) );
  XOR U2611 ( .A(n2461), .B(n2764), .Z(n2465) );
  XOR U2612 ( .A(n6148), .B(n6337), .Z(n6152) );
  XOR U2613 ( .A(n4708), .B(n4921), .Z(n4712) );
  XOR U2614 ( .A(n16685), .B(n16808), .Z(n16689) );
  XOR U2615 ( .A(n12287), .B(n12412), .Z(n12291) );
  XOR U2616 ( .A(n46088), .B(n46204), .Z(n46092) );
  XOR U2617 ( .A(n45824), .B(n45940), .Z(n45828) );
  XOR U2618 ( .A(n17892), .B(n18009), .Z(n17896) );
  XOR U2619 ( .A(n8972), .B(n9089), .Z(n8976) );
  XOR U2620 ( .A(n7602), .B(n7719), .Z(n7606) );
  XOR U2621 ( .A(n6178), .B(n6331), .Z(n6182) );
  XOR U2622 ( .A(n4738), .B(n4915), .Z(n4742) );
  XOR U2623 ( .A(n3965), .B(n4208), .Z(n3969) );
  XOR U2624 ( .A(n2491), .B(n2758), .Z(n2495) );
  XOR U2625 ( .A(n2446), .B(n2767), .Z(n2450) );
  XOR U2626 ( .A(n45688), .B(n45798), .Z(n45692) );
  XOR U2627 ( .A(n45388), .B(n45498), .Z(n45392) );
  XOR U2628 ( .A(n45064), .B(n45174), .Z(n45068) );
  XOR U2629 ( .A(n44716), .B(n44826), .Z(n44720) );
  XOR U2630 ( .A(n44344), .B(n44454), .Z(n44348) );
  XOR U2631 ( .A(n43948), .B(n44058), .Z(n43952) );
  XOR U2632 ( .A(n43528), .B(n43638), .Z(n43532) );
  XOR U2633 ( .A(n43084), .B(n43194), .Z(n43088) );
  XOR U2634 ( .A(n42616), .B(n42726), .Z(n42620) );
  XOR U2635 ( .A(n42124), .B(n42234), .Z(n42128) );
  XOR U2636 ( .A(n41608), .B(n41718), .Z(n41612) );
  XOR U2637 ( .A(n41068), .B(n41178), .Z(n41072) );
  XOR U2638 ( .A(n40504), .B(n40614), .Z(n40508) );
  XOR U2639 ( .A(n39916), .B(n40026), .Z(n39920) );
  XOR U2640 ( .A(n39304), .B(n39414), .Z(n39308) );
  XOR U2641 ( .A(n38668), .B(n38778), .Z(n38672) );
  XOR U2642 ( .A(n38008), .B(n38118), .Z(n38012) );
  XOR U2643 ( .A(n37324), .B(n37434), .Z(n37328) );
  XOR U2644 ( .A(n36616), .B(n36726), .Z(n36620) );
  XOR U2645 ( .A(n35884), .B(n35994), .Z(n35888) );
  XOR U2646 ( .A(n35128), .B(n35238), .Z(n35132) );
  XOR U2647 ( .A(n34348), .B(n34458), .Z(n34352) );
  XOR U2648 ( .A(n33544), .B(n33654), .Z(n33548) );
  XOR U2649 ( .A(n32716), .B(n32826), .Z(n32720) );
  XOR U2650 ( .A(n31864), .B(n31974), .Z(n31868) );
  XOR U2651 ( .A(n30988), .B(n31098), .Z(n30992) );
  XOR U2652 ( .A(n30088), .B(n30198), .Z(n30092) );
  XOR U2653 ( .A(n29164), .B(n29274), .Z(n29168) );
  XOR U2654 ( .A(n28216), .B(n28326), .Z(n28220) );
  XOR U2655 ( .A(n27244), .B(n27354), .Z(n27248) );
  XOR U2656 ( .A(n26246), .B(n26356), .Z(n26250) );
  XOR U2657 ( .A(n25224), .B(n25334), .Z(n25228) );
  XOR U2658 ( .A(n24176), .B(n24286), .Z(n24180) );
  XOR U2659 ( .A(n23107), .B(n23217), .Z(n23111) );
  XOR U2660 ( .A(n22014), .B(n22124), .Z(n22018) );
  XOR U2661 ( .A(n20897), .B(n21007), .Z(n20901) );
  XOR U2662 ( .A(n19757), .B(n19867), .Z(n19761) );
  XOR U2663 ( .A(n16085), .B(n16196), .Z(n16089) );
  XOR U2664 ( .A(n2476), .B(n2761), .Z(n2480) );
  XOR U2665 ( .A(n3995), .B(n4202), .Z(n3999) );
  XOR U2666 ( .A(n2521), .B(n2752), .Z(n2525) );
  XOR U2667 ( .A(n6208), .B(n6325), .Z(n6212) );
  XOR U2668 ( .A(n4768), .B(n4909), .Z(n4772) );
  XOR U2669 ( .A(n17304), .B(n17409), .Z(n17308) );
  XOR U2670 ( .A(n14852), .B(n14957), .Z(n14856) );
  XOR U2671 ( .A(n12950), .B(n13055), .Z(n12954) );
  XOR U2672 ( .A(n10992), .B(n11097), .Z(n10996) );
  XOR U2673 ( .A(n46454), .B(n46552), .Z(n46458) );
  XOR U2674 ( .A(n46226), .B(n46324), .Z(n46230) );
  XOR U2675 ( .A(n18499), .B(n18619), .Z(n18503) );
  XOR U2676 ( .A(n10333), .B(n10432), .Z(n10337) );
  XOR U2677 ( .A(n8987), .B(n9086), .Z(n8991) );
  XOR U2678 ( .A(n7617), .B(n7716), .Z(n7621) );
  XOR U2679 ( .A(n4798), .B(n4903), .Z(n4802) );
  XOR U2680 ( .A(n4025), .B(n4196), .Z(n4029) );
  XOR U2681 ( .A(n2551), .B(n2746), .Z(n2555) );
  XOR U2682 ( .A(n2506), .B(n2755), .Z(n2510) );
  XNOR U2683 ( .A(n46354), .B(n46234), .Z(n46236) );
  XOR U2684 ( .A(n45979), .B(n46071), .Z(n45983) );
  XOR U2685 ( .A(n45703), .B(n45795), .Z(n45707) );
  XOR U2686 ( .A(n45403), .B(n45495), .Z(n45407) );
  XOR U2687 ( .A(n45079), .B(n45171), .Z(n45083) );
  XOR U2688 ( .A(n44731), .B(n44823), .Z(n44735) );
  XOR U2689 ( .A(n44359), .B(n44451), .Z(n44363) );
  XOR U2690 ( .A(n43963), .B(n44055), .Z(n43967) );
  XOR U2691 ( .A(n43543), .B(n43635), .Z(n43547) );
  XOR U2692 ( .A(n43099), .B(n43191), .Z(n43103) );
  XOR U2693 ( .A(n42631), .B(n42723), .Z(n42635) );
  XOR U2694 ( .A(n42139), .B(n42231), .Z(n42143) );
  XOR U2695 ( .A(n41623), .B(n41715), .Z(n41627) );
  XOR U2696 ( .A(n41083), .B(n41175), .Z(n41087) );
  XOR U2697 ( .A(n40519), .B(n40611), .Z(n40523) );
  XOR U2698 ( .A(n39931), .B(n40023), .Z(n39935) );
  XOR U2699 ( .A(n39319), .B(n39411), .Z(n39323) );
  XOR U2700 ( .A(n38683), .B(n38775), .Z(n38687) );
  XOR U2701 ( .A(n38023), .B(n38115), .Z(n38027) );
  XOR U2702 ( .A(n37339), .B(n37431), .Z(n37343) );
  XOR U2703 ( .A(n36631), .B(n36723), .Z(n36635) );
  XOR U2704 ( .A(n35899), .B(n35991), .Z(n35903) );
  XOR U2705 ( .A(n35143), .B(n35235), .Z(n35147) );
  XOR U2706 ( .A(n34363), .B(n34455), .Z(n34367) );
  XOR U2707 ( .A(n33559), .B(n33651), .Z(n33563) );
  XOR U2708 ( .A(n32731), .B(n32823), .Z(n32735) );
  XOR U2709 ( .A(n31879), .B(n31971), .Z(n31883) );
  XOR U2710 ( .A(n31003), .B(n31095), .Z(n31007) );
  XOR U2711 ( .A(n30103), .B(n30195), .Z(n30107) );
  XOR U2712 ( .A(n29179), .B(n29271), .Z(n29183) );
  XOR U2713 ( .A(n28231), .B(n28323), .Z(n28235) );
  XOR U2714 ( .A(n27259), .B(n27351), .Z(n27263) );
  XOR U2715 ( .A(n26261), .B(n26353), .Z(n26265) );
  XOR U2716 ( .A(n25239), .B(n25331), .Z(n25243) );
  XOR U2717 ( .A(n24191), .B(n24283), .Z(n24195) );
  XOR U2718 ( .A(n23122), .B(n23214), .Z(n23126) );
  XOR U2719 ( .A(n22029), .B(n22121), .Z(n22033) );
  XOR U2720 ( .A(n20912), .B(n21004), .Z(n20916) );
  XOR U2721 ( .A(n19772), .B(n19864), .Z(n19776) );
  XOR U2722 ( .A(n2536), .B(n2749), .Z(n2540) );
  XOR U2723 ( .A(n4055), .B(n4190), .Z(n4059) );
  XOR U2724 ( .A(n2581), .B(n2740), .Z(n2585) );
  XOR U2725 ( .A(n17917), .B(n18004), .Z(n17921) );
  XOR U2726 ( .A(n16715), .B(n16802), .Z(n16719) );
  XOR U2727 ( .A(n15489), .B(n15576), .Z(n15493) );
  XOR U2728 ( .A(n14239), .B(n14326), .Z(n14243) );
  XOR U2729 ( .A(n12965), .B(n13052), .Z(n12969) );
  XOR U2730 ( .A(n46766), .B(n46846), .Z(n46770) );
  XOR U2731 ( .A(n46574), .B(n46654), .Z(n46578) );
  XOR U2732 ( .A(n12322), .B(n12405), .Z(n12326) );
  XOR U2733 ( .A(n11012), .B(n11093), .Z(n11016) );
  XOR U2734 ( .A(n9678), .B(n9759), .Z(n9682) );
  XOR U2735 ( .A(n8320), .B(n8401), .Z(n8324) );
  XOR U2736 ( .A(n6938), .B(n7019), .Z(n6942) );
  XOR U2737 ( .A(n5530), .B(n5613), .Z(n5534) );
  XOR U2738 ( .A(n4085), .B(n4184), .Z(n4089) );
  XOR U2739 ( .A(n2611), .B(n2734), .Z(n2615) );
  XOR U2740 ( .A(n2566), .B(n2743), .Z(n2570) );
  XOR U2741 ( .A(n46474), .B(n46548), .Z(n46478) );
  XOR U2742 ( .A(n46246), .B(n46320), .Z(n46250) );
  XOR U2743 ( .A(n45994), .B(n46068), .Z(n45998) );
  XOR U2744 ( .A(n45718), .B(n45792), .Z(n45722) );
  XOR U2745 ( .A(n45418), .B(n45492), .Z(n45422) );
  XOR U2746 ( .A(n45094), .B(n45168), .Z(n45098) );
  XOR U2747 ( .A(n44746), .B(n44820), .Z(n44750) );
  XOR U2748 ( .A(n44374), .B(n44448), .Z(n44378) );
  XOR U2749 ( .A(n43978), .B(n44052), .Z(n43982) );
  XOR U2750 ( .A(n43558), .B(n43632), .Z(n43562) );
  XOR U2751 ( .A(n43114), .B(n43188), .Z(n43118) );
  XOR U2752 ( .A(n42646), .B(n42720), .Z(n42650) );
  XOR U2753 ( .A(n42154), .B(n42228), .Z(n42158) );
  XOR U2754 ( .A(n41638), .B(n41712), .Z(n41642) );
  XOR U2755 ( .A(n41098), .B(n41172), .Z(n41102) );
  XOR U2756 ( .A(n40534), .B(n40608), .Z(n40538) );
  XOR U2757 ( .A(n39946), .B(n40020), .Z(n39950) );
  XOR U2758 ( .A(n39334), .B(n39408), .Z(n39338) );
  XOR U2759 ( .A(n38698), .B(n38772), .Z(n38702) );
  XOR U2760 ( .A(n38038), .B(n38112), .Z(n38042) );
  XOR U2761 ( .A(n37354), .B(n37428), .Z(n37358) );
  XOR U2762 ( .A(n36646), .B(n36720), .Z(n36650) );
  XOR U2763 ( .A(n35914), .B(n35988), .Z(n35918) );
  XOR U2764 ( .A(n35158), .B(n35232), .Z(n35162) );
  XOR U2765 ( .A(n34378), .B(n34452), .Z(n34382) );
  XOR U2766 ( .A(n33574), .B(n33648), .Z(n33578) );
  XOR U2767 ( .A(n32746), .B(n32820), .Z(n32750) );
  XOR U2768 ( .A(n31894), .B(n31968), .Z(n31898) );
  XOR U2769 ( .A(n31018), .B(n31092), .Z(n31022) );
  XOR U2770 ( .A(n30118), .B(n30192), .Z(n30122) );
  XOR U2771 ( .A(n29194), .B(n29268), .Z(n29198) );
  XOR U2772 ( .A(n28246), .B(n28320), .Z(n28250) );
  XOR U2773 ( .A(n27274), .B(n27348), .Z(n27278) );
  XOR U2774 ( .A(n26276), .B(n26350), .Z(n26280) );
  XOR U2775 ( .A(n25254), .B(n25328), .Z(n25258) );
  XOR U2776 ( .A(n24206), .B(n24280), .Z(n24210) );
  XOR U2777 ( .A(n23137), .B(n23211), .Z(n23141) );
  XOR U2778 ( .A(n22044), .B(n22118), .Z(n22048) );
  XOR U2779 ( .A(n20927), .B(n21001), .Z(n20931) );
  XOR U2780 ( .A(n19787), .B(n19861), .Z(n19791) );
  XOR U2781 ( .A(n2596), .B(n2737), .Z(n2600) );
  XOR U2782 ( .A(n17932), .B(n18001), .Z(n17936) );
  XOR U2783 ( .A(n16730), .B(n16799), .Z(n16734) );
  XOR U2784 ( .A(n15504), .B(n15573), .Z(n15508) );
  XOR U2785 ( .A(n14254), .B(n14323), .Z(n14258) );
  XOR U2786 ( .A(n4110), .B(n4179), .Z(n4114) );
  XOR U2787 ( .A(n47024), .B(n47086), .Z(n47028) );
  XOR U2788 ( .A(n46868), .B(n46930), .Z(n46872) );
  XOR U2789 ( .A(n13625), .B(n13688), .Z(n13629) );
  XOR U2790 ( .A(n12337), .B(n12402), .Z(n12341) );
  XOR U2791 ( .A(n11027), .B(n11090), .Z(n11031) );
  XOR U2792 ( .A(n9693), .B(n9756), .Z(n9697) );
  XOR U2793 ( .A(n8335), .B(n8398), .Z(n8339) );
  XOR U2794 ( .A(n6953), .B(n7016), .Z(n6957) );
  XOR U2795 ( .A(n5545), .B(n5610), .Z(n5549) );
  XOR U2796 ( .A(n2626), .B(n2731), .Z(n2630) );
  XOR U2797 ( .A(n3391), .B(n3454), .Z(n3395) );
  XNOR U2798 ( .A(n46960), .B(n46876), .Z(n46878) );
  XOR U2799 ( .A(n46693), .B(n46749), .Z(n46697) );
  XOR U2800 ( .A(n46489), .B(n46545), .Z(n46493) );
  XOR U2801 ( .A(n46261), .B(n46317), .Z(n46265) );
  XOR U2802 ( .A(n46009), .B(n46065), .Z(n46013) );
  XOR U2803 ( .A(n45733), .B(n45789), .Z(n45737) );
  XOR U2804 ( .A(n45433), .B(n45489), .Z(n45437) );
  XOR U2805 ( .A(n45109), .B(n45165), .Z(n45113) );
  XOR U2806 ( .A(n44761), .B(n44817), .Z(n44765) );
  XOR U2807 ( .A(n44389), .B(n44445), .Z(n44393) );
  XOR U2808 ( .A(n43993), .B(n44049), .Z(n43997) );
  XOR U2809 ( .A(n43573), .B(n43629), .Z(n43577) );
  XOR U2810 ( .A(n43129), .B(n43185), .Z(n43133) );
  XOR U2811 ( .A(n42661), .B(n42717), .Z(n42665) );
  XOR U2812 ( .A(n42169), .B(n42225), .Z(n42173) );
  XOR U2813 ( .A(n41653), .B(n41709), .Z(n41657) );
  XOR U2814 ( .A(n41113), .B(n41169), .Z(n41117) );
  XOR U2815 ( .A(n40549), .B(n40605), .Z(n40553) );
  XOR U2816 ( .A(n39961), .B(n40017), .Z(n39965) );
  XOR U2817 ( .A(n39349), .B(n39405), .Z(n39353) );
  XOR U2818 ( .A(n38713), .B(n38769), .Z(n38717) );
  XOR U2819 ( .A(n38053), .B(n38109), .Z(n38057) );
  XOR U2820 ( .A(n37369), .B(n37425), .Z(n37373) );
  XOR U2821 ( .A(n36661), .B(n36717), .Z(n36665) );
  XOR U2822 ( .A(n35929), .B(n35985), .Z(n35933) );
  XOR U2823 ( .A(n35173), .B(n35229), .Z(n35177) );
  XOR U2824 ( .A(n34393), .B(n34449), .Z(n34397) );
  XOR U2825 ( .A(n33589), .B(n33645), .Z(n33593) );
  XOR U2826 ( .A(n32761), .B(n32817), .Z(n32765) );
  XOR U2827 ( .A(n31909), .B(n31965), .Z(n31913) );
  XOR U2828 ( .A(n31033), .B(n31089), .Z(n31037) );
  XOR U2829 ( .A(n30133), .B(n30189), .Z(n30137) );
  XOR U2830 ( .A(n29209), .B(n29265), .Z(n29213) );
  XOR U2831 ( .A(n28261), .B(n28317), .Z(n28265) );
  XOR U2832 ( .A(n27289), .B(n27345), .Z(n27293) );
  XOR U2833 ( .A(n26291), .B(n26347), .Z(n26295) );
  XOR U2834 ( .A(n25269), .B(n25325), .Z(n25273) );
  XOR U2835 ( .A(n24221), .B(n24277), .Z(n24225) );
  XOR U2836 ( .A(n23152), .B(n23208), .Z(n23156) );
  XOR U2837 ( .A(n22059), .B(n22115), .Z(n22063) );
  XOR U2838 ( .A(n20942), .B(n20998), .Z(n20946) );
  XOR U2839 ( .A(n19802), .B(n19858), .Z(n19806) );
  XOR U2840 ( .A(n17947), .B(n17998), .Z(n17951) );
  XOR U2841 ( .A(n15519), .B(n15570), .Z(n15523) );
  XOR U2842 ( .A(n47227), .B(n47271), .Z(n47231) );
  XOR U2843 ( .A(n47108), .B(n47152), .Z(n47112) );
  XOR U2844 ( .A(n14902), .B(n14947), .Z(n14906) );
  XOR U2845 ( .A(n13640), .B(n13685), .Z(n13644) );
  XOR U2846 ( .A(n12352), .B(n12399), .Z(n12356) );
  XOR U2847 ( .A(n11042), .B(n11087), .Z(n11046) );
  XOR U2848 ( .A(n9708), .B(n9753), .Z(n9712) );
  XOR U2849 ( .A(n8350), .B(n8395), .Z(n8354) );
  XOR U2850 ( .A(n6968), .B(n7013), .Z(n6972) );
  XOR U2851 ( .A(n5560), .B(n5607), .Z(n5564) );
  XOR U2852 ( .A(n4130), .B(n4175), .Z(n4134) );
  XOR U2853 ( .A(n2676), .B(n2721), .Z(n2680) );
  XOR U2854 ( .A(n47328), .B(n47366), .Z(n47332) );
  XOR U2855 ( .A(n47044), .B(n47082), .Z(n47048) );
  XOR U2856 ( .A(n46888), .B(n46926), .Z(n46892) );
  XOR U2857 ( .A(n46708), .B(n46746), .Z(n46712) );
  XOR U2858 ( .A(n46504), .B(n46542), .Z(n46508) );
  XOR U2859 ( .A(n46276), .B(n46314), .Z(n46280) );
  XOR U2860 ( .A(n46024), .B(n46062), .Z(n46028) );
  XOR U2861 ( .A(n45748), .B(n45786), .Z(n45752) );
  XOR U2862 ( .A(n45448), .B(n45486), .Z(n45452) );
  XOR U2863 ( .A(n45124), .B(n45162), .Z(n45128) );
  XOR U2864 ( .A(n44776), .B(n44814), .Z(n44780) );
  XOR U2865 ( .A(n44404), .B(n44442), .Z(n44408) );
  XOR U2866 ( .A(n44008), .B(n44046), .Z(n44012) );
  XOR U2867 ( .A(n43588), .B(n43626), .Z(n43592) );
  XOR U2868 ( .A(n43144), .B(n43182), .Z(n43148) );
  XOR U2869 ( .A(n42676), .B(n42714), .Z(n42680) );
  XOR U2870 ( .A(n42184), .B(n42222), .Z(n42188) );
  XOR U2871 ( .A(n41668), .B(n41706), .Z(n41672) );
  XOR U2872 ( .A(n41128), .B(n41166), .Z(n41132) );
  XOR U2873 ( .A(n40564), .B(n40602), .Z(n40568) );
  XOR U2874 ( .A(n39976), .B(n40014), .Z(n39980) );
  XOR U2875 ( .A(n39364), .B(n39402), .Z(n39368) );
  XOR U2876 ( .A(n38728), .B(n38766), .Z(n38732) );
  XOR U2877 ( .A(n38068), .B(n38106), .Z(n38072) );
  XOR U2878 ( .A(n37384), .B(n37422), .Z(n37388) );
  XOR U2879 ( .A(n36676), .B(n36714), .Z(n36680) );
  XOR U2880 ( .A(n35944), .B(n35982), .Z(n35948) );
  XOR U2881 ( .A(n35188), .B(n35226), .Z(n35192) );
  XOR U2882 ( .A(n34408), .B(n34446), .Z(n34412) );
  XOR U2883 ( .A(n33604), .B(n33642), .Z(n33608) );
  XOR U2884 ( .A(n32776), .B(n32814), .Z(n32780) );
  XOR U2885 ( .A(n31924), .B(n31962), .Z(n31928) );
  XOR U2886 ( .A(n31048), .B(n31086), .Z(n31052) );
  XOR U2887 ( .A(n30148), .B(n30186), .Z(n30152) );
  XOR U2888 ( .A(n29224), .B(n29262), .Z(n29228) );
  XOR U2889 ( .A(n28276), .B(n28314), .Z(n28280) );
  XOR U2890 ( .A(n27304), .B(n27342), .Z(n27308) );
  XOR U2891 ( .A(n26306), .B(n26344), .Z(n26310) );
  XOR U2892 ( .A(n25284), .B(n25322), .Z(n25288) );
  XOR U2893 ( .A(n24236), .B(n24274), .Z(n24240) );
  XOR U2894 ( .A(n23167), .B(n23205), .Z(n23171) );
  XOR U2895 ( .A(n22074), .B(n22112), .Z(n22078) );
  XOR U2896 ( .A(n20957), .B(n20995), .Z(n20961) );
  XOR U2897 ( .A(n19817), .B(n19855), .Z(n19821) );
  XOR U2898 ( .A(n16760), .B(n16793), .Z(n16764) );
  XOR U2899 ( .A(n47293), .B(n47319), .Z(n47297) );
  XOR U2900 ( .A(n17967), .B(n17994), .Z(n17971) );
  XOR U2901 ( .A(n16155), .B(n16182), .Z(n16159) );
  XOR U2902 ( .A(n14917), .B(n14944), .Z(n14921) );
  XOR U2903 ( .A(n13655), .B(n13682), .Z(n13659) );
  XOR U2904 ( .A(n12367), .B(n12396), .Z(n12371) );
  XOR U2905 ( .A(n11057), .B(n11084), .Z(n11061) );
  XOR U2906 ( .A(n9723), .B(n9750), .Z(n9727) );
  XOR U2907 ( .A(n8365), .B(n8392), .Z(n8369) );
  XOR U2908 ( .A(n6983), .B(n7010), .Z(n6987) );
  XOR U2909 ( .A(n5575), .B(n5604), .Z(n5579) );
  XOR U2910 ( .A(n4145), .B(n4172), .Z(n4149) );
  XOR U2911 ( .A(n2691), .B(n2718), .Z(n2695) );
  XOR U2912 ( .A(n47442), .B(n47462), .Z(n47446) );
  XOR U2913 ( .A(n47382), .B(n47402), .Z(n47386) );
  XOR U2914 ( .A(n47247), .B(n47267), .Z(n47251) );
  XOR U2915 ( .A(n47128), .B(n47148), .Z(n47132) );
  XOR U2916 ( .A(n46984), .B(n47004), .Z(n46988) );
  XOR U2917 ( .A(n46816), .B(n46836), .Z(n46820) );
  XOR U2918 ( .A(n46624), .B(n46644), .Z(n46628) );
  XOR U2919 ( .A(n46408), .B(n46428), .Z(n46412) );
  XOR U2920 ( .A(n46168), .B(n46188), .Z(n46172) );
  XOR U2921 ( .A(n45904), .B(n45924), .Z(n45908) );
  XOR U2922 ( .A(n45616), .B(n45636), .Z(n45620) );
  XOR U2923 ( .A(n45304), .B(n45324), .Z(n45308) );
  XOR U2924 ( .A(n44968), .B(n44988), .Z(n44972) );
  XOR U2925 ( .A(n44608), .B(n44628), .Z(n44612) );
  XOR U2926 ( .A(n44224), .B(n44244), .Z(n44228) );
  XOR U2927 ( .A(n43816), .B(n43836), .Z(n43820) );
  XOR U2928 ( .A(n43384), .B(n43404), .Z(n43388) );
  XOR U2929 ( .A(n42928), .B(n42948), .Z(n42932) );
  XOR U2930 ( .A(n42448), .B(n42468), .Z(n42452) );
  XOR U2931 ( .A(n41944), .B(n41964), .Z(n41948) );
  XOR U2932 ( .A(n41416), .B(n41436), .Z(n41420) );
  XOR U2933 ( .A(n40864), .B(n40884), .Z(n40868) );
  XOR U2934 ( .A(n40288), .B(n40308), .Z(n40292) );
  XOR U2935 ( .A(n39688), .B(n39708), .Z(n39692) );
  XOR U2936 ( .A(n39064), .B(n39084), .Z(n39068) );
  XOR U2937 ( .A(n38416), .B(n38436), .Z(n38420) );
  XOR U2938 ( .A(n37744), .B(n37764), .Z(n37748) );
  XOR U2939 ( .A(n37048), .B(n37068), .Z(n37052) );
  XOR U2940 ( .A(n36328), .B(n36348), .Z(n36332) );
  XOR U2941 ( .A(n35584), .B(n35604), .Z(n35588) );
  XOR U2942 ( .A(n34816), .B(n34836), .Z(n34820) );
  XOR U2943 ( .A(n34024), .B(n34044), .Z(n34028) );
  XOR U2944 ( .A(n33208), .B(n33228), .Z(n33212) );
  XOR U2945 ( .A(n32368), .B(n32388), .Z(n32372) );
  XOR U2946 ( .A(n31504), .B(n31524), .Z(n31508) );
  XOR U2947 ( .A(n30616), .B(n30636), .Z(n30620) );
  XOR U2948 ( .A(n29704), .B(n29724), .Z(n29708) );
  XOR U2949 ( .A(n28768), .B(n28788), .Z(n28772) );
  XOR U2950 ( .A(n27808), .B(n27828), .Z(n27812) );
  XOR U2951 ( .A(n26822), .B(n26842), .Z(n26826) );
  XOR U2952 ( .A(n25813), .B(n25833), .Z(n25817) );
  XOR U2953 ( .A(n24776), .B(n24796), .Z(n24780) );
  XOR U2954 ( .A(n23720), .B(n23740), .Z(n23724) );
  XOR U2955 ( .A(n22638), .B(n22658), .Z(n22642) );
  XOR U2956 ( .A(n21534), .B(n21554), .Z(n21538) );
  XOR U2957 ( .A(n20405), .B(n20425), .Z(n20409) );
  XOR U2958 ( .A(n19253), .B(n19273), .Z(n19257) );
  XNOR U2959 ( .A(n28870), .B(n28396), .Z(n28398) );
  XNOR U2960 ( .A(n28399), .B(n27919), .Z(n27921) );
  XOR U2961 ( .A(n26944), .B(n27414), .Z(n26948) );
  XOR U2962 ( .A(n25926), .B(n26420), .Z(n25930) );
  XNOR U2963 ( .A(n30262), .B(n29806), .Z(n29808) );
  XNOR U2964 ( .A(n29809), .B(n29347), .Z(n29349) );
  XNOR U2965 ( .A(n29350), .B(n28882), .Z(n28884) );
  XNOR U2966 ( .A(n28885), .B(n28411), .Z(n28413) );
  XNOR U2967 ( .A(n28414), .B(n27934), .Z(n27936) );
  XOR U2968 ( .A(n26959), .B(n27411), .Z(n26963) );
  XOR U2969 ( .A(n25438), .B(n25909), .Z(n25442) );
  XOR U2970 ( .A(n25961), .B(n26413), .Z(n25965) );
  XOR U2971 ( .A(n25941), .B(n26417), .Z(n25945) );
  XOR U2972 ( .A(n24898), .B(n25400), .Z(n24902) );
  XNOR U2973 ( .A(n31600), .B(n31162), .Z(n31164) );
  XNOR U2974 ( .A(n31165), .B(n30721), .Z(n30723) );
  XNOR U2975 ( .A(n30724), .B(n30274), .Z(n30276) );
  XNOR U2976 ( .A(n30277), .B(n29821), .Z(n29823) );
  XOR U2977 ( .A(n28894), .B(n29328), .Z(n28898) );
  XOR U2978 ( .A(n27946), .B(n28380), .Z(n27950) );
  XOR U2979 ( .A(n26974), .B(n27408), .Z(n26978) );
  XOR U2980 ( .A(n23836), .B(n24354), .Z(n23840) );
  XOR U2981 ( .A(n24948), .B(n25390), .Z(n24952) );
  XOR U2982 ( .A(n23861), .B(n24349), .Z(n23865) );
  XNOR U2983 ( .A(n23296), .B(n22755), .Z(n22757) );
  XOR U2984 ( .A(n25458), .B(n25905), .Z(n25462) );
  XOR U2985 ( .A(n24401), .B(n24874), .Z(n24405) );
  XOR U2986 ( .A(n24381), .B(n24878), .Z(n24385) );
  XNOR U2987 ( .A(n32884), .B(n32464), .Z(n32466) );
  XNOR U2988 ( .A(n32467), .B(n32041), .Z(n32043) );
  XNOR U2989 ( .A(n32044), .B(n31612), .Z(n31614) );
  XNOR U2990 ( .A(n31615), .B(n31177), .Z(n31179) );
  XNOR U2991 ( .A(n31180), .B(n30736), .Z(n30738) );
  XOR U2992 ( .A(n29833), .B(n30249), .Z(n29837) );
  XOR U2993 ( .A(n28909), .B(n29325), .Z(n28913) );
  XOR U2994 ( .A(n27961), .B(n28377), .Z(n27965) );
  XOR U2995 ( .A(n26989), .B(n27405), .Z(n26993) );
  XOR U2996 ( .A(n25991), .B(n26407), .Z(n25995) );
  XNOR U2997 ( .A(n24974), .B(n24449), .Z(n24451) );
  XOR U2998 ( .A(n23310), .B(n23822), .Z(n23314) );
  XNOR U2999 ( .A(n25484), .B(n24966), .Z(n24968) );
  XOR U3000 ( .A(n23896), .B(n24342), .Z(n23900) );
  XOR U3001 ( .A(n22787), .B(n23282), .Z(n22791) );
  XOR U3002 ( .A(n22213), .B(n22744), .Z(n22217) );
  XNOR U3003 ( .A(n21650), .B(n21092), .Z(n21094) );
  XOR U3004 ( .A(n22812), .B(n23277), .Z(n22816) );
  XOR U3005 ( .A(n23881), .B(n24345), .Z(n23885) );
  XNOR U3006 ( .A(n34114), .B(n33712), .Z(n33714) );
  XNOR U3007 ( .A(n33715), .B(n33307), .Z(n33309) );
  XNOR U3008 ( .A(n33310), .B(n32896), .Z(n32898) );
  XNOR U3009 ( .A(n32899), .B(n32479), .Z(n32481) );
  XOR U3010 ( .A(n31624), .B(n32022), .Z(n31628) );
  XOR U3011 ( .A(n30748), .B(n31146), .Z(n30752) );
  XOR U3012 ( .A(n29848), .B(n30246), .Z(n29852) );
  XOR U3013 ( .A(n28924), .B(n29322), .Z(n28928) );
  XOR U3014 ( .A(n27976), .B(n28374), .Z(n27980) );
  XOR U3015 ( .A(n27004), .B(n27402), .Z(n27008) );
  XOR U3016 ( .A(n26006), .B(n26404), .Z(n26010) );
  XOR U3017 ( .A(n24983), .B(n25382), .Z(n24987) );
  XOR U3018 ( .A(n23911), .B(n24339), .Z(n23915) );
  XOR U3019 ( .A(n23395), .B(n23805), .Z(n23399) );
  XOR U3020 ( .A(n21689), .B(n22189), .Z(n21693) );
  XOR U3021 ( .A(n20552), .B(n21077), .Z(n20556) );
  XOR U3022 ( .A(n21669), .B(n22193), .Z(n21673) );
  XNOR U3023 ( .A(n19951), .B(n19375), .Z(n19377) );
  XOR U3024 ( .A(n22827), .B(n23274), .Z(n22831) );
  XOR U3025 ( .A(n20577), .B(n21072), .Z(n20581) );
  XOR U3026 ( .A(n22298), .B(n22727), .Z(n22302) );
  XOR U3027 ( .A(n22253), .B(n22736), .Z(n22257) );
  XOR U3028 ( .A(n20537), .B(n21080), .Z(n20541) );
  XNOR U3029 ( .A(n19956), .B(n19380), .Z(n19382) );
  XOR U3030 ( .A(n21154), .B(n21630), .Z(n21158) );
  XNOR U3031 ( .A(n35290), .B(n34906), .Z(n34908) );
  XNOR U3032 ( .A(n34909), .B(n34519), .Z(n34521) );
  XNOR U3033 ( .A(n34522), .B(n34126), .Z(n34128) );
  XNOR U3034 ( .A(n34129), .B(n33727), .Z(n33729) );
  XNOR U3035 ( .A(n33730), .B(n33322), .Z(n33324) );
  XOR U3036 ( .A(n32491), .B(n32871), .Z(n32495) );
  XOR U3037 ( .A(n31639), .B(n32019), .Z(n31643) );
  XOR U3038 ( .A(n30763), .B(n31143), .Z(n30767) );
  XOR U3039 ( .A(n29863), .B(n30243), .Z(n29867) );
  XOR U3040 ( .A(n28939), .B(n29319), .Z(n28943) );
  XOR U3041 ( .A(n27991), .B(n28371), .Z(n27995) );
  XOR U3042 ( .A(n27019), .B(n27399), .Z(n27023) );
  XOR U3043 ( .A(n26021), .B(n26401), .Z(n26025) );
  XOR U3044 ( .A(n24999), .B(n25379), .Z(n25003) );
  XOR U3045 ( .A(n24476), .B(n24856), .Z(n24480) );
  XOR U3046 ( .A(n23420), .B(n23800), .Z(n23424) );
  XOR U3047 ( .A(n21179), .B(n21625), .Z(n21183) );
  XNOR U3048 ( .A(n21695), .B(n21137), .Z(n21139) );
  XOR U3049 ( .A(n19990), .B(n20508), .Z(n19994) );
  XOR U3050 ( .A(n21729), .B(n22181), .Z(n21733) );
  XNOR U3051 ( .A(n20011), .B(n19435), .Z(n19437) );
  XOR U3052 ( .A(n22333), .B(n22720), .Z(n22337) );
  XOR U3053 ( .A(n21209), .B(n21619), .Z(n21213) );
  XOR U3054 ( .A(n22313), .B(n22724), .Z(n22317) );
  XOR U3055 ( .A(n18823), .B(n19359), .Z(n18827) );
  XOR U3056 ( .A(n19392), .B(n19940), .Z(n19396) );
  XOR U3057 ( .A(n20597), .B(n21068), .Z(n20601) );
  XNOR U3058 ( .A(n20016), .B(n19440), .Z(n19442) );
  XNOR U3059 ( .A(n36412), .B(n36046), .Z(n36048) );
  XNOR U3060 ( .A(n36049), .B(n35677), .Z(n35679) );
  XNOR U3061 ( .A(n35680), .B(n35302), .Z(n35304) );
  XNOR U3062 ( .A(n35305), .B(n34921), .Z(n34923) );
  XOR U3063 ( .A(n34138), .B(n34500), .Z(n34142) );
  XOR U3064 ( .A(n33334), .B(n33696), .Z(n33338) );
  XOR U3065 ( .A(n32506), .B(n32868), .Z(n32510) );
  XOR U3066 ( .A(n31654), .B(n32016), .Z(n31658) );
  XOR U3067 ( .A(n30778), .B(n31140), .Z(n30782) );
  XOR U3068 ( .A(n29878), .B(n30240), .Z(n29882) );
  XOR U3069 ( .A(n28954), .B(n29316), .Z(n28958) );
  XOR U3070 ( .A(n28006), .B(n28368), .Z(n28010) );
  XOR U3071 ( .A(n27034), .B(n27396), .Z(n27038) );
  XOR U3072 ( .A(n26036), .B(n26398), .Z(n26040) );
  XOR U3073 ( .A(n25014), .B(n25376), .Z(n25018) );
  XOR U3074 ( .A(n23966), .B(n24328), .Z(n23970) );
  XOR U3075 ( .A(n23435), .B(n23797), .Z(n23439) );
  XOR U3076 ( .A(n22897), .B(n23259), .Z(n22901) );
  XOR U3077 ( .A(n21239), .B(n21613), .Z(n21243) );
  XNOR U3078 ( .A(n21755), .B(n21197), .Z(n21199) );
  XOR U3079 ( .A(n20622), .B(n21063), .Z(n20626) );
  XOR U3080 ( .A(n17522), .B(n18083), .Z(n17526) );
  XOR U3081 ( .A(n18104), .B(n18777), .Z(n18108) );
  XOR U3082 ( .A(n18149), .B(n18759), .Z(n18153) );
  XOR U3083 ( .A(n19467), .B(n19925), .Z(n19471) );
  XOR U3084 ( .A(n19422), .B(n19934), .Z(n19426) );
  XOR U3085 ( .A(n21789), .B(n22169), .Z(n21793) );
  XOR U3086 ( .A(n20075), .B(n20491), .Z(n20079) );
  XOR U3087 ( .A(n18134), .B(n18765), .Z(n18138) );
  XOR U3088 ( .A(n19452), .B(n19928), .Z(n19456) );
  XOR U3089 ( .A(n20657), .B(n21056), .Z(n20661) );
  XOR U3090 ( .A(n18908), .B(n19342), .Z(n18912) );
  XNOR U3091 ( .A(n37480), .B(n37132), .Z(n37134) );
  XNOR U3092 ( .A(n37135), .B(n36781), .Z(n36783) );
  XNOR U3093 ( .A(n36784), .B(n36424), .Z(n36426) );
  XNOR U3094 ( .A(n36427), .B(n36061), .Z(n36063) );
  XOR U3095 ( .A(n35314), .B(n35658), .Z(n35318) );
  XOR U3096 ( .A(n34546), .B(n34890), .Z(n34550) );
  XOR U3097 ( .A(n33754), .B(n34098), .Z(n33758) );
  XOR U3098 ( .A(n32938), .B(n33282), .Z(n32942) );
  XOR U3099 ( .A(n32098), .B(n32442), .Z(n32102) );
  XOR U3100 ( .A(n31234), .B(n31578), .Z(n31238) );
  XOR U3101 ( .A(n30346), .B(n30690), .Z(n30350) );
  XOR U3102 ( .A(n29434), .B(n29778), .Z(n29438) );
  XOR U3103 ( .A(n28498), .B(n28842), .Z(n28502) );
  XOR U3104 ( .A(n27538), .B(n27882), .Z(n27542) );
  XOR U3105 ( .A(n26552), .B(n26896), .Z(n26556) );
  XOR U3106 ( .A(n25543), .B(n25887), .Z(n25547) );
  XOR U3107 ( .A(n24506), .B(n24850), .Z(n24510) );
  XOR U3108 ( .A(n23450), .B(n23794), .Z(n23454) );
  XOR U3109 ( .A(n22368), .B(n22712), .Z(n22372) );
  XNOR U3110 ( .A(n22374), .B(n21822), .Z(n21824) );
  XOR U3111 ( .A(n20105), .B(n20485), .Z(n20109) );
  XOR U3112 ( .A(n20060), .B(n20494), .Z(n20064) );
  XOR U3113 ( .A(n17582), .B(n18071), .Z(n17586) );
  XOR U3114 ( .A(n15695), .B(n16274), .Z(n15699) );
  XOR U3115 ( .A(n16295), .B(n16886), .Z(n16299) );
  XOR U3116 ( .A(n18164), .B(n18753), .Z(n18168) );
  XOR U3117 ( .A(n16340), .B(n16877), .Z(n16344) );
  XOR U3118 ( .A(n20687), .B(n21050), .Z(n20691) );
  XOR U3119 ( .A(n18938), .B(n19336), .Z(n18942) );
  XOR U3120 ( .A(n18893), .B(n19345), .Z(n18897) );
  XOR U3121 ( .A(n17612), .B(n18065), .Z(n17616) );
  XOR U3122 ( .A(n20135), .B(n20479), .Z(n20139) );
  XOR U3123 ( .A(n16325), .B(n16880), .Z(n16329) );
  XOR U3124 ( .A(n19512), .B(n19916), .Z(n19516) );
  XOR U3125 ( .A(n18968), .B(n19330), .Z(n18972) );
  XNOR U3126 ( .A(n38494), .B(n38164), .Z(n38166) );
  XNOR U3127 ( .A(n38167), .B(n37831), .Z(n37833) );
  XNOR U3128 ( .A(n37834), .B(n37492), .Z(n37494) );
  XNOR U3129 ( .A(n37495), .B(n37147), .Z(n37149) );
  XNOR U3130 ( .A(n37150), .B(n36796), .Z(n36798) );
  XOR U3131 ( .A(n36073), .B(n36399), .Z(n36077) );
  XOR U3132 ( .A(n35329), .B(n35655), .Z(n35333) );
  XOR U3133 ( .A(n34561), .B(n34887), .Z(n34565) );
  XOR U3134 ( .A(n33769), .B(n34095), .Z(n33773) );
  XOR U3135 ( .A(n32953), .B(n33279), .Z(n32957) );
  XOR U3136 ( .A(n32113), .B(n32439), .Z(n32117) );
  XOR U3137 ( .A(n31249), .B(n31575), .Z(n31253) );
  XOR U3138 ( .A(n30361), .B(n30687), .Z(n30365) );
  XOR U3139 ( .A(n29449), .B(n29775), .Z(n29453) );
  XOR U3140 ( .A(n28513), .B(n28839), .Z(n28517) );
  XOR U3141 ( .A(n27553), .B(n27879), .Z(n27557) );
  XOR U3142 ( .A(n26567), .B(n26893), .Z(n26571) );
  XOR U3143 ( .A(n25558), .B(n25884), .Z(n25562) );
  XOR U3144 ( .A(n24521), .B(n24847), .Z(n24525) );
  XOR U3145 ( .A(n23465), .B(n23791), .Z(n23469) );
  XOR U3146 ( .A(n22383), .B(n22709), .Z(n22387) );
  XOR U3147 ( .A(n21279), .B(n21605), .Z(n21283) );
  XNOR U3148 ( .A(n21285), .B(n20720), .Z(n20722) );
  XNOR U3149 ( .A(n20156), .B(n19580), .Z(n19582) );
  XOR U3150 ( .A(n17642), .B(n18059), .Z(n17646) );
  XOR U3151 ( .A(n17597), .B(n18068), .Z(n17601) );
  XOR U3152 ( .A(n16375), .B(n16870), .Z(n16379) );
  XOR U3153 ( .A(n13814), .B(n14411), .Z(n13818) );
  XOR U3154 ( .A(n14432), .B(n15041), .Z(n14436) );
  XOR U3155 ( .A(n16355), .B(n16874), .Z(n16359) );
  XOR U3156 ( .A(n14477), .B(n15032), .Z(n14481) );
  XOR U3157 ( .A(n19542), .B(n19910), .Z(n19546) );
  XOR U3158 ( .A(n18229), .B(n18727), .Z(n18233) );
  XOR U3159 ( .A(n17019), .B(n17466), .Z(n17023) );
  XOR U3160 ( .A(n15785), .B(n16256), .Z(n15789) );
  XOR U3161 ( .A(n17672), .B(n18053), .Z(n17676) );
  XOR U3162 ( .A(n14507), .B(n15026), .Z(n14511) );
  XOR U3163 ( .A(n14462), .B(n15035), .Z(n14466) );
  XOR U3164 ( .A(n19572), .B(n19904), .Z(n19576) );
  XNOR U3165 ( .A(n39454), .B(n39142), .Z(n39144) );
  XNOR U3166 ( .A(n39145), .B(n38827), .Z(n38829) );
  XNOR U3167 ( .A(n38830), .B(n38506), .Z(n38508) );
  XNOR U3168 ( .A(n38509), .B(n38179), .Z(n38181) );
  XOR U3169 ( .A(n37504), .B(n37812), .Z(n37508) );
  XOR U3170 ( .A(n36808), .B(n37116), .Z(n36812) );
  XOR U3171 ( .A(n36088), .B(n36396), .Z(n36092) );
  XOR U3172 ( .A(n35344), .B(n35652), .Z(n35348) );
  XOR U3173 ( .A(n34576), .B(n34884), .Z(n34580) );
  XOR U3174 ( .A(n33784), .B(n34092), .Z(n33788) );
  XOR U3175 ( .A(n32968), .B(n33276), .Z(n32972) );
  XOR U3176 ( .A(n32128), .B(n32436), .Z(n32132) );
  XOR U3177 ( .A(n31264), .B(n31572), .Z(n31268) );
  XOR U3178 ( .A(n30376), .B(n30684), .Z(n30380) );
  XOR U3179 ( .A(n29464), .B(n29772), .Z(n29468) );
  XOR U3180 ( .A(n28528), .B(n28836), .Z(n28532) );
  XOR U3181 ( .A(n27568), .B(n27876), .Z(n27572) );
  XOR U3182 ( .A(n26582), .B(n26890), .Z(n26586) );
  XOR U3183 ( .A(n25573), .B(n25881), .Z(n25577) );
  XOR U3184 ( .A(n24536), .B(n24844), .Z(n24540) );
  XOR U3185 ( .A(n23480), .B(n23788), .Z(n23484) );
  XOR U3186 ( .A(n22398), .B(n22706), .Z(n22402) );
  XOR U3187 ( .A(n21294), .B(n21602), .Z(n21298) );
  XOR U3188 ( .A(n20165), .B(n20473), .Z(n20169) );
  XOR U3189 ( .A(n19008), .B(n19322), .Z(n19012) );
  XOR U3190 ( .A(n17702), .B(n18047), .Z(n17706) );
  XOR U3191 ( .A(n18259), .B(n18715), .Z(n18263) );
  XOR U3192 ( .A(n17049), .B(n17460), .Z(n17053) );
  XOR U3193 ( .A(n15815), .B(n16250), .Z(n15819) );
  XOR U3194 ( .A(n16390), .B(n16867), .Z(n16394) );
  XOR U3195 ( .A(n15144), .B(n15645), .Z(n15148) );
  XOR U3196 ( .A(n11877), .B(n12494), .Z(n11881) );
  XOR U3197 ( .A(n12515), .B(n13142), .Z(n12519) );
  XOR U3198 ( .A(n14492), .B(n15029), .Z(n14496) );
  XOR U3199 ( .A(n12560), .B(n13133), .Z(n12564) );
  XOR U3200 ( .A(n16420), .B(n16861), .Z(n16424) );
  XOR U3201 ( .A(n15174), .B(n15639), .Z(n15178) );
  XOR U3202 ( .A(n13904), .B(n14393), .Z(n13908) );
  XOR U3203 ( .A(n18289), .B(n18703), .Z(n18293) );
  XOR U3204 ( .A(n17079), .B(n17454), .Z(n17083) );
  XOR U3205 ( .A(n15845), .B(n16244), .Z(n15849) );
  XOR U3206 ( .A(n17732), .B(n18041), .Z(n17736) );
  XOR U3207 ( .A(n12590), .B(n13127), .Z(n12594) );
  XOR U3208 ( .A(n12545), .B(n13136), .Z(n12549) );
  XNOR U3209 ( .A(n40360), .B(n40066), .Z(n40068) );
  XNOR U3210 ( .A(n40069), .B(n39769), .Z(n39771) );
  XNOR U3211 ( .A(n39772), .B(n39466), .Z(n39468) );
  XNOR U3212 ( .A(n39469), .B(n39157), .Z(n39159) );
  XNOR U3213 ( .A(n39160), .B(n38842), .Z(n38844) );
  XOR U3214 ( .A(n38191), .B(n38481), .Z(n38195) );
  XOR U3215 ( .A(n37519), .B(n37809), .Z(n37523) );
  XOR U3216 ( .A(n36823), .B(n37113), .Z(n36827) );
  XOR U3217 ( .A(n36103), .B(n36393), .Z(n36107) );
  XOR U3218 ( .A(n35359), .B(n35649), .Z(n35363) );
  XOR U3219 ( .A(n34591), .B(n34881), .Z(n34595) );
  XOR U3220 ( .A(n33799), .B(n34089), .Z(n33803) );
  XOR U3221 ( .A(n32983), .B(n33273), .Z(n32987) );
  XOR U3222 ( .A(n32143), .B(n32433), .Z(n32147) );
  XOR U3223 ( .A(n31279), .B(n31569), .Z(n31283) );
  XOR U3224 ( .A(n30391), .B(n30681), .Z(n30395) );
  XOR U3225 ( .A(n29479), .B(n29769), .Z(n29483) );
  XOR U3226 ( .A(n28543), .B(n28833), .Z(n28547) );
  XOR U3227 ( .A(n27583), .B(n27873), .Z(n27587) );
  XOR U3228 ( .A(n26597), .B(n26887), .Z(n26601) );
  XOR U3229 ( .A(n25588), .B(n25878), .Z(n25592) );
  XOR U3230 ( .A(n24551), .B(n24841), .Z(n24555) );
  XOR U3231 ( .A(n23495), .B(n23785), .Z(n23499) );
  XOR U3232 ( .A(n22413), .B(n22703), .Z(n22417) );
  XOR U3233 ( .A(n21309), .B(n21599), .Z(n21313) );
  XOR U3234 ( .A(n20180), .B(n20470), .Z(n20184) );
  XOR U3235 ( .A(n19028), .B(n19318), .Z(n19032) );
  XOR U3236 ( .A(n18319), .B(n18691), .Z(n18323) );
  XOR U3237 ( .A(n17109), .B(n17448), .Z(n17113) );
  XOR U3238 ( .A(n15875), .B(n16238), .Z(n15879) );
  XOR U3239 ( .A(n16450), .B(n16855), .Z(n16454) );
  XOR U3240 ( .A(n15204), .B(n15633), .Z(n15208) );
  XOR U3241 ( .A(n13934), .B(n14387), .Z(n13938) );
  XOR U3242 ( .A(n14527), .B(n15022), .Z(n14531) );
  XOR U3243 ( .A(n9888), .B(n10521), .Z(n9892) );
  XOR U3244 ( .A(n10542), .B(n11187), .Z(n10546) );
  XOR U3245 ( .A(n13225), .B(n13768), .Z(n13229) );
  XOR U3246 ( .A(n11917), .B(n12486), .Z(n11921) );
  XOR U3247 ( .A(n9918), .B(n10515), .Z(n9922) );
  XOR U3248 ( .A(n14557), .B(n15016), .Z(n14561) );
  XOR U3249 ( .A(n13275), .B(n13758), .Z(n13279) );
  XOR U3250 ( .A(n16480), .B(n16849), .Z(n16484) );
  XOR U3251 ( .A(n15234), .B(n15627), .Z(n15238) );
  XOR U3252 ( .A(n13964), .B(n14381), .Z(n13968) );
  XOR U3253 ( .A(n17139), .B(n17442), .Z(n17143) );
  XOR U3254 ( .A(n15905), .B(n16232), .Z(n15909) );
  XOR U3255 ( .A(n11947), .B(n12480), .Z(n11951) );
  XOR U3256 ( .A(n10617), .B(n11172), .Z(n10621) );
  XOR U3257 ( .A(n10572), .B(n11181), .Z(n10576) );
  XNOR U3258 ( .A(n41212), .B(n40936), .Z(n40938) );
  XNOR U3259 ( .A(n40939), .B(n40657), .Z(n40659) );
  XNOR U3260 ( .A(n40660), .B(n40372), .Z(n40374) );
  XNOR U3261 ( .A(n40375), .B(n40081), .Z(n40083) );
  XOR U3262 ( .A(n39478), .B(n39750), .Z(n39482) );
  XOR U3263 ( .A(n38854), .B(n39126), .Z(n38858) );
  XOR U3264 ( .A(n38206), .B(n38478), .Z(n38210) );
  XOR U3265 ( .A(n37534), .B(n37806), .Z(n37538) );
  XOR U3266 ( .A(n36838), .B(n37110), .Z(n36842) );
  XOR U3267 ( .A(n36118), .B(n36390), .Z(n36122) );
  XOR U3268 ( .A(n35374), .B(n35646), .Z(n35378) );
  XOR U3269 ( .A(n34606), .B(n34878), .Z(n34610) );
  XOR U3270 ( .A(n33814), .B(n34086), .Z(n33818) );
  XOR U3271 ( .A(n32998), .B(n33270), .Z(n33002) );
  XOR U3272 ( .A(n32158), .B(n32430), .Z(n32162) );
  XOR U3273 ( .A(n31294), .B(n31566), .Z(n31298) );
  XOR U3274 ( .A(n30406), .B(n30678), .Z(n30410) );
  XOR U3275 ( .A(n29494), .B(n29766), .Z(n29498) );
  XOR U3276 ( .A(n28558), .B(n28830), .Z(n28562) );
  XOR U3277 ( .A(n27598), .B(n27870), .Z(n27602) );
  XOR U3278 ( .A(n26612), .B(n26884), .Z(n26616) );
  XOR U3279 ( .A(n25603), .B(n25875), .Z(n25607) );
  XOR U3280 ( .A(n24566), .B(n24838), .Z(n24570) );
  XOR U3281 ( .A(n23510), .B(n23782), .Z(n23514) );
  XOR U3282 ( .A(n22428), .B(n22700), .Z(n22432) );
  XOR U3283 ( .A(n21324), .B(n21596), .Z(n21328) );
  XOR U3284 ( .A(n20195), .B(n20467), .Z(n20199) );
  XOR U3285 ( .A(n19043), .B(n19315), .Z(n19047) );
  XOR U3286 ( .A(n15935), .B(n16226), .Z(n15939) );
  XOR U3287 ( .A(n16510), .B(n16843), .Z(n16514) );
  XOR U3288 ( .A(n15264), .B(n15621), .Z(n15268) );
  XOR U3289 ( .A(n13994), .B(n14375), .Z(n13998) );
  XOR U3290 ( .A(n14587), .B(n15010), .Z(n14591) );
  XOR U3291 ( .A(n13305), .B(n13752), .Z(n13309) );
  XOR U3292 ( .A(n12610), .B(n13123), .Z(n12614) );
  XOR U3293 ( .A(n7845), .B(n8496), .Z(n7849) );
  XOR U3294 ( .A(n8517), .B(n9180), .Z(n8521) );
  XOR U3295 ( .A(n11270), .B(n11831), .Z(n11274) );
  XOR U3296 ( .A(n11315), .B(n11822), .Z(n11319) );
  XOR U3297 ( .A(n17757), .B(n18036), .Z(n17761) );
  XOR U3298 ( .A(n9253), .B(n9844), .Z(n9257) );
  XOR U3299 ( .A(n7875), .B(n8490), .Z(n7879) );
  XOR U3300 ( .A(n12640), .B(n13117), .Z(n12644) );
  XOR U3301 ( .A(n14617), .B(n15004), .Z(n14621) );
  XOR U3302 ( .A(n13335), .B(n13746), .Z(n13339) );
  XOR U3303 ( .A(n16540), .B(n16837), .Z(n16544) );
  XOR U3304 ( .A(n15294), .B(n15615), .Z(n15298) );
  XOR U3305 ( .A(n14024), .B(n14369), .Z(n14028) );
  XOR U3306 ( .A(n11345), .B(n11816), .Z(n11349) );
  XOR U3307 ( .A(n9278), .B(n9839), .Z(n9282) );
  XOR U3308 ( .A(n8547), .B(n9174), .Z(n8551) );
  XNOR U3309 ( .A(n42010), .B(n41752), .Z(n41754) );
  XNOR U3310 ( .A(n41755), .B(n41491), .Z(n41493) );
  XNOR U3311 ( .A(n41494), .B(n41224), .Z(n41226) );
  XNOR U3312 ( .A(n41227), .B(n40951), .Z(n40953) );
  XNOR U3313 ( .A(n40954), .B(n40672), .Z(n40674) );
  XOR U3314 ( .A(n40093), .B(n40347), .Z(n40097) );
  XOR U3315 ( .A(n39493), .B(n39747), .Z(n39497) );
  XOR U3316 ( .A(n38869), .B(n39123), .Z(n38873) );
  XOR U3317 ( .A(n38221), .B(n38475), .Z(n38225) );
  XOR U3318 ( .A(n37549), .B(n37803), .Z(n37553) );
  XOR U3319 ( .A(n36853), .B(n37107), .Z(n36857) );
  XOR U3320 ( .A(n36133), .B(n36387), .Z(n36137) );
  XOR U3321 ( .A(n35389), .B(n35643), .Z(n35393) );
  XOR U3322 ( .A(n34621), .B(n34875), .Z(n34625) );
  XOR U3323 ( .A(n33829), .B(n34083), .Z(n33833) );
  XOR U3324 ( .A(n33013), .B(n33267), .Z(n33017) );
  XOR U3325 ( .A(n32173), .B(n32427), .Z(n32177) );
  XOR U3326 ( .A(n31309), .B(n31563), .Z(n31313) );
  XOR U3327 ( .A(n30421), .B(n30675), .Z(n30425) );
  XOR U3328 ( .A(n29509), .B(n29763), .Z(n29513) );
  XOR U3329 ( .A(n28573), .B(n28827), .Z(n28577) );
  XOR U3330 ( .A(n27613), .B(n27867), .Z(n27617) );
  XOR U3331 ( .A(n26627), .B(n26881), .Z(n26631) );
  XOR U3332 ( .A(n25618), .B(n25872), .Z(n25622) );
  XOR U3333 ( .A(n24581), .B(n24835), .Z(n24585) );
  XOR U3334 ( .A(n23525), .B(n23779), .Z(n23529) );
  XOR U3335 ( .A(n22443), .B(n22697), .Z(n22447) );
  XOR U3336 ( .A(n21339), .B(n21593), .Z(n21343) );
  XOR U3337 ( .A(n20210), .B(n20464), .Z(n20214) );
  XOR U3338 ( .A(n19058), .B(n19312), .Z(n19062) );
  XOR U3339 ( .A(n18369), .B(n18671), .Z(n18373) );
  XOR U3340 ( .A(n15965), .B(n16220), .Z(n15969) );
  XOR U3341 ( .A(n16570), .B(n16831), .Z(n16574) );
  XOR U3342 ( .A(n15324), .B(n15609), .Z(n15328) );
  XOR U3343 ( .A(n14054), .B(n14363), .Z(n14058) );
  XOR U3344 ( .A(n14647), .B(n14998), .Z(n14651) );
  XOR U3345 ( .A(n13365), .B(n13740), .Z(n13369) );
  XOR U3346 ( .A(n12670), .B(n13111), .Z(n12674) );
  XOR U3347 ( .A(n10637), .B(n11168), .Z(n10641) );
  XOR U3348 ( .A(n7905), .B(n8484), .Z(n7909) );
  XOR U3349 ( .A(n5748), .B(n6417), .Z(n5752) );
  XOR U3350 ( .A(n6438), .B(n7119), .Z(n6442) );
  XOR U3351 ( .A(n9308), .B(n9833), .Z(n9312) );
  XOR U3352 ( .A(n11375), .B(n11810), .Z(n11379) );
  XOR U3353 ( .A(n8582), .B(n9167), .Z(n8586) );
  XOR U3354 ( .A(n7192), .B(n7801), .Z(n7196) );
  XOR U3355 ( .A(n5778), .B(n6411), .Z(n5782) );
  XOR U3356 ( .A(n10667), .B(n11162), .Z(n10671) );
  XOR U3357 ( .A(n7935), .B(n8478), .Z(n7939) );
  XOR U3358 ( .A(n12700), .B(n13105), .Z(n12704) );
  XOR U3359 ( .A(n14677), .B(n14992), .Z(n14681) );
  XOR U3360 ( .A(n13395), .B(n13734), .Z(n13399) );
  XOR U3361 ( .A(n14084), .B(n14357), .Z(n14088) );
  XOR U3362 ( .A(n11405), .B(n11804), .Z(n11409) );
  XOR U3363 ( .A(n9338), .B(n9827), .Z(n9342) );
  XOR U3364 ( .A(n7172), .B(n7805), .Z(n7176) );
  XOR U3365 ( .A(n3570), .B(n4287), .Z(n3574) );
  XNOR U3366 ( .A(n42754), .B(n42514), .Z(n42516) );
  XNOR U3367 ( .A(n42517), .B(n42271), .Z(n42273) );
  XNOR U3368 ( .A(n42274), .B(n42022), .Z(n42024) );
  XNOR U3369 ( .A(n42025), .B(n41767), .Z(n41769) );
  XOR U3370 ( .A(n41236), .B(n41472), .Z(n41240) );
  XOR U3371 ( .A(n40684), .B(n40920), .Z(n40688) );
  XOR U3372 ( .A(n40108), .B(n40344), .Z(n40112) );
  XOR U3373 ( .A(n39508), .B(n39744), .Z(n39512) );
  XOR U3374 ( .A(n38884), .B(n39120), .Z(n38888) );
  XOR U3375 ( .A(n38236), .B(n38472), .Z(n38240) );
  XOR U3376 ( .A(n37564), .B(n37800), .Z(n37568) );
  XOR U3377 ( .A(n36868), .B(n37104), .Z(n36872) );
  XOR U3378 ( .A(n36148), .B(n36384), .Z(n36152) );
  XOR U3379 ( .A(n35404), .B(n35640), .Z(n35408) );
  XOR U3380 ( .A(n34636), .B(n34872), .Z(n34640) );
  XOR U3381 ( .A(n33844), .B(n34080), .Z(n33848) );
  XOR U3382 ( .A(n33028), .B(n33264), .Z(n33032) );
  XOR U3383 ( .A(n32188), .B(n32424), .Z(n32192) );
  XOR U3384 ( .A(n31324), .B(n31560), .Z(n31328) );
  XOR U3385 ( .A(n30436), .B(n30672), .Z(n30440) );
  XOR U3386 ( .A(n29524), .B(n29760), .Z(n29528) );
  XOR U3387 ( .A(n28588), .B(n28824), .Z(n28592) );
  XOR U3388 ( .A(n27628), .B(n27864), .Z(n27632) );
  XOR U3389 ( .A(n26642), .B(n26878), .Z(n26646) );
  XOR U3390 ( .A(n25633), .B(n25869), .Z(n25637) );
  XOR U3391 ( .A(n24596), .B(n24832), .Z(n24600) );
  XOR U3392 ( .A(n23540), .B(n23776), .Z(n23544) );
  XOR U3393 ( .A(n22458), .B(n22694), .Z(n22462) );
  XOR U3394 ( .A(n21354), .B(n21590), .Z(n21358) );
  XOR U3395 ( .A(n20225), .B(n20461), .Z(n20229) );
  XOR U3396 ( .A(n19073), .B(n19309), .Z(n19077) );
  XOR U3397 ( .A(n18384), .B(n18665), .Z(n18388) );
  XOR U3398 ( .A(n17194), .B(n17431), .Z(n17198) );
  XOR U3399 ( .A(n15980), .B(n16217), .Z(n15984) );
  XOR U3400 ( .A(n14707), .B(n14986), .Z(n14711) );
  XOR U3401 ( .A(n13425), .B(n13728), .Z(n13429) );
  XOR U3402 ( .A(n12730), .B(n13099), .Z(n12734) );
  XOR U3403 ( .A(n10697), .B(n11156), .Z(n10701) );
  XOR U3404 ( .A(n7965), .B(n8472), .Z(n7969) );
  XOR U3405 ( .A(n8612), .B(n9161), .Z(n8616) );
  XOR U3406 ( .A(n7222), .B(n7795), .Z(n7226) );
  XOR U3407 ( .A(n5808), .B(n6405), .Z(n5812) );
  XOR U3408 ( .A(n5763), .B(n6414), .Z(n5767) );
  XOR U3409 ( .A(n4323), .B(n4998), .Z(n4327) );
  XOR U3410 ( .A(n4303), .B(n5002), .Z(n4307) );
  XOR U3411 ( .A(n9368), .B(n9821), .Z(n9372) );
  XOR U3412 ( .A(n11435), .B(n11798), .Z(n11439) );
  XOR U3413 ( .A(n6503), .B(n7106), .Z(n6507) );
  XOR U3414 ( .A(n5075), .B(n5704), .Z(n5079) );
  XOR U3415 ( .A(n3625), .B(n4276), .Z(n3629) );
  XOR U3416 ( .A(n8642), .B(n9155), .Z(n8646) );
  XOR U3417 ( .A(n7252), .B(n7789), .Z(n7256) );
  XOR U3418 ( .A(n5838), .B(n6399), .Z(n5842) );
  XOR U3419 ( .A(n10727), .B(n11150), .Z(n10731) );
  XOR U3420 ( .A(n7995), .B(n8466), .Z(n7999) );
  XOR U3421 ( .A(n12760), .B(n13093), .Z(n12764) );
  XOR U3422 ( .A(n14737), .B(n14980), .Z(n14741) );
  XOR U3423 ( .A(n13455), .B(n13722), .Z(n13459) );
  XOR U3424 ( .A(n14752), .B(n14977), .Z(n14756) );
  XOR U3425 ( .A(n11465), .B(n11792), .Z(n11469) );
  XOR U3426 ( .A(n9398), .B(n9815), .Z(n9402) );
  XOR U3427 ( .A(n2131), .B(n2830), .Z(n2135) );
  XNOR U3428 ( .A(n43444), .B(n43222), .Z(n43224) );
  XNOR U3429 ( .A(n43225), .B(n42997), .Z(n42999) );
  XNOR U3430 ( .A(n43000), .B(n42766), .Z(n42768) );
  XNOR U3431 ( .A(n42769), .B(n42529), .Z(n42531) );
  XNOR U3432 ( .A(n42532), .B(n42286), .Z(n42288) );
  XOR U3433 ( .A(n41779), .B(n41997), .Z(n41783) );
  XOR U3434 ( .A(n41251), .B(n41469), .Z(n41255) );
  XOR U3435 ( .A(n40699), .B(n40917), .Z(n40703) );
  XOR U3436 ( .A(n40123), .B(n40341), .Z(n40127) );
  XOR U3437 ( .A(n39523), .B(n39741), .Z(n39527) );
  XOR U3438 ( .A(n38899), .B(n39117), .Z(n38903) );
  XOR U3439 ( .A(n38251), .B(n38469), .Z(n38255) );
  XOR U3440 ( .A(n37579), .B(n37797), .Z(n37583) );
  XOR U3441 ( .A(n36883), .B(n37101), .Z(n36887) );
  XOR U3442 ( .A(n36163), .B(n36381), .Z(n36167) );
  XOR U3443 ( .A(n35419), .B(n35637), .Z(n35423) );
  XOR U3444 ( .A(n34651), .B(n34869), .Z(n34655) );
  XOR U3445 ( .A(n33859), .B(n34077), .Z(n33863) );
  XOR U3446 ( .A(n33043), .B(n33261), .Z(n33047) );
  XOR U3447 ( .A(n32203), .B(n32421), .Z(n32207) );
  XOR U3448 ( .A(n31339), .B(n31557), .Z(n31343) );
  XOR U3449 ( .A(n30451), .B(n30669), .Z(n30455) );
  XOR U3450 ( .A(n29539), .B(n29757), .Z(n29543) );
  XOR U3451 ( .A(n28603), .B(n28821), .Z(n28607) );
  XOR U3452 ( .A(n27643), .B(n27861), .Z(n27647) );
  XOR U3453 ( .A(n26657), .B(n26875), .Z(n26661) );
  XOR U3454 ( .A(n25648), .B(n25866), .Z(n25652) );
  XOR U3455 ( .A(n24611), .B(n24829), .Z(n24615) );
  XOR U3456 ( .A(n23555), .B(n23773), .Z(n23559) );
  XOR U3457 ( .A(n22473), .B(n22691), .Z(n22477) );
  XOR U3458 ( .A(n21369), .B(n21587), .Z(n21373) );
  XOR U3459 ( .A(n20240), .B(n20458), .Z(n20244) );
  XOR U3460 ( .A(n19088), .B(n19306), .Z(n19092) );
  XOR U3461 ( .A(n18399), .B(n18659), .Z(n18403) );
  XOR U3462 ( .A(n17209), .B(n17428), .Z(n17213) );
  XOR U3463 ( .A(n15995), .B(n16214), .Z(n15999) );
  XOR U3464 ( .A(n13485), .B(n13716), .Z(n13489) );
  XOR U3465 ( .A(n12790), .B(n13087), .Z(n12794) );
  XOR U3466 ( .A(n10757), .B(n11144), .Z(n10761) );
  XOR U3467 ( .A(n8025), .B(n8460), .Z(n8029) );
  XOR U3468 ( .A(n8672), .B(n9149), .Z(n8676) );
  XOR U3469 ( .A(n7282), .B(n7783), .Z(n7286) );
  XOR U3470 ( .A(n5868), .B(n6393), .Z(n5872) );
  XOR U3471 ( .A(n6533), .B(n7100), .Z(n6537) );
  XOR U3472 ( .A(n5105), .B(n5698), .Z(n5109) );
  XOR U3473 ( .A(n3655), .B(n4270), .Z(n3659) );
  XOR U3474 ( .A(n4338), .B(n4995), .Z(n4342) );
  XOR U3475 ( .A(n2876), .B(n3557), .Z(n2880) );
  XOR U3476 ( .A(n2116), .B(n2833), .Z(n2120) );
  XOR U3477 ( .A(n9428), .B(n9809), .Z(n9432) );
  XOR U3478 ( .A(n11495), .B(n11786), .Z(n11499) );
  XOR U3479 ( .A(n4368), .B(n4989), .Z(n4372) );
  XOR U3480 ( .A(n2906), .B(n3551), .Z(n2910) );
  XOR U3481 ( .A(n1420), .B(n2089), .Z(n1424) );
  XOR U3482 ( .A(n6563), .B(n7094), .Z(n6567) );
  XOR U3483 ( .A(n5135), .B(n5692), .Z(n5139) );
  XOR U3484 ( .A(n3685), .B(n4264), .Z(n3689) );
  XOR U3485 ( .A(n8702), .B(n9143), .Z(n8706) );
  XOR U3486 ( .A(n7312), .B(n7777), .Z(n7316) );
  XOR U3487 ( .A(n5898), .B(n6387), .Z(n5902) );
  XOR U3488 ( .A(n10787), .B(n11138), .Z(n10791) );
  XOR U3489 ( .A(n8055), .B(n8454), .Z(n8059) );
  XOR U3490 ( .A(n12820), .B(n13081), .Z(n12824) );
  XOR U3491 ( .A(n11525), .B(n11780), .Z(n11529) );
  XOR U3492 ( .A(n9458), .B(n9803), .Z(n9462) );
  XNOR U3493 ( .A(n44080), .B(n43876), .Z(n43878) );
  XNOR U3494 ( .A(n43879), .B(n43669), .Z(n43671) );
  XNOR U3495 ( .A(n43672), .B(n43456), .Z(n43458) );
  XNOR U3496 ( .A(n43459), .B(n43237), .Z(n43239) );
  XOR U3497 ( .A(n42778), .B(n42978), .Z(n42782) );
  XOR U3498 ( .A(n42298), .B(n42498), .Z(n42302) );
  XOR U3499 ( .A(n41794), .B(n41994), .Z(n41798) );
  XOR U3500 ( .A(n41266), .B(n41466), .Z(n41270) );
  XOR U3501 ( .A(n40714), .B(n40914), .Z(n40718) );
  XOR U3502 ( .A(n40138), .B(n40338), .Z(n40142) );
  XOR U3503 ( .A(n39538), .B(n39738), .Z(n39542) );
  XOR U3504 ( .A(n38914), .B(n39114), .Z(n38918) );
  XOR U3505 ( .A(n38266), .B(n38466), .Z(n38270) );
  XOR U3506 ( .A(n37594), .B(n37794), .Z(n37598) );
  XOR U3507 ( .A(n36898), .B(n37098), .Z(n36902) );
  XOR U3508 ( .A(n36178), .B(n36378), .Z(n36182) );
  XOR U3509 ( .A(n35434), .B(n35634), .Z(n35438) );
  XOR U3510 ( .A(n34666), .B(n34866), .Z(n34670) );
  XOR U3511 ( .A(n33874), .B(n34074), .Z(n33878) );
  XOR U3512 ( .A(n33058), .B(n33258), .Z(n33062) );
  XOR U3513 ( .A(n32218), .B(n32418), .Z(n32222) );
  XOR U3514 ( .A(n31354), .B(n31554), .Z(n31358) );
  XOR U3515 ( .A(n30466), .B(n30666), .Z(n30470) );
  XOR U3516 ( .A(n29554), .B(n29754), .Z(n29558) );
  XOR U3517 ( .A(n28618), .B(n28818), .Z(n28622) );
  XOR U3518 ( .A(n27658), .B(n27858), .Z(n27662) );
  XOR U3519 ( .A(n26672), .B(n26872), .Z(n26676) );
  XOR U3520 ( .A(n25663), .B(n25863), .Z(n25667) );
  XOR U3521 ( .A(n24626), .B(n24826), .Z(n24630) );
  XOR U3522 ( .A(n23570), .B(n23770), .Z(n23574) );
  XOR U3523 ( .A(n22488), .B(n22688), .Z(n22492) );
  XOR U3524 ( .A(n21384), .B(n21584), .Z(n21388) );
  XOR U3525 ( .A(n20255), .B(n20455), .Z(n20259) );
  XOR U3526 ( .A(n19103), .B(n19303), .Z(n19107) );
  XOR U3527 ( .A(n17822), .B(n18023), .Z(n17826) );
  XOR U3528 ( .A(n16620), .B(n16821), .Z(n16624) );
  XOR U3529 ( .A(n15394), .B(n15595), .Z(n15398) );
  XOR U3530 ( .A(n14144), .B(n14345), .Z(n14148) );
  XOR U3531 ( .A(n12850), .B(n13075), .Z(n12854) );
  XOR U3532 ( .A(n10817), .B(n11132), .Z(n10821) );
  XOR U3533 ( .A(n8085), .B(n8448), .Z(n8089) );
  XOR U3534 ( .A(n8732), .B(n9137), .Z(n8736) );
  XOR U3535 ( .A(n7342), .B(n7771), .Z(n7346) );
  XOR U3536 ( .A(n5928), .B(n6381), .Z(n5932) );
  XOR U3537 ( .A(n6593), .B(n7088), .Z(n6597) );
  XOR U3538 ( .A(n5165), .B(n5686), .Z(n5169) );
  XOR U3539 ( .A(n3715), .B(n4258), .Z(n3719) );
  XOR U3540 ( .A(n4398), .B(n4983), .Z(n4402) );
  XOR U3541 ( .A(n2936), .B(n3545), .Z(n2940) );
  XOR U3542 ( .A(n1450), .B(n2083), .Z(n1454) );
  XOR U3543 ( .A(n2151), .B(n2826), .Z(n2155) );
  XOR U3544 ( .A(n9488), .B(n9797), .Z(n9492) );
  XOR U3545 ( .A(n11555), .B(n11774), .Z(n11559) );
  XOR U3546 ( .A(n2181), .B(n2820), .Z(n2185) );
  XOR U3547 ( .A(n4428), .B(n4977), .Z(n4432) );
  XOR U3548 ( .A(n2966), .B(n3539), .Z(n2970) );
  XOR U3549 ( .A(n1480), .B(n2077), .Z(n1484) );
  XOR U3550 ( .A(n6623), .B(n7082), .Z(n6627) );
  XOR U3551 ( .A(n5195), .B(n5680), .Z(n5199) );
  XOR U3552 ( .A(n3745), .B(n4252), .Z(n3749) );
  XOR U3553 ( .A(n8762), .B(n9131), .Z(n8766) );
  XOR U3554 ( .A(n7372), .B(n7765), .Z(n7376) );
  XOR U3555 ( .A(n5958), .B(n6375), .Z(n5962) );
  XOR U3556 ( .A(n10847), .B(n11126), .Z(n10851) );
  XOR U3557 ( .A(n8115), .B(n8442), .Z(n8119) );
  XOR U3558 ( .A(n12222), .B(n12425), .Z(n12226) );
  XOR U3559 ( .A(n9518), .B(n9791), .Z(n9522) );
  XNOR U3560 ( .A(n44662), .B(n44476), .Z(n44478) );
  XNOR U3561 ( .A(n44479), .B(n44287), .Z(n44289) );
  XNOR U3562 ( .A(n44290), .B(n44092), .Z(n44094) );
  XNOR U3563 ( .A(n44095), .B(n43891), .Z(n43893) );
  XNOR U3564 ( .A(n43894), .B(n43684), .Z(n43686) );
  XOR U3565 ( .A(n43249), .B(n43431), .Z(n43253) );
  XOR U3566 ( .A(n42793), .B(n42975), .Z(n42797) );
  XOR U3567 ( .A(n42313), .B(n42495), .Z(n42317) );
  XOR U3568 ( .A(n41809), .B(n41991), .Z(n41813) );
  XOR U3569 ( .A(n41281), .B(n41463), .Z(n41285) );
  XOR U3570 ( .A(n40729), .B(n40911), .Z(n40733) );
  XOR U3571 ( .A(n40153), .B(n40335), .Z(n40157) );
  XOR U3572 ( .A(n39553), .B(n39735), .Z(n39557) );
  XOR U3573 ( .A(n38929), .B(n39111), .Z(n38933) );
  XOR U3574 ( .A(n38281), .B(n38463), .Z(n38285) );
  XOR U3575 ( .A(n37609), .B(n37791), .Z(n37613) );
  XOR U3576 ( .A(n36913), .B(n37095), .Z(n36917) );
  XOR U3577 ( .A(n36193), .B(n36375), .Z(n36197) );
  XOR U3578 ( .A(n35449), .B(n35631), .Z(n35453) );
  XOR U3579 ( .A(n34681), .B(n34863), .Z(n34685) );
  XOR U3580 ( .A(n33889), .B(n34071), .Z(n33893) );
  XOR U3581 ( .A(n33073), .B(n33255), .Z(n33077) );
  XOR U3582 ( .A(n32233), .B(n32415), .Z(n32237) );
  XOR U3583 ( .A(n31369), .B(n31551), .Z(n31373) );
  XOR U3584 ( .A(n30481), .B(n30663), .Z(n30485) );
  XOR U3585 ( .A(n29569), .B(n29751), .Z(n29573) );
  XOR U3586 ( .A(n28633), .B(n28815), .Z(n28637) );
  XOR U3587 ( .A(n27673), .B(n27855), .Z(n27677) );
  XOR U3588 ( .A(n26687), .B(n26869), .Z(n26691) );
  XOR U3589 ( .A(n25678), .B(n25860), .Z(n25682) );
  XOR U3590 ( .A(n24641), .B(n24823), .Z(n24645) );
  XOR U3591 ( .A(n23585), .B(n23767), .Z(n23589) );
  XOR U3592 ( .A(n22503), .B(n22685), .Z(n22507) );
  XOR U3593 ( .A(n21399), .B(n21581), .Z(n21403) );
  XOR U3594 ( .A(n20270), .B(n20452), .Z(n20274) );
  XOR U3595 ( .A(n19118), .B(n19300), .Z(n19122) );
  XOR U3596 ( .A(n17837), .B(n18020), .Z(n17841) );
  XOR U3597 ( .A(n16635), .B(n16818), .Z(n16639) );
  XOR U3598 ( .A(n15409), .B(n15592), .Z(n15413) );
  XOR U3599 ( .A(n14159), .B(n14342), .Z(n14163) );
  XOR U3600 ( .A(n12885), .B(n13068), .Z(n12889) );
  XOR U3601 ( .A(n10877), .B(n11120), .Z(n10881) );
  XOR U3602 ( .A(n8145), .B(n8436), .Z(n8149) );
  XOR U3603 ( .A(n8792), .B(n9125), .Z(n8796) );
  XOR U3604 ( .A(n7402), .B(n7759), .Z(n7406) );
  XOR U3605 ( .A(n5988), .B(n6369), .Z(n5992) );
  XOR U3606 ( .A(n6653), .B(n7076), .Z(n6657) );
  XOR U3607 ( .A(n5225), .B(n5674), .Z(n5229) );
  XOR U3608 ( .A(n3775), .B(n4246), .Z(n3779) );
  XOR U3609 ( .A(n4458), .B(n4971), .Z(n4462) );
  XOR U3610 ( .A(n2996), .B(n3533), .Z(n3000) );
  XOR U3611 ( .A(n1510), .B(n2071), .Z(n1514) );
  XOR U3612 ( .A(n2211), .B(n2814), .Z(n2215) );
  XOR U3613 ( .A(n9548), .B(n9785), .Z(n9552) );
  XOR U3614 ( .A(n12242), .B(n12421), .Z(n12246) );
  XOR U3615 ( .A(n2241), .B(n2808), .Z(n2245) );
  XOR U3616 ( .A(n4488), .B(n4965), .Z(n4492) );
  XOR U3617 ( .A(n3026), .B(n3527), .Z(n3030) );
  XOR U3618 ( .A(n1540), .B(n2065), .Z(n1544) );
  XOR U3619 ( .A(n6683), .B(n7070), .Z(n6687) );
  XOR U3620 ( .A(n5255), .B(n5668), .Z(n5259) );
  XOR U3621 ( .A(n3805), .B(n4240), .Z(n3809) );
  XOR U3622 ( .A(n8822), .B(n9119), .Z(n8826) );
  XOR U3623 ( .A(n7432), .B(n7753), .Z(n7436) );
  XOR U3624 ( .A(n6018), .B(n6363), .Z(n6022) );
  XOR U3625 ( .A(n10907), .B(n11114), .Z(n10911) );
  XOR U3626 ( .A(n8175), .B(n8430), .Z(n8179) );
  XOR U3627 ( .A(n9578), .B(n9779), .Z(n9582) );
  XNOR U3628 ( .A(n45190), .B(n45022), .Z(n45024) );
  XNOR U3629 ( .A(n45025), .B(n44851), .Z(n44853) );
  XNOR U3630 ( .A(n44854), .B(n44674), .Z(n44676) );
  XNOR U3631 ( .A(n44677), .B(n44491), .Z(n44493) );
  XOR U3632 ( .A(n44104), .B(n44268), .Z(n44108) );
  XOR U3633 ( .A(n43696), .B(n43860), .Z(n43700) );
  XOR U3634 ( .A(n43264), .B(n43428), .Z(n43268) );
  XOR U3635 ( .A(n42808), .B(n42972), .Z(n42812) );
  XOR U3636 ( .A(n42328), .B(n42492), .Z(n42332) );
  XOR U3637 ( .A(n41824), .B(n41988), .Z(n41828) );
  XOR U3638 ( .A(n41296), .B(n41460), .Z(n41300) );
  XOR U3639 ( .A(n40744), .B(n40908), .Z(n40748) );
  XOR U3640 ( .A(n40168), .B(n40332), .Z(n40172) );
  XOR U3641 ( .A(n39568), .B(n39732), .Z(n39572) );
  XOR U3642 ( .A(n38944), .B(n39108), .Z(n38948) );
  XOR U3643 ( .A(n38296), .B(n38460), .Z(n38300) );
  XOR U3644 ( .A(n37624), .B(n37788), .Z(n37628) );
  XOR U3645 ( .A(n36928), .B(n37092), .Z(n36932) );
  XOR U3646 ( .A(n36208), .B(n36372), .Z(n36212) );
  XOR U3647 ( .A(n35464), .B(n35628), .Z(n35468) );
  XOR U3648 ( .A(n34696), .B(n34860), .Z(n34700) );
  XOR U3649 ( .A(n33904), .B(n34068), .Z(n33908) );
  XOR U3650 ( .A(n33088), .B(n33252), .Z(n33092) );
  XOR U3651 ( .A(n32248), .B(n32412), .Z(n32252) );
  XOR U3652 ( .A(n31384), .B(n31548), .Z(n31388) );
  XOR U3653 ( .A(n30496), .B(n30660), .Z(n30500) );
  XOR U3654 ( .A(n29584), .B(n29748), .Z(n29588) );
  XOR U3655 ( .A(n28648), .B(n28812), .Z(n28652) );
  XOR U3656 ( .A(n27688), .B(n27852), .Z(n27692) );
  XOR U3657 ( .A(n26702), .B(n26866), .Z(n26706) );
  XOR U3658 ( .A(n25693), .B(n25857), .Z(n25697) );
  XOR U3659 ( .A(n24656), .B(n24820), .Z(n24660) );
  XOR U3660 ( .A(n23600), .B(n23764), .Z(n23604) );
  XOR U3661 ( .A(n22518), .B(n22682), .Z(n22522) );
  XOR U3662 ( .A(n21414), .B(n21578), .Z(n21418) );
  XOR U3663 ( .A(n20285), .B(n20449), .Z(n20289) );
  XOR U3664 ( .A(n19133), .B(n19297), .Z(n19137) );
  XOR U3665 ( .A(n17852), .B(n18017), .Z(n17856) );
  XOR U3666 ( .A(n16650), .B(n16815), .Z(n16654) );
  XOR U3667 ( .A(n15424), .B(n15589), .Z(n15428) );
  XOR U3668 ( .A(n14174), .B(n14339), .Z(n14178) );
  XOR U3669 ( .A(n10937), .B(n11108), .Z(n10941) );
  XOR U3670 ( .A(n8205), .B(n8424), .Z(n8209) );
  XOR U3671 ( .A(n8852), .B(n9113), .Z(n8856) );
  XOR U3672 ( .A(n7462), .B(n7747), .Z(n7466) );
  XOR U3673 ( .A(n6048), .B(n6357), .Z(n6052) );
  XOR U3674 ( .A(n6713), .B(n7064), .Z(n6717) );
  XOR U3675 ( .A(n5285), .B(n5662), .Z(n5289) );
  XOR U3676 ( .A(n3835), .B(n4234), .Z(n3839) );
  XOR U3677 ( .A(n4518), .B(n4959), .Z(n4522) );
  XOR U3678 ( .A(n3056), .B(n3521), .Z(n3060) );
  XOR U3679 ( .A(n1570), .B(n2059), .Z(n1574) );
  XOR U3680 ( .A(n2271), .B(n2802), .Z(n2275) );
  XOR U3681 ( .A(n9608), .B(n9773), .Z(n9612) );
  XOR U3682 ( .A(n12905), .B(n13064), .Z(n12909) );
  XOR U3683 ( .A(n2301), .B(n2796), .Z(n2305) );
  XOR U3684 ( .A(n4548), .B(n4953), .Z(n4552) );
  XOR U3685 ( .A(n3086), .B(n3515), .Z(n3090) );
  XOR U3686 ( .A(n1600), .B(n2053), .Z(n1604) );
  XOR U3687 ( .A(n6743), .B(n7058), .Z(n6747) );
  XOR U3688 ( .A(n5315), .B(n5656), .Z(n5319) );
  XOR U3689 ( .A(n3865), .B(n4228), .Z(n3869) );
  XOR U3690 ( .A(n8882), .B(n9107), .Z(n8886) );
  XOR U3691 ( .A(n7492), .B(n7741), .Z(n7496) );
  XOR U3692 ( .A(n6078), .B(n6351), .Z(n6082) );
  XOR U3693 ( .A(n8235), .B(n8418), .Z(n8239) );
  XNOR U3694 ( .A(n45664), .B(n45514), .Z(n45516) );
  XNOR U3695 ( .A(n45517), .B(n45361), .Z(n45363) );
  XNOR U3696 ( .A(n45364), .B(n45202), .Z(n45204) );
  XNOR U3697 ( .A(n45205), .B(n45037), .Z(n45039) );
  XNOR U3698 ( .A(n45040), .B(n44866), .Z(n44868) );
  XOR U3699 ( .A(n44503), .B(n44649), .Z(n44507) );
  XOR U3700 ( .A(n44119), .B(n44265), .Z(n44123) );
  XOR U3701 ( .A(n43711), .B(n43857), .Z(n43715) );
  XOR U3702 ( .A(n43279), .B(n43425), .Z(n43283) );
  XOR U3703 ( .A(n42823), .B(n42969), .Z(n42827) );
  XOR U3704 ( .A(n42343), .B(n42489), .Z(n42347) );
  XOR U3705 ( .A(n41839), .B(n41985), .Z(n41843) );
  XOR U3706 ( .A(n41311), .B(n41457), .Z(n41315) );
  XOR U3707 ( .A(n40759), .B(n40905), .Z(n40763) );
  XOR U3708 ( .A(n40183), .B(n40329), .Z(n40187) );
  XOR U3709 ( .A(n39583), .B(n39729), .Z(n39587) );
  XOR U3710 ( .A(n38959), .B(n39105), .Z(n38963) );
  XOR U3711 ( .A(n38311), .B(n38457), .Z(n38315) );
  XOR U3712 ( .A(n37639), .B(n37785), .Z(n37643) );
  XOR U3713 ( .A(n36943), .B(n37089), .Z(n36947) );
  XOR U3714 ( .A(n36223), .B(n36369), .Z(n36227) );
  XOR U3715 ( .A(n35479), .B(n35625), .Z(n35483) );
  XOR U3716 ( .A(n34711), .B(n34857), .Z(n34715) );
  XOR U3717 ( .A(n33919), .B(n34065), .Z(n33923) );
  XOR U3718 ( .A(n33103), .B(n33249), .Z(n33107) );
  XOR U3719 ( .A(n32263), .B(n32409), .Z(n32267) );
  XOR U3720 ( .A(n31399), .B(n31545), .Z(n31403) );
  XOR U3721 ( .A(n30511), .B(n30657), .Z(n30515) );
  XOR U3722 ( .A(n29599), .B(n29745), .Z(n29603) );
  XOR U3723 ( .A(n28663), .B(n28809), .Z(n28667) );
  XOR U3724 ( .A(n27703), .B(n27849), .Z(n27707) );
  XOR U3725 ( .A(n26717), .B(n26863), .Z(n26721) );
  XOR U3726 ( .A(n25708), .B(n25854), .Z(n25712) );
  XOR U3727 ( .A(n24671), .B(n24817), .Z(n24675) );
  XOR U3728 ( .A(n23615), .B(n23761), .Z(n23619) );
  XOR U3729 ( .A(n22533), .B(n22679), .Z(n22537) );
  XOR U3730 ( .A(n21429), .B(n21575), .Z(n21433) );
  XOR U3731 ( .A(n20300), .B(n20446), .Z(n20304) );
  XOR U3732 ( .A(n19148), .B(n19294), .Z(n19152) );
  XOR U3733 ( .A(n17867), .B(n18014), .Z(n17871) );
  XOR U3734 ( .A(n16665), .B(n16812), .Z(n16669) );
  XOR U3735 ( .A(n15439), .B(n15586), .Z(n15443) );
  XOR U3736 ( .A(n11615), .B(n11762), .Z(n11619) );
  XOR U3737 ( .A(n8265), .B(n8412), .Z(n8269) );
  XOR U3738 ( .A(n8912), .B(n9101), .Z(n8916) );
  XOR U3739 ( .A(n7522), .B(n7735), .Z(n7526) );
  XOR U3740 ( .A(n6108), .B(n6345), .Z(n6112) );
  XOR U3741 ( .A(n6773), .B(n7052), .Z(n6777) );
  XOR U3742 ( .A(n5345), .B(n5650), .Z(n5349) );
  XOR U3743 ( .A(n3895), .B(n4222), .Z(n3899) );
  XOR U3744 ( .A(n4578), .B(n4947), .Z(n4582) );
  XOR U3745 ( .A(n3116), .B(n3509), .Z(n3120) );
  XOR U3746 ( .A(n1630), .B(n2047), .Z(n1634) );
  XOR U3747 ( .A(n2331), .B(n2790), .Z(n2335) );
  XOR U3748 ( .A(n14194), .B(n14335), .Z(n14198) );
  XOR U3749 ( .A(n12920), .B(n13061), .Z(n12924) );
  XOR U3750 ( .A(n10962), .B(n11103), .Z(n10966) );
  XOR U3751 ( .A(n2361), .B(n2784), .Z(n2365) );
  XOR U3752 ( .A(n4608), .B(n4941), .Z(n4612) );
  XOR U3753 ( .A(n3146), .B(n3503), .Z(n3150) );
  XOR U3754 ( .A(n1660), .B(n2041), .Z(n1664) );
  XOR U3755 ( .A(n6803), .B(n7046), .Z(n6807) );
  XOR U3756 ( .A(n5375), .B(n5644), .Z(n5379) );
  XOR U3757 ( .A(n3925), .B(n4216), .Z(n3929) );
  XOR U3758 ( .A(n8942), .B(n9095), .Z(n8946) );
  XOR U3759 ( .A(n7552), .B(n7729), .Z(n7556) );
  XOR U3760 ( .A(n6138), .B(n6339), .Z(n6142) );
  XNOR U3761 ( .A(n46084), .B(n45952), .Z(n45954) );
  XNOR U3762 ( .A(n45955), .B(n45817), .Z(n45819) );
  XNOR U3763 ( .A(n45820), .B(n45676), .Z(n45678) );
  XNOR U3764 ( .A(n45679), .B(n45529), .Z(n45531) );
  XOR U3765 ( .A(n45214), .B(n45342), .Z(n45218) );
  XOR U3766 ( .A(n44878), .B(n45006), .Z(n44882) );
  XOR U3767 ( .A(n44518), .B(n44646), .Z(n44522) );
  XOR U3768 ( .A(n44134), .B(n44262), .Z(n44138) );
  XOR U3769 ( .A(n43726), .B(n43854), .Z(n43730) );
  XOR U3770 ( .A(n43294), .B(n43422), .Z(n43298) );
  XOR U3771 ( .A(n42838), .B(n42966), .Z(n42842) );
  XOR U3772 ( .A(n42358), .B(n42486), .Z(n42362) );
  XOR U3773 ( .A(n41854), .B(n41982), .Z(n41858) );
  XOR U3774 ( .A(n41326), .B(n41454), .Z(n41330) );
  XOR U3775 ( .A(n40774), .B(n40902), .Z(n40778) );
  XOR U3776 ( .A(n40198), .B(n40326), .Z(n40202) );
  XOR U3777 ( .A(n39598), .B(n39726), .Z(n39602) );
  XOR U3778 ( .A(n38974), .B(n39102), .Z(n38978) );
  XOR U3779 ( .A(n38326), .B(n38454), .Z(n38330) );
  XOR U3780 ( .A(n37654), .B(n37782), .Z(n37658) );
  XOR U3781 ( .A(n36958), .B(n37086), .Z(n36962) );
  XOR U3782 ( .A(n36238), .B(n36366), .Z(n36242) );
  XOR U3783 ( .A(n35494), .B(n35622), .Z(n35498) );
  XOR U3784 ( .A(n34726), .B(n34854), .Z(n34730) );
  XOR U3785 ( .A(n33934), .B(n34062), .Z(n33938) );
  XOR U3786 ( .A(n33118), .B(n33246), .Z(n33122) );
  XOR U3787 ( .A(n32278), .B(n32406), .Z(n32282) );
  XOR U3788 ( .A(n31414), .B(n31542), .Z(n31418) );
  XOR U3789 ( .A(n30526), .B(n30654), .Z(n30530) );
  XOR U3790 ( .A(n29614), .B(n29742), .Z(n29618) );
  XOR U3791 ( .A(n28678), .B(n28806), .Z(n28682) );
  XOR U3792 ( .A(n27718), .B(n27846), .Z(n27722) );
  XOR U3793 ( .A(n26732), .B(n26860), .Z(n26736) );
  XOR U3794 ( .A(n25723), .B(n25851), .Z(n25727) );
  XOR U3795 ( .A(n24686), .B(n24814), .Z(n24690) );
  XOR U3796 ( .A(n23630), .B(n23758), .Z(n23634) );
  XOR U3797 ( .A(n22548), .B(n22676), .Z(n22552) );
  XOR U3798 ( .A(n21444), .B(n21572), .Z(n21448) );
  XOR U3799 ( .A(n20315), .B(n20443), .Z(n20319) );
  XOR U3800 ( .A(n19163), .B(n19291), .Z(n19167) );
  XOR U3801 ( .A(n17882), .B(n18011), .Z(n17886) );
  XOR U3802 ( .A(n16680), .B(n16809), .Z(n16684) );
  XOR U3803 ( .A(n7582), .B(n7723), .Z(n7586) );
  XOR U3804 ( .A(n6168), .B(n6333), .Z(n6172) );
  XOR U3805 ( .A(n6833), .B(n7040), .Z(n6837) );
  XOR U3806 ( .A(n5405), .B(n5638), .Z(n5409) );
  XOR U3807 ( .A(n3955), .B(n4210), .Z(n3959) );
  XOR U3808 ( .A(n4638), .B(n4935), .Z(n4642) );
  XOR U3809 ( .A(n3176), .B(n3497), .Z(n3180) );
  XOR U3810 ( .A(n1690), .B(n2035), .Z(n1694) );
  XOR U3811 ( .A(n2391), .B(n2778), .Z(n2395) );
  XOR U3812 ( .A(n15459), .B(n15582), .Z(n15463) );
  XOR U3813 ( .A(n14209), .B(n14332), .Z(n14213) );
  XOR U3814 ( .A(n12935), .B(n13058), .Z(n12939) );
  XOR U3815 ( .A(n11635), .B(n11758), .Z(n11639) );
  XOR U3816 ( .A(n9643), .B(n9766), .Z(n9647) );
  XOR U3817 ( .A(n2421), .B(n2772), .Z(n2425) );
  XOR U3818 ( .A(n4668), .B(n4929), .Z(n4672) );
  XOR U3819 ( .A(n3206), .B(n3491), .Z(n3210) );
  XOR U3820 ( .A(n1720), .B(n2029), .Z(n1724) );
  XOR U3821 ( .A(n6863), .B(n7034), .Z(n6867) );
  XOR U3822 ( .A(n5435), .B(n5632), .Z(n5439) );
  XOR U3823 ( .A(n3985), .B(n4204), .Z(n3989) );
  XOR U3824 ( .A(n6198), .B(n6327), .Z(n6202) );
  XOR U3825 ( .A(n10982), .B(n11099), .Z(n10986) );
  XOR U3826 ( .A(n8290), .B(n8407), .Z(n8294) );
  XNOR U3827 ( .A(n46450), .B(n46336), .Z(n46338) );
  XNOR U3828 ( .A(n46339), .B(n46219), .Z(n46221) );
  XNOR U3829 ( .A(n46222), .B(n46096), .Z(n46098) );
  XNOR U3830 ( .A(n46099), .B(n45967), .Z(n45969) );
  XNOR U3831 ( .A(n45970), .B(n45832), .Z(n45834) );
  XOR U3832 ( .A(n45541), .B(n45651), .Z(n45545) );
  XOR U3833 ( .A(n45229), .B(n45339), .Z(n45233) );
  XOR U3834 ( .A(n44893), .B(n45003), .Z(n44897) );
  XOR U3835 ( .A(n44533), .B(n44643), .Z(n44537) );
  XOR U3836 ( .A(n44149), .B(n44259), .Z(n44153) );
  XOR U3837 ( .A(n43741), .B(n43851), .Z(n43745) );
  XOR U3838 ( .A(n43309), .B(n43419), .Z(n43313) );
  XOR U3839 ( .A(n42853), .B(n42963), .Z(n42857) );
  XOR U3840 ( .A(n42373), .B(n42483), .Z(n42377) );
  XOR U3841 ( .A(n41869), .B(n41979), .Z(n41873) );
  XOR U3842 ( .A(n41341), .B(n41451), .Z(n41345) );
  XOR U3843 ( .A(n40789), .B(n40899), .Z(n40793) );
  XOR U3844 ( .A(n40213), .B(n40323), .Z(n40217) );
  XOR U3845 ( .A(n39613), .B(n39723), .Z(n39617) );
  XOR U3846 ( .A(n38989), .B(n39099), .Z(n38993) );
  XOR U3847 ( .A(n38341), .B(n38451), .Z(n38345) );
  XOR U3848 ( .A(n37669), .B(n37779), .Z(n37673) );
  XOR U3849 ( .A(n36973), .B(n37083), .Z(n36977) );
  XOR U3850 ( .A(n36253), .B(n36363), .Z(n36257) );
  XOR U3851 ( .A(n35509), .B(n35619), .Z(n35513) );
  XOR U3852 ( .A(n34741), .B(n34851), .Z(n34745) );
  XOR U3853 ( .A(n33949), .B(n34059), .Z(n33953) );
  XOR U3854 ( .A(n33133), .B(n33243), .Z(n33137) );
  XOR U3855 ( .A(n32293), .B(n32403), .Z(n32297) );
  XOR U3856 ( .A(n31429), .B(n31539), .Z(n31433) );
  XOR U3857 ( .A(n30541), .B(n30651), .Z(n30545) );
  XOR U3858 ( .A(n29629), .B(n29739), .Z(n29633) );
  XOR U3859 ( .A(n28693), .B(n28803), .Z(n28697) );
  XOR U3860 ( .A(n27733), .B(n27843), .Z(n27737) );
  XOR U3861 ( .A(n26747), .B(n26857), .Z(n26751) );
  XOR U3862 ( .A(n25738), .B(n25848), .Z(n25742) );
  XOR U3863 ( .A(n24701), .B(n24811), .Z(n24705) );
  XOR U3864 ( .A(n23645), .B(n23755), .Z(n23649) );
  XOR U3865 ( .A(n22563), .B(n22673), .Z(n22567) );
  XOR U3866 ( .A(n21459), .B(n21569), .Z(n21463) );
  XOR U3867 ( .A(n20330), .B(n20440), .Z(n20334) );
  XOR U3868 ( .A(n19178), .B(n19288), .Z(n19182) );
  XOR U3869 ( .A(n18489), .B(n18623), .Z(n18493) );
  XOR U3870 ( .A(n17299), .B(n17410), .Z(n17303) );
  XOR U3871 ( .A(n6893), .B(n7028), .Z(n6897) );
  XOR U3872 ( .A(n5465), .B(n5626), .Z(n5469) );
  XOR U3873 ( .A(n4015), .B(n4198), .Z(n4019) );
  XOR U3874 ( .A(n4698), .B(n4923), .Z(n4702) );
  XOR U3875 ( .A(n3236), .B(n3485), .Z(n3240) );
  XOR U3876 ( .A(n1750), .B(n2023), .Z(n1754) );
  XOR U3877 ( .A(n2451), .B(n2766), .Z(n2455) );
  XOR U3878 ( .A(n16090), .B(n16195), .Z(n16094) );
  XOR U3879 ( .A(n2481), .B(n2760), .Z(n2485) );
  XOR U3880 ( .A(n4728), .B(n4917), .Z(n4732) );
  XOR U3881 ( .A(n3266), .B(n3479), .Z(n3270) );
  XOR U3882 ( .A(n1780), .B(n2017), .Z(n1784) );
  XOR U3883 ( .A(n5495), .B(n5620), .Z(n5499) );
  XOR U3884 ( .A(n4045), .B(n4192), .Z(n4049) );
  XOR U3885 ( .A(n14857), .B(n14956), .Z(n14861) );
  XOR U3886 ( .A(n13595), .B(n13694), .Z(n13599) );
  XOR U3887 ( .A(n12307), .B(n12408), .Z(n12311) );
  XOR U3888 ( .A(n10997), .B(n11096), .Z(n11001) );
  XOR U3889 ( .A(n9663), .B(n9762), .Z(n9667) );
  XOR U3890 ( .A(n8305), .B(n8404), .Z(n8309) );
  XOR U3891 ( .A(n6923), .B(n7022), .Z(n6927) );
  XNOR U3892 ( .A(n46762), .B(n46666), .Z(n46668) );
  XNOR U3893 ( .A(n46669), .B(n46567), .Z(n46569) );
  XNOR U3894 ( .A(n46570), .B(n46462), .Z(n46464) );
  XNOR U3895 ( .A(n46465), .B(n46351), .Z(n46353) );
  XOR U3896 ( .A(n46108), .B(n46200), .Z(n46112) );
  XOR U3897 ( .A(n45844), .B(n45936), .Z(n45848) );
  XOR U3898 ( .A(n45556), .B(n45648), .Z(n45560) );
  XOR U3899 ( .A(n45244), .B(n45336), .Z(n45248) );
  XOR U3900 ( .A(n44908), .B(n45000), .Z(n44912) );
  XOR U3901 ( .A(n44548), .B(n44640), .Z(n44552) );
  XOR U3902 ( .A(n44164), .B(n44256), .Z(n44168) );
  XOR U3903 ( .A(n43756), .B(n43848), .Z(n43760) );
  XOR U3904 ( .A(n43324), .B(n43416), .Z(n43328) );
  XOR U3905 ( .A(n42868), .B(n42960), .Z(n42872) );
  XOR U3906 ( .A(n42388), .B(n42480), .Z(n42392) );
  XOR U3907 ( .A(n41884), .B(n41976), .Z(n41888) );
  XOR U3908 ( .A(n41356), .B(n41448), .Z(n41360) );
  XOR U3909 ( .A(n40804), .B(n40896), .Z(n40808) );
  XOR U3910 ( .A(n40228), .B(n40320), .Z(n40232) );
  XOR U3911 ( .A(n39628), .B(n39720), .Z(n39632) );
  XOR U3912 ( .A(n39004), .B(n39096), .Z(n39008) );
  XOR U3913 ( .A(n38356), .B(n38448), .Z(n38360) );
  XOR U3914 ( .A(n37684), .B(n37776), .Z(n37688) );
  XOR U3915 ( .A(n36988), .B(n37080), .Z(n36992) );
  XOR U3916 ( .A(n36268), .B(n36360), .Z(n36272) );
  XOR U3917 ( .A(n35524), .B(n35616), .Z(n35528) );
  XOR U3918 ( .A(n34756), .B(n34848), .Z(n34760) );
  XOR U3919 ( .A(n33964), .B(n34056), .Z(n33968) );
  XOR U3920 ( .A(n33148), .B(n33240), .Z(n33152) );
  XOR U3921 ( .A(n32308), .B(n32400), .Z(n32312) );
  XOR U3922 ( .A(n31444), .B(n31536), .Z(n31448) );
  XOR U3923 ( .A(n30556), .B(n30648), .Z(n30560) );
  XOR U3924 ( .A(n29644), .B(n29736), .Z(n29648) );
  XOR U3925 ( .A(n28708), .B(n28800), .Z(n28712) );
  XOR U3926 ( .A(n27748), .B(n27840), .Z(n27752) );
  XOR U3927 ( .A(n26762), .B(n26854), .Z(n26766) );
  XOR U3928 ( .A(n25753), .B(n25845), .Z(n25757) );
  XOR U3929 ( .A(n24716), .B(n24808), .Z(n24720) );
  XOR U3930 ( .A(n23660), .B(n23752), .Z(n23664) );
  XOR U3931 ( .A(n22578), .B(n22670), .Z(n22582) );
  XOR U3932 ( .A(n21474), .B(n21566), .Z(n21478) );
  XOR U3933 ( .A(n20345), .B(n20437), .Z(n20349) );
  XOR U3934 ( .A(n19193), .B(n19285), .Z(n19197) );
  XOR U3935 ( .A(n17912), .B(n18005), .Z(n17916) );
  XOR U3936 ( .A(n4075), .B(n4186), .Z(n4079) );
  XOR U3937 ( .A(n4758), .B(n4911), .Z(n4762) );
  XOR U3938 ( .A(n3296), .B(n3473), .Z(n3300) );
  XOR U3939 ( .A(n1810), .B(n2011), .Z(n1814) );
  XOR U3940 ( .A(n2511), .B(n2754), .Z(n2515) );
  XOR U3941 ( .A(n2541), .B(n2748), .Z(n2545) );
  XOR U3942 ( .A(n4788), .B(n4905), .Z(n4792) );
  XOR U3943 ( .A(n3326), .B(n3467), .Z(n3330) );
  XOR U3944 ( .A(n1840), .B(n2005), .Z(n1844) );
  XOR U3945 ( .A(n16720), .B(n16801), .Z(n16724) );
  XOR U3946 ( .A(n15494), .B(n15575), .Z(n15498) );
  XOR U3947 ( .A(n14244), .B(n14325), .Z(n14248) );
  XOR U3948 ( .A(n12970), .B(n13051), .Z(n12974) );
  XOR U3949 ( .A(n11670), .B(n11751), .Z(n11674) );
  XOR U3950 ( .A(n10348), .B(n10429), .Z(n10352) );
  XOR U3951 ( .A(n9002), .B(n9083), .Z(n9006) );
  XOR U3952 ( .A(n7632), .B(n7713), .Z(n7636) );
  XOR U3953 ( .A(n6238), .B(n6319), .Z(n6242) );
  XNOR U3954 ( .A(n47020), .B(n46942), .Z(n46944) );
  XNOR U3955 ( .A(n46945), .B(n46861), .Z(n46863) );
  XNOR U3956 ( .A(n46864), .B(n46774), .Z(n46776) );
  XNOR U3957 ( .A(n46777), .B(n46681), .Z(n46683) );
  XNOR U3958 ( .A(n46684), .B(n46582), .Z(n46584) );
  XOR U3959 ( .A(n46363), .B(n46437), .Z(n46367) );
  XOR U3960 ( .A(n46123), .B(n46197), .Z(n46127) );
  XOR U3961 ( .A(n45859), .B(n45933), .Z(n45863) );
  XOR U3962 ( .A(n45571), .B(n45645), .Z(n45575) );
  XOR U3963 ( .A(n45259), .B(n45333), .Z(n45263) );
  XOR U3964 ( .A(n44923), .B(n44997), .Z(n44927) );
  XOR U3965 ( .A(n44563), .B(n44637), .Z(n44567) );
  XOR U3966 ( .A(n44179), .B(n44253), .Z(n44183) );
  XOR U3967 ( .A(n43771), .B(n43845), .Z(n43775) );
  XOR U3968 ( .A(n43339), .B(n43413), .Z(n43343) );
  XOR U3969 ( .A(n42883), .B(n42957), .Z(n42887) );
  XOR U3970 ( .A(n42403), .B(n42477), .Z(n42407) );
  XOR U3971 ( .A(n41899), .B(n41973), .Z(n41903) );
  XOR U3972 ( .A(n41371), .B(n41445), .Z(n41375) );
  XOR U3973 ( .A(n40819), .B(n40893), .Z(n40823) );
  XOR U3974 ( .A(n40243), .B(n40317), .Z(n40247) );
  XOR U3975 ( .A(n39643), .B(n39717), .Z(n39647) );
  XOR U3976 ( .A(n39019), .B(n39093), .Z(n39023) );
  XOR U3977 ( .A(n38371), .B(n38445), .Z(n38375) );
  XOR U3978 ( .A(n37699), .B(n37773), .Z(n37703) );
  XOR U3979 ( .A(n37003), .B(n37077), .Z(n37007) );
  XOR U3980 ( .A(n36283), .B(n36357), .Z(n36287) );
  XOR U3981 ( .A(n35539), .B(n35613), .Z(n35543) );
  XOR U3982 ( .A(n34771), .B(n34845), .Z(n34775) );
  XOR U3983 ( .A(n33979), .B(n34053), .Z(n33983) );
  XOR U3984 ( .A(n33163), .B(n33237), .Z(n33167) );
  XOR U3985 ( .A(n32323), .B(n32397), .Z(n32327) );
  XOR U3986 ( .A(n31459), .B(n31533), .Z(n31463) );
  XOR U3987 ( .A(n30571), .B(n30645), .Z(n30575) );
  XOR U3988 ( .A(n29659), .B(n29733), .Z(n29663) );
  XOR U3989 ( .A(n28723), .B(n28797), .Z(n28727) );
  XOR U3990 ( .A(n27763), .B(n27837), .Z(n27767) );
  XOR U3991 ( .A(n26777), .B(n26851), .Z(n26781) );
  XOR U3992 ( .A(n25768), .B(n25842), .Z(n25772) );
  XOR U3993 ( .A(n24731), .B(n24805), .Z(n24735) );
  XOR U3994 ( .A(n23675), .B(n23749), .Z(n23679) );
  XOR U3995 ( .A(n22593), .B(n22667), .Z(n22597) );
  XOR U3996 ( .A(n21489), .B(n21563), .Z(n21493) );
  XOR U3997 ( .A(n20360), .B(n20434), .Z(n20364) );
  XOR U3998 ( .A(n19208), .B(n19282), .Z(n19212) );
  XOR U3999 ( .A(n18519), .B(n18611), .Z(n18523) );
  XOR U4000 ( .A(n4818), .B(n4899), .Z(n4822) );
  XOR U4001 ( .A(n3356), .B(n3461), .Z(n3360) );
  XOR U4002 ( .A(n1870), .B(n1999), .Z(n1874) );
  XOR U4003 ( .A(n2571), .B(n2742), .Z(n2575) );
  XOR U4004 ( .A(n2601), .B(n2736), .Z(n2605) );
  XOR U4005 ( .A(n1900), .B(n1993), .Z(n1904) );
  XOR U4006 ( .A(n17937), .B(n18000), .Z(n17941) );
  XOR U4007 ( .A(n16735), .B(n16798), .Z(n16739) );
  XOR U4008 ( .A(n14259), .B(n14322), .Z(n14263) );
  XOR U4009 ( .A(n12985), .B(n13048), .Z(n12989) );
  XOR U4010 ( .A(n11685), .B(n11748), .Z(n11689) );
  XOR U4011 ( .A(n10363), .B(n10426), .Z(n10367) );
  XOR U4012 ( .A(n9017), .B(n9080), .Z(n9021) );
  XOR U4013 ( .A(n7647), .B(n7710), .Z(n7651) );
  XOR U4014 ( .A(n6253), .B(n6316), .Z(n6257) );
  XOR U4015 ( .A(n4833), .B(n4896), .Z(n4837) );
  XOR U4016 ( .A(n2651), .B(n2726), .Z(n2655) );
  XNOR U4017 ( .A(n47223), .B(n47164), .Z(n47166) );
  XNOR U4018 ( .A(n47167), .B(n47101), .Z(n47103) );
  XNOR U4019 ( .A(n47104), .B(n47032), .Z(n47034) );
  XNOR U4020 ( .A(n47035), .B(n46957), .Z(n46959) );
  XOR U4021 ( .A(n46786), .B(n46842), .Z(n46790) );
  XOR U4022 ( .A(n46594), .B(n46650), .Z(n46598) );
  XOR U4023 ( .A(n46378), .B(n46434), .Z(n46382) );
  XOR U4024 ( .A(n46138), .B(n46194), .Z(n46142) );
  XOR U4025 ( .A(n45874), .B(n45930), .Z(n45878) );
  XOR U4026 ( .A(n45586), .B(n45642), .Z(n45590) );
  XOR U4027 ( .A(n45274), .B(n45330), .Z(n45278) );
  XOR U4028 ( .A(n44938), .B(n44994), .Z(n44942) );
  XOR U4029 ( .A(n44578), .B(n44634), .Z(n44582) );
  XOR U4030 ( .A(n44194), .B(n44250), .Z(n44198) );
  XOR U4031 ( .A(n43786), .B(n43842), .Z(n43790) );
  XOR U4032 ( .A(n43354), .B(n43410), .Z(n43358) );
  XOR U4033 ( .A(n42898), .B(n42954), .Z(n42902) );
  XOR U4034 ( .A(n42418), .B(n42474), .Z(n42422) );
  XOR U4035 ( .A(n41914), .B(n41970), .Z(n41918) );
  XOR U4036 ( .A(n41386), .B(n41442), .Z(n41390) );
  XOR U4037 ( .A(n40834), .B(n40890), .Z(n40838) );
  XOR U4038 ( .A(n40258), .B(n40314), .Z(n40262) );
  XOR U4039 ( .A(n39658), .B(n39714), .Z(n39662) );
  XOR U4040 ( .A(n39034), .B(n39090), .Z(n39038) );
  XOR U4041 ( .A(n38386), .B(n38442), .Z(n38390) );
  XOR U4042 ( .A(n37714), .B(n37770), .Z(n37718) );
  XOR U4043 ( .A(n37018), .B(n37074), .Z(n37022) );
  XOR U4044 ( .A(n36298), .B(n36354), .Z(n36302) );
  XOR U4045 ( .A(n35554), .B(n35610), .Z(n35558) );
  XOR U4046 ( .A(n34786), .B(n34842), .Z(n34790) );
  XOR U4047 ( .A(n33994), .B(n34050), .Z(n33998) );
  XOR U4048 ( .A(n33178), .B(n33234), .Z(n33182) );
  XOR U4049 ( .A(n32338), .B(n32394), .Z(n32342) );
  XOR U4050 ( .A(n31474), .B(n31530), .Z(n31478) );
  XOR U4051 ( .A(n30586), .B(n30642), .Z(n30590) );
  XOR U4052 ( .A(n29674), .B(n29730), .Z(n29678) );
  XOR U4053 ( .A(n28738), .B(n28794), .Z(n28742) );
  XOR U4054 ( .A(n27778), .B(n27834), .Z(n27782) );
  XOR U4055 ( .A(n26792), .B(n26848), .Z(n26796) );
  XOR U4056 ( .A(n25783), .B(n25839), .Z(n25787) );
  XOR U4057 ( .A(n24746), .B(n24802), .Z(n24750) );
  XOR U4058 ( .A(n23690), .B(n23746), .Z(n23694) );
  XOR U4059 ( .A(n22608), .B(n22664), .Z(n22612) );
  XOR U4060 ( .A(n21504), .B(n21560), .Z(n21508) );
  XOR U4061 ( .A(n20375), .B(n20431), .Z(n20379) );
  XOR U4062 ( .A(n19223), .B(n19279), .Z(n19227) );
  XOR U4063 ( .A(n16130), .B(n16187), .Z(n16134) );
  XOR U4064 ( .A(n2631), .B(n2730), .Z(n2635) );
  XOR U4065 ( .A(n17952), .B(n17997), .Z(n17956) );
  XOR U4066 ( .A(n15524), .B(n15569), .Z(n15528) );
  XOR U4067 ( .A(n14274), .B(n14319), .Z(n14278) );
  XOR U4068 ( .A(n13000), .B(n13045), .Z(n13004) );
  XOR U4069 ( .A(n11700), .B(n11745), .Z(n11704) );
  XOR U4070 ( .A(n10378), .B(n10423), .Z(n10382) );
  XOR U4071 ( .A(n9032), .B(n9077), .Z(n9036) );
  XOR U4072 ( .A(n7662), .B(n7707), .Z(n7666) );
  XOR U4073 ( .A(n6268), .B(n6313), .Z(n6272) );
  XOR U4074 ( .A(n4848), .B(n4893), .Z(n4852) );
  XOR U4075 ( .A(n3406), .B(n3451), .Z(n3410) );
  XOR U4076 ( .A(n1940), .B(n1985), .Z(n1944) );
  XOR U4077 ( .A(n47283), .B(n47321), .Z(n47287) );
  XNOR U4078 ( .A(n47289), .B(n47235), .Z(n47237) );
  XNOR U4079 ( .A(n47238), .B(n47179), .Z(n47181) );
  XOR U4080 ( .A(n46969), .B(n47007), .Z(n46973) );
  XOR U4081 ( .A(n46801), .B(n46839), .Z(n46805) );
  XOR U4082 ( .A(n46609), .B(n46647), .Z(n46613) );
  XOR U4083 ( .A(n46393), .B(n46431), .Z(n46397) );
  XOR U4084 ( .A(n46153), .B(n46191), .Z(n46157) );
  XOR U4085 ( .A(n45889), .B(n45927), .Z(n45893) );
  XOR U4086 ( .A(n45601), .B(n45639), .Z(n45605) );
  XOR U4087 ( .A(n45289), .B(n45327), .Z(n45293) );
  XOR U4088 ( .A(n44953), .B(n44991), .Z(n44957) );
  XOR U4089 ( .A(n44593), .B(n44631), .Z(n44597) );
  XOR U4090 ( .A(n44209), .B(n44247), .Z(n44213) );
  XOR U4091 ( .A(n43801), .B(n43839), .Z(n43805) );
  XOR U4092 ( .A(n43369), .B(n43407), .Z(n43373) );
  XOR U4093 ( .A(n42913), .B(n42951), .Z(n42917) );
  XOR U4094 ( .A(n42433), .B(n42471), .Z(n42437) );
  XOR U4095 ( .A(n41929), .B(n41967), .Z(n41933) );
  XOR U4096 ( .A(n41401), .B(n41439), .Z(n41405) );
  XOR U4097 ( .A(n40849), .B(n40887), .Z(n40853) );
  XOR U4098 ( .A(n40273), .B(n40311), .Z(n40277) );
  XOR U4099 ( .A(n39673), .B(n39711), .Z(n39677) );
  XOR U4100 ( .A(n39049), .B(n39087), .Z(n39053) );
  XOR U4101 ( .A(n38401), .B(n38439), .Z(n38405) );
  XOR U4102 ( .A(n37729), .B(n37767), .Z(n37733) );
  XOR U4103 ( .A(n37033), .B(n37071), .Z(n37037) );
  XOR U4104 ( .A(n36313), .B(n36351), .Z(n36317) );
  XOR U4105 ( .A(n35569), .B(n35607), .Z(n35573) );
  XOR U4106 ( .A(n34801), .B(n34839), .Z(n34805) );
  XOR U4107 ( .A(n34009), .B(n34047), .Z(n34013) );
  XOR U4108 ( .A(n33193), .B(n33231), .Z(n33197) );
  XOR U4109 ( .A(n32353), .B(n32391), .Z(n32357) );
  XOR U4110 ( .A(n31489), .B(n31527), .Z(n31493) );
  XOR U4111 ( .A(n30601), .B(n30639), .Z(n30605) );
  XOR U4112 ( .A(n29689), .B(n29727), .Z(n29693) );
  XOR U4113 ( .A(n28753), .B(n28791), .Z(n28757) );
  XOR U4114 ( .A(n27793), .B(n27831), .Z(n27797) );
  XOR U4115 ( .A(n26807), .B(n26845), .Z(n26811) );
  XOR U4116 ( .A(n25798), .B(n25836), .Z(n25802) );
  XOR U4117 ( .A(n24761), .B(n24799), .Z(n24765) );
  XOR U4118 ( .A(n23705), .B(n23743), .Z(n23709) );
  XOR U4119 ( .A(n22623), .B(n22661), .Z(n22627) );
  XOR U4120 ( .A(n21519), .B(n21557), .Z(n21523) );
  XOR U4121 ( .A(n20390), .B(n20428), .Z(n20394) );
  XOR U4122 ( .A(n19238), .B(n19276), .Z(n19242) );
  XOR U4123 ( .A(n17359), .B(n17398), .Z(n17363) );
  XOR U4124 ( .A(n47118), .B(n47150), .Z(n47122) );
  XOR U4125 ( .A(n16765), .B(n16792), .Z(n16769) );
  XOR U4126 ( .A(n15539), .B(n15566), .Z(n15543) );
  XOR U4127 ( .A(n14289), .B(n14316), .Z(n14293) );
  XOR U4128 ( .A(n13015), .B(n13042), .Z(n13019) );
  XOR U4129 ( .A(n11715), .B(n11742), .Z(n11719) );
  XOR U4130 ( .A(n10393), .B(n10420), .Z(n10397) );
  XOR U4131 ( .A(n9047), .B(n9074), .Z(n9051) );
  XOR U4132 ( .A(n7677), .B(n7704), .Z(n7681) );
  XOR U4133 ( .A(n6283), .B(n6310), .Z(n6287) );
  XOR U4134 ( .A(n4863), .B(n4890), .Z(n4867) );
  XOR U4135 ( .A(n3421), .B(n3448), .Z(n3425) );
  XOR U4136 ( .A(n1955), .B(n1982), .Z(n1959) );
  XOR U4137 ( .A(n47415), .B(n47435), .Z(n47419) );
  XOR U4138 ( .A(n47343), .B(n47363), .Z(n47347) );
  XNOR U4139 ( .A(n47349), .B(n47301), .Z(n47303) );
  XNOR U4140 ( .A(n47253), .B(n47194), .Z(n47196) );
  XOR U4141 ( .A(n47059), .B(n47079), .Z(n47063) );
  XOR U4142 ( .A(n46903), .B(n46923), .Z(n46907) );
  XOR U4143 ( .A(n46723), .B(n46743), .Z(n46727) );
  XOR U4144 ( .A(n46519), .B(n46539), .Z(n46523) );
  XOR U4145 ( .A(n46291), .B(n46311), .Z(n46295) );
  XOR U4146 ( .A(n46039), .B(n46059), .Z(n46043) );
  XOR U4147 ( .A(n45763), .B(n45783), .Z(n45767) );
  XOR U4148 ( .A(n45463), .B(n45483), .Z(n45467) );
  XOR U4149 ( .A(n45139), .B(n45159), .Z(n45143) );
  XOR U4150 ( .A(n44791), .B(n44811), .Z(n44795) );
  XOR U4151 ( .A(n44419), .B(n44439), .Z(n44423) );
  XOR U4152 ( .A(n44023), .B(n44043), .Z(n44027) );
  XOR U4153 ( .A(n43603), .B(n43623), .Z(n43607) );
  XOR U4154 ( .A(n43159), .B(n43179), .Z(n43163) );
  XOR U4155 ( .A(n42691), .B(n42711), .Z(n42695) );
  XOR U4156 ( .A(n42199), .B(n42219), .Z(n42203) );
  XOR U4157 ( .A(n41683), .B(n41703), .Z(n41687) );
  XOR U4158 ( .A(n41143), .B(n41163), .Z(n41147) );
  XOR U4159 ( .A(n40579), .B(n40599), .Z(n40583) );
  XOR U4160 ( .A(n39991), .B(n40011), .Z(n39995) );
  XOR U4161 ( .A(n39379), .B(n39399), .Z(n39383) );
  XOR U4162 ( .A(n38743), .B(n38763), .Z(n38747) );
  XOR U4163 ( .A(n38083), .B(n38103), .Z(n38087) );
  XOR U4164 ( .A(n37399), .B(n37419), .Z(n37403) );
  XOR U4165 ( .A(n36691), .B(n36711), .Z(n36695) );
  XOR U4166 ( .A(n35959), .B(n35979), .Z(n35963) );
  XOR U4167 ( .A(n35203), .B(n35223), .Z(n35207) );
  XOR U4168 ( .A(n34423), .B(n34443), .Z(n34427) );
  XOR U4169 ( .A(n33619), .B(n33639), .Z(n33623) );
  XOR U4170 ( .A(n32791), .B(n32811), .Z(n32795) );
  XOR U4171 ( .A(n31939), .B(n31959), .Z(n31943) );
  XOR U4172 ( .A(n31063), .B(n31083), .Z(n31067) );
  XOR U4173 ( .A(n30163), .B(n30183), .Z(n30167) );
  XOR U4174 ( .A(n29239), .B(n29259), .Z(n29243) );
  XOR U4175 ( .A(n28291), .B(n28311), .Z(n28295) );
  XOR U4176 ( .A(n27319), .B(n27339), .Z(n27323) );
  XOR U4177 ( .A(n26321), .B(n26341), .Z(n26325) );
  XOR U4178 ( .A(n25299), .B(n25319), .Z(n25303) );
  XOR U4179 ( .A(n24251), .B(n24271), .Z(n24255) );
  XOR U4180 ( .A(n23182), .B(n23202), .Z(n23186) );
  XOR U4181 ( .A(n22089), .B(n22109), .Z(n22093) );
  XOR U4182 ( .A(n20972), .B(n20992), .Z(n20976) );
  XOR U4183 ( .A(n19832), .B(n19852), .Z(n19836) );
  XNOR U4184 ( .A(n19838), .B(n19256), .Z(n19258) );
  XOR U4185 ( .A(n18564), .B(n18593), .Z(n18568) );
  XNOR U4186 ( .A(n47307), .B(n47306), .Z(n47264) );
  XNOR U4187 ( .A(n28394), .B(n27914), .Z(n27916) );
  XOR U4188 ( .A(n26934), .B(n27416), .Z(n26938) );
  XNOR U4189 ( .A(n26428), .B(n25924), .Z(n25926) );
  XOR U4190 ( .A(n29339), .B(n29797), .Z(n29343) );
  XOR U4191 ( .A(n28403), .B(n28861), .Z(n28407) );
  XNOR U4192 ( .A(n28409), .B(n27929), .Z(n27931) );
  XNOR U4193 ( .A(n27454), .B(n26962), .Z(n26964) );
  XOR U4194 ( .A(n26949), .B(n27413), .Z(n26953) );
  XNOR U4195 ( .A(n28419), .B(n27939), .Z(n27941) );
  XOR U4196 ( .A(n25936), .B(n26418), .Z(n25940) );
  XOR U4197 ( .A(n24893), .B(n25401), .Z(n24897) );
  XOR U4198 ( .A(n30713), .B(n31153), .Z(n30717) );
  XOR U4199 ( .A(n29813), .B(n30253), .Z(n29817) );
  XOR U4200 ( .A(n28889), .B(n29329), .Z(n28893) );
  XOR U4201 ( .A(n25443), .B(n25908), .Z(n25447) );
  XNOR U4202 ( .A(n28900), .B(n28426), .Z(n28428) );
  XNOR U4203 ( .A(n28429), .B(n27949), .Z(n27951) );
  XNOR U4204 ( .A(n27952), .B(n27466), .Z(n27468) );
  XNOR U4205 ( .A(n27469), .B(n26977), .Z(n26979) );
  XNOR U4206 ( .A(n26483), .B(n25979), .Z(n25981) );
  XOR U4207 ( .A(n24391), .B(n24876), .Z(n24395) );
  XOR U4208 ( .A(n23295), .B(n23825), .Z(n23299) );
  XNOR U4209 ( .A(n29829), .B(n29367), .Z(n29369) );
  XOR U4210 ( .A(n25971), .B(n26411), .Z(n25975) );
  XNOR U4211 ( .A(n25449), .B(n24931), .Z(n24933) );
  XOR U4212 ( .A(n24908), .B(n25398), .Z(n24912) );
  XOR U4213 ( .A(n23841), .B(n24353), .Z(n23845) );
  XNOR U4214 ( .A(n24949), .B(n24424), .Z(n24426) );
  XOR U4215 ( .A(n32033), .B(n32455), .Z(n32037) );
  XOR U4216 ( .A(n31169), .B(n31591), .Z(n31173) );
  XOR U4217 ( .A(n30281), .B(n30703), .Z(n30285) );
  XOR U4218 ( .A(n22757), .B(n23288), .Z(n22761) );
  XNOR U4219 ( .A(n23887), .B(n23353), .Z(n23355) );
  XNOR U4220 ( .A(n30292), .B(n29836), .Z(n29838) );
  XNOR U4221 ( .A(n29839), .B(n29377), .Z(n29379) );
  XNOR U4222 ( .A(n29380), .B(n28912), .Z(n28914) );
  XNOR U4223 ( .A(n28915), .B(n28441), .Z(n28443) );
  XNOR U4224 ( .A(n28444), .B(n27964), .Z(n27966) );
  XNOR U4225 ( .A(n27967), .B(n27481), .Z(n27483) );
  XNOR U4226 ( .A(n27484), .B(n26992), .Z(n26994) );
  XNOR U4227 ( .A(n26995), .B(n26495), .Z(n26497) );
  XNOR U4228 ( .A(n26498), .B(n25994), .Z(n25996) );
  XOR U4229 ( .A(n23330), .B(n23818), .Z(n23334) );
  XOR U4230 ( .A(n21649), .B(n22197), .Z(n21653) );
  XNOR U4231 ( .A(n31185), .B(n30741), .Z(n30743) );
  XNOR U4232 ( .A(n23917), .B(n23383), .Z(n23385) );
  XOR U4233 ( .A(n24411), .B(n24872), .Z(n24415) );
  XNOR U4234 ( .A(n23872), .B(n23338), .Z(n23340) );
  XOR U4235 ( .A(n22233), .B(n22740), .Z(n22237) );
  XOR U4236 ( .A(n23315), .B(n23821), .Z(n23319) );
  XNOR U4237 ( .A(n25489), .B(n24971), .Z(n24973) );
  XNOR U4238 ( .A(n24964), .B(n24439), .Z(n24441) );
  XNOR U4239 ( .A(n23897), .B(n23363), .Z(n23365) );
  XNOR U4240 ( .A(n23356), .B(n22815), .Z(n22817) );
  XOR U4241 ( .A(n33299), .B(n33703), .Z(n33303) );
  XOR U4242 ( .A(n32471), .B(n32875), .Z(n32475) );
  XOR U4243 ( .A(n31619), .B(n32023), .Z(n31623) );
  XOR U4244 ( .A(n22218), .B(n22743), .Z(n22222) );
  XOR U4245 ( .A(n21094), .B(n21642), .Z(n21098) );
  XNOR U4246 ( .A(n23902), .B(n23368), .Z(n23370) );
  XNOR U4247 ( .A(n22259), .B(n21707), .Z(n21709) );
  XNOR U4248 ( .A(n31630), .B(n31192), .Z(n31194) );
  XNOR U4249 ( .A(n31195), .B(n30751), .Z(n30753) );
  XNOR U4250 ( .A(n30754), .B(n30304), .Z(n30306) );
  XNOR U4251 ( .A(n30307), .B(n29851), .Z(n29853) );
  XNOR U4252 ( .A(n29854), .B(n29392), .Z(n29394) );
  XNOR U4253 ( .A(n29395), .B(n28927), .Z(n28929) );
  XNOR U4254 ( .A(n28930), .B(n28456), .Z(n28458) );
  XNOR U4255 ( .A(n28459), .B(n27979), .Z(n27981) );
  XNOR U4256 ( .A(n27982), .B(n27496), .Z(n27498) );
  XNOR U4257 ( .A(n27499), .B(n27007), .Z(n27009) );
  XNOR U4258 ( .A(n27010), .B(n26510), .Z(n26512) );
  XNOR U4259 ( .A(n26513), .B(n26009), .Z(n26011) );
  XNOR U4260 ( .A(n26012), .B(n25501), .Z(n25503) );
  XNOR U4261 ( .A(n25504), .B(n24986), .Z(n24988) );
  XNOR U4262 ( .A(n23386), .B(n22845), .Z(n22847) );
  XOR U4263 ( .A(n19950), .B(n20516), .Z(n19954) );
  XNOR U4264 ( .A(n23411), .B(n22870), .Z(n22872) );
  XNOR U4265 ( .A(n32487), .B(n32061), .Z(n32063) );
  XNOR U4266 ( .A(n23932), .B(n23398), .Z(n23400) );
  XNOR U4267 ( .A(n23391), .B(n22850), .Z(n22852) );
  XNOR U4268 ( .A(n22289), .B(n21737), .Z(n21739) );
  XOR U4269 ( .A(n22802), .B(n23279), .Z(n22806) );
  XNOR U4270 ( .A(n22244), .B(n21692), .Z(n21694) );
  XOR U4271 ( .A(n21124), .B(n21636), .Z(n21128) );
  XNOR U4272 ( .A(n23912), .B(n23378), .Z(n23380) );
  XNOR U4273 ( .A(n23371), .B(n22830), .Z(n22832) );
  XNOR U4274 ( .A(n22269), .B(n21717), .Z(n21719) );
  XNOR U4275 ( .A(n21710), .B(n21152), .Z(n21154) );
  XOR U4276 ( .A(n34511), .B(n34897), .Z(n34515) );
  XOR U4277 ( .A(n33719), .B(n34105), .Z(n33723) );
  XOR U4278 ( .A(n32903), .B(n33289), .Z(n32907) );
  XOR U4279 ( .A(n19980), .B(n20510), .Z(n19984) );
  XOR U4280 ( .A(n21109), .B(n21639), .Z(n21113) );
  XNOR U4281 ( .A(n22274), .B(n21722), .Z(n21724) );
  XNOR U4282 ( .A(n20578), .B(n20008), .Z(n20010) );
  XNOR U4283 ( .A(n32914), .B(n32494), .Z(n32496) );
  XNOR U4284 ( .A(n32497), .B(n32071), .Z(n32073) );
  XNOR U4285 ( .A(n32074), .B(n31642), .Z(n31644) );
  XNOR U4286 ( .A(n31645), .B(n31207), .Z(n31209) );
  XNOR U4287 ( .A(n31210), .B(n30766), .Z(n30768) );
  XNOR U4288 ( .A(n30769), .B(n30319), .Z(n30321) );
  XNOR U4289 ( .A(n30322), .B(n29866), .Z(n29868) );
  XNOR U4290 ( .A(n29869), .B(n29407), .Z(n29409) );
  XNOR U4291 ( .A(n29410), .B(n28942), .Z(n28944) );
  XNOR U4292 ( .A(n28945), .B(n28471), .Z(n28473) );
  XNOR U4293 ( .A(n28474), .B(n27994), .Z(n27996) );
  XNOR U4294 ( .A(n27997), .B(n27511), .Z(n27513) );
  XNOR U4295 ( .A(n27514), .B(n27022), .Z(n27024) );
  XNOR U4296 ( .A(n27025), .B(n26525), .Z(n26527) );
  XNOR U4297 ( .A(n26528), .B(n26024), .Z(n26026) );
  XNOR U4298 ( .A(n26027), .B(n25516), .Z(n25518) );
  XNOR U4299 ( .A(n25519), .B(n25002), .Z(n25004) );
  XNOR U4300 ( .A(n25005), .B(n24479), .Z(n24481) );
  XNOR U4301 ( .A(n24482), .B(n23954), .Z(n23956) );
  XNOR U4302 ( .A(n23957), .B(n23423), .Z(n23425) );
  XNOR U4303 ( .A(n21740), .B(n21182), .Z(n21184) );
  XOR U4304 ( .A(n19965), .B(n20513), .Z(n19969) );
  XNOR U4305 ( .A(n33735), .B(n33327), .Z(n33329) );
  XOR U4306 ( .A(n22862), .B(n23267), .Z(n22866) );
  XNOR U4307 ( .A(n22304), .B(n21752), .Z(n21754) );
  XNOR U4308 ( .A(n21745), .B(n21187), .Z(n21189) );
  XNOR U4309 ( .A(n20608), .B(n20038), .Z(n20040) );
  XOR U4310 ( .A(n21139), .B(n21633), .Z(n21143) );
  XNOR U4311 ( .A(n20563), .B(n19993), .Z(n19995) );
  XOR U4312 ( .A(n19407), .B(n19937), .Z(n19411) );
  XOR U4313 ( .A(n18094), .B(n18781), .Z(n18098) );
  XOR U4314 ( .A(n18798), .B(n19364), .Z(n18802) );
  XNOR U4315 ( .A(n22284), .B(n21732), .Z(n21734) );
  XNOR U4316 ( .A(n21725), .B(n21167), .Z(n21169) );
  XNOR U4317 ( .A(n20588), .B(n20018), .Z(n20020) );
  XNOR U4318 ( .A(n22329), .B(n21777), .Z(n21779) );
  XNOR U4319 ( .A(n21770), .B(n21212), .Z(n21214) );
  XOR U4320 ( .A(n35669), .B(n36037), .Z(n35673) );
  XOR U4321 ( .A(n34913), .B(n35281), .Z(n34917) );
  XOR U4322 ( .A(n34133), .B(n34501), .Z(n34137) );
  XNOR U4323 ( .A(n19971), .B(n19395), .Z(n19397) );
  XNOR U4324 ( .A(n20593), .B(n20023), .Z(n20025) );
  XOR U4325 ( .A(n18848), .B(n19354), .Z(n18852) );
  XOR U4326 ( .A(n22338), .B(n22719), .Z(n22342) );
  XNOR U4327 ( .A(n20638), .B(n20068), .Z(n20070) );
  XNOR U4328 ( .A(n34144), .B(n33742), .Z(n33744) );
  XNOR U4329 ( .A(n33745), .B(n33337), .Z(n33339) );
  XNOR U4330 ( .A(n33340), .B(n32926), .Z(n32928) );
  XNOR U4331 ( .A(n32929), .B(n32509), .Z(n32511) );
  XNOR U4332 ( .A(n32512), .B(n32086), .Z(n32088) );
  XNOR U4333 ( .A(n32089), .B(n31657), .Z(n31659) );
  XNOR U4334 ( .A(n31660), .B(n31222), .Z(n31224) );
  XNOR U4335 ( .A(n31225), .B(n30781), .Z(n30783) );
  XNOR U4336 ( .A(n30784), .B(n30334), .Z(n30336) );
  XNOR U4337 ( .A(n30337), .B(n29881), .Z(n29883) );
  XNOR U4338 ( .A(n29884), .B(n29422), .Z(n29424) );
  XNOR U4339 ( .A(n29425), .B(n28957), .Z(n28959) );
  XNOR U4340 ( .A(n28960), .B(n28486), .Z(n28488) );
  XNOR U4341 ( .A(n28489), .B(n28009), .Z(n28011) );
  XNOR U4342 ( .A(n28012), .B(n27526), .Z(n27528) );
  XNOR U4343 ( .A(n27529), .B(n27037), .Z(n27039) );
  XNOR U4344 ( .A(n27040), .B(n26540), .Z(n26542) );
  XNOR U4345 ( .A(n26543), .B(n26039), .Z(n26041) );
  XNOR U4346 ( .A(n26042), .B(n25531), .Z(n25533) );
  XNOR U4347 ( .A(n25534), .B(n25017), .Z(n25019) );
  XNOR U4348 ( .A(n25020), .B(n24494), .Z(n24496) );
  XNOR U4349 ( .A(n24497), .B(n23969), .Z(n23971) );
  XNOR U4350 ( .A(n23972), .B(n23438), .Z(n23440) );
  XNOR U4351 ( .A(n23441), .B(n22900), .Z(n22902) );
  XNOR U4352 ( .A(n22359), .B(n21807), .Z(n21809) );
  XNOR U4353 ( .A(n21800), .B(n21242), .Z(n21244) );
  XNOR U4354 ( .A(n34929), .B(n34539), .Z(n34541) );
  XNOR U4355 ( .A(n20668), .B(n20098), .Z(n20100) );
  XOR U4356 ( .A(n21199), .B(n21621), .Z(n21203) );
  XNOR U4357 ( .A(n20623), .B(n20053), .Z(n20055) );
  XNOR U4358 ( .A(n20046), .B(n19470), .Z(n19472) );
  XOR U4359 ( .A(n18878), .B(n19348), .Z(n18882) );
  XNOR U4360 ( .A(n20001), .B(n19425), .Z(n19427) );
  XOR U4361 ( .A(n18833), .B(n19357), .Z(n18837) );
  XOR U4362 ( .A(n17527), .B(n18082), .Z(n17531) );
  XOR U4363 ( .A(n18109), .B(n18775), .Z(n18113) );
  XOR U4364 ( .A(n16899), .B(n17490), .Z(n16903) );
  XNOR U4365 ( .A(n20603), .B(n20033), .Z(n20035) );
  XNOR U4366 ( .A(n20648), .B(n20078), .Z(n20080) );
  XNOR U4367 ( .A(n20071), .B(n19495), .Z(n19497) );
  XOR U4368 ( .A(n36773), .B(n37123), .Z(n36777) );
  XOR U4369 ( .A(n36053), .B(n36403), .Z(n36057) );
  XOR U4370 ( .A(n35309), .B(n35659), .Z(n35313) );
  XOR U4371 ( .A(n15670), .B(n16279), .Z(n15674) );
  XOR U4372 ( .A(n18863), .B(n19351), .Z(n18867) );
  XOR U4373 ( .A(n18159), .B(n18755), .Z(n18163) );
  XOR U4374 ( .A(n21229), .B(n21615), .Z(n21233) );
  XNOR U4375 ( .A(n35320), .B(n34936), .Z(n34938) );
  XNOR U4376 ( .A(n34939), .B(n34549), .Z(n34551) );
  XNOR U4377 ( .A(n34552), .B(n34156), .Z(n34158) );
  XNOR U4378 ( .A(n34159), .B(n33757), .Z(n33759) );
  XNOR U4379 ( .A(n33760), .B(n33352), .Z(n33354) );
  XNOR U4380 ( .A(n33355), .B(n32941), .Z(n32943) );
  XNOR U4381 ( .A(n32944), .B(n32524), .Z(n32526) );
  XNOR U4382 ( .A(n32527), .B(n32101), .Z(n32103) );
  XNOR U4383 ( .A(n32104), .B(n31672), .Z(n31674) );
  XNOR U4384 ( .A(n31675), .B(n31237), .Z(n31239) );
  XNOR U4385 ( .A(n31240), .B(n30796), .Z(n30798) );
  XNOR U4386 ( .A(n30799), .B(n30349), .Z(n30351) );
  XNOR U4387 ( .A(n30352), .B(n29896), .Z(n29898) );
  XNOR U4388 ( .A(n29899), .B(n29437), .Z(n29439) );
  XNOR U4389 ( .A(n29440), .B(n28972), .Z(n28974) );
  XNOR U4390 ( .A(n28975), .B(n28501), .Z(n28503) );
  XNOR U4391 ( .A(n28504), .B(n28024), .Z(n28026) );
  XNOR U4392 ( .A(n28027), .B(n27541), .Z(n27543) );
  XNOR U4393 ( .A(n27544), .B(n27052), .Z(n27054) );
  XNOR U4394 ( .A(n27055), .B(n26555), .Z(n26557) );
  XNOR U4395 ( .A(n26558), .B(n26054), .Z(n26056) );
  XNOR U4396 ( .A(n26057), .B(n25546), .Z(n25548) );
  XNOR U4397 ( .A(n25549), .B(n25032), .Z(n25034) );
  XNOR U4398 ( .A(n25035), .B(n24509), .Z(n24511) );
  XNOR U4399 ( .A(n24512), .B(n23984), .Z(n23986) );
  XNOR U4400 ( .A(n23987), .B(n23453), .Z(n23455) );
  XNOR U4401 ( .A(n23456), .B(n22915), .Z(n22917) );
  XNOR U4402 ( .A(n22918), .B(n22371), .Z(n22373) );
  XNOR U4403 ( .A(n21825), .B(n21267), .Z(n21269) );
  XNOR U4404 ( .A(n20678), .B(n20108), .Z(n20110) );
  XNOR U4405 ( .A(n20101), .B(n19525), .Z(n19527) );
  XNOR U4406 ( .A(n20056), .B(n19480), .Z(n19482) );
  XOR U4407 ( .A(n16954), .B(n17479), .Z(n16958) );
  XOR U4408 ( .A(n18209), .B(n18735), .Z(n18213) );
  XNOR U4409 ( .A(n36069), .B(n35697), .Z(n35699) );
  XOR U4410 ( .A(n21259), .B(n21609), .Z(n21263) );
  XNOR U4411 ( .A(n20061), .B(n19485), .Z(n19487) );
  XOR U4412 ( .A(n17542), .B(n18079), .Z(n17546) );
  XOR U4413 ( .A(n16320), .B(n16881), .Z(n16324) );
  XOR U4414 ( .A(n16914), .B(n17487), .Z(n16918) );
  XNOR U4415 ( .A(n20086), .B(n19510), .Z(n19512) );
  XOR U4416 ( .A(n18918), .B(n19340), .Z(n18922) );
  XNOR U4417 ( .A(n20708), .B(n20138), .Z(n20140) );
  XNOR U4418 ( .A(n20131), .B(n19555), .Z(n19557) );
  XOR U4419 ( .A(n37823), .B(n38155), .Z(n37827) );
  XOR U4420 ( .A(n37139), .B(n37471), .Z(n37143) );
  XOR U4421 ( .A(n36431), .B(n36763), .Z(n36435) );
  XOR U4422 ( .A(n18239), .B(n18723), .Z(n18243) );
  XOR U4423 ( .A(n18194), .B(n18741), .Z(n18198) );
  XOR U4424 ( .A(n16984), .B(n17473), .Z(n16988) );
  XOR U4425 ( .A(n15079), .B(n15658), .Z(n15083) );
  XOR U4426 ( .A(n15685), .B(n16276), .Z(n15689) );
  XOR U4427 ( .A(n14427), .B(n15042), .Z(n14431) );
  XOR U4428 ( .A(n18174), .B(n18749), .Z(n18178) );
  XNOR U4429 ( .A(n20091), .B(n19515), .Z(n19517) );
  XNOR U4430 ( .A(n36442), .B(n36076), .Z(n36078) );
  XNOR U4431 ( .A(n36079), .B(n35707), .Z(n35709) );
  XNOR U4432 ( .A(n35710), .B(n35332), .Z(n35334) );
  XNOR U4433 ( .A(n35335), .B(n34951), .Z(n34953) );
  XNOR U4434 ( .A(n34954), .B(n34564), .Z(n34566) );
  XNOR U4435 ( .A(n34567), .B(n34171), .Z(n34173) );
  XNOR U4436 ( .A(n34174), .B(n33772), .Z(n33774) );
  XNOR U4437 ( .A(n33775), .B(n33367), .Z(n33369) );
  XNOR U4438 ( .A(n33370), .B(n32956), .Z(n32958) );
  XNOR U4439 ( .A(n32959), .B(n32539), .Z(n32541) );
  XNOR U4440 ( .A(n32542), .B(n32116), .Z(n32118) );
  XNOR U4441 ( .A(n32119), .B(n31687), .Z(n31689) );
  XNOR U4442 ( .A(n31690), .B(n31252), .Z(n31254) );
  XNOR U4443 ( .A(n31255), .B(n30811), .Z(n30813) );
  XNOR U4444 ( .A(n30814), .B(n30364), .Z(n30366) );
  XNOR U4445 ( .A(n30367), .B(n29911), .Z(n29913) );
  XNOR U4446 ( .A(n29914), .B(n29452), .Z(n29454) );
  XNOR U4447 ( .A(n29455), .B(n28987), .Z(n28989) );
  XNOR U4448 ( .A(n28990), .B(n28516), .Z(n28518) );
  XNOR U4449 ( .A(n28519), .B(n28039), .Z(n28041) );
  XNOR U4450 ( .A(n28042), .B(n27556), .Z(n27558) );
  XNOR U4451 ( .A(n27559), .B(n27067), .Z(n27069) );
  XNOR U4452 ( .A(n27070), .B(n26570), .Z(n26572) );
  XNOR U4453 ( .A(n26573), .B(n26069), .Z(n26071) );
  XNOR U4454 ( .A(n26072), .B(n25561), .Z(n25563) );
  XNOR U4455 ( .A(n25564), .B(n25047), .Z(n25049) );
  XNOR U4456 ( .A(n25050), .B(n24524), .Z(n24526) );
  XNOR U4457 ( .A(n24527), .B(n23999), .Z(n24001) );
  XNOR U4458 ( .A(n24002), .B(n23468), .Z(n23470) );
  XNOR U4459 ( .A(n23471), .B(n22930), .Z(n22932) );
  XNOR U4460 ( .A(n22933), .B(n22386), .Z(n22388) );
  XNOR U4461 ( .A(n22389), .B(n21837), .Z(n21839) );
  XNOR U4462 ( .A(n21840), .B(n21282), .Z(n21284) );
  XNOR U4463 ( .A(n20116), .B(n19540), .Z(n19542) );
  XOR U4464 ( .A(n18948), .B(n19334), .Z(n18952) );
  XOR U4465 ( .A(n13150), .B(n13783), .Z(n13154) );
  XOR U4466 ( .A(n16969), .B(n17476), .Z(n16973) );
  XOR U4467 ( .A(n15735), .B(n16266), .Z(n15739) );
  XOR U4468 ( .A(n17622), .B(n18063), .Z(n17626) );
  XOR U4469 ( .A(n16400), .B(n16865), .Z(n16404) );
  XOR U4470 ( .A(n18269), .B(n18711), .Z(n18273) );
  XNOR U4471 ( .A(n37155), .B(n36801), .Z(n36803) );
  XNOR U4472 ( .A(n20121), .B(n19545), .Z(n19547) );
  XOR U4473 ( .A(n16335), .B(n16878), .Z(n16339) );
  XOR U4474 ( .A(n14482), .B(n15031), .Z(n14486) );
  XNOR U4475 ( .A(n20146), .B(n19570), .Z(n19572) );
  XOR U4476 ( .A(n18978), .B(n19328), .Z(n18982) );
  XOR U4477 ( .A(n38819), .B(n39133), .Z(n38823) );
  XOR U4478 ( .A(n38171), .B(n38485), .Z(n38175) );
  XOR U4479 ( .A(n37499), .B(n37813), .Z(n37503) );
  XOR U4480 ( .A(n18299), .B(n18699), .Z(n18303) );
  XOR U4481 ( .A(n17652), .B(n18057), .Z(n17656) );
  XOR U4482 ( .A(n16430), .B(n16859), .Z(n16434) );
  XOR U4483 ( .A(n16999), .B(n17470), .Z(n17003) );
  XOR U4484 ( .A(n15765), .B(n16260), .Z(n15769) );
  XOR U4485 ( .A(n15094), .B(n15655), .Z(n15098) );
  XOR U4486 ( .A(n13824), .B(n14409), .Z(n13828) );
  XOR U4487 ( .A(n14442), .B(n15039), .Z(n14446) );
  XNOR U4488 ( .A(n20151), .B(n19575), .Z(n19577) );
  XNOR U4489 ( .A(n37510), .B(n37162), .Z(n37164) );
  XNOR U4490 ( .A(n37165), .B(n36811), .Z(n36813) );
  XNOR U4491 ( .A(n36814), .B(n36454), .Z(n36456) );
  XNOR U4492 ( .A(n36457), .B(n36091), .Z(n36093) );
  XNOR U4493 ( .A(n36094), .B(n35722), .Z(n35724) );
  XNOR U4494 ( .A(n35725), .B(n35347), .Z(n35349) );
  XNOR U4495 ( .A(n35350), .B(n34966), .Z(n34968) );
  XNOR U4496 ( .A(n34969), .B(n34579), .Z(n34581) );
  XNOR U4497 ( .A(n34582), .B(n34186), .Z(n34188) );
  XNOR U4498 ( .A(n34189), .B(n33787), .Z(n33789) );
  XNOR U4499 ( .A(n33790), .B(n33382), .Z(n33384) );
  XNOR U4500 ( .A(n33385), .B(n32971), .Z(n32973) );
  XNOR U4501 ( .A(n32974), .B(n32554), .Z(n32556) );
  XNOR U4502 ( .A(n32557), .B(n32131), .Z(n32133) );
  XNOR U4503 ( .A(n32134), .B(n31702), .Z(n31704) );
  XNOR U4504 ( .A(n31705), .B(n31267), .Z(n31269) );
  XNOR U4505 ( .A(n31270), .B(n30826), .Z(n30828) );
  XNOR U4506 ( .A(n30829), .B(n30379), .Z(n30381) );
  XNOR U4507 ( .A(n30382), .B(n29926), .Z(n29928) );
  XNOR U4508 ( .A(n29929), .B(n29467), .Z(n29469) );
  XNOR U4509 ( .A(n29470), .B(n29002), .Z(n29004) );
  XNOR U4510 ( .A(n29005), .B(n28531), .Z(n28533) );
  XNOR U4511 ( .A(n28534), .B(n28054), .Z(n28056) );
  XNOR U4512 ( .A(n28057), .B(n27571), .Z(n27573) );
  XNOR U4513 ( .A(n27574), .B(n27082), .Z(n27084) );
  XNOR U4514 ( .A(n27085), .B(n26585), .Z(n26587) );
  XNOR U4515 ( .A(n26588), .B(n26084), .Z(n26086) );
  XNOR U4516 ( .A(n26087), .B(n25576), .Z(n25578) );
  XNOR U4517 ( .A(n25579), .B(n25062), .Z(n25064) );
  XNOR U4518 ( .A(n25065), .B(n24539), .Z(n24541) );
  XNOR U4519 ( .A(n24542), .B(n24014), .Z(n24016) );
  XNOR U4520 ( .A(n24017), .B(n23483), .Z(n23485) );
  XNOR U4521 ( .A(n23486), .B(n22945), .Z(n22947) );
  XNOR U4522 ( .A(n22948), .B(n22401), .Z(n22403) );
  XNOR U4523 ( .A(n22404), .B(n21852), .Z(n21854) );
  XNOR U4524 ( .A(n21855), .B(n21297), .Z(n21299) );
  XNOR U4525 ( .A(n21300), .B(n20735), .Z(n20737) );
  XNOR U4526 ( .A(n20738), .B(n20168), .Z(n20170) );
  XOR U4527 ( .A(n12535), .B(n13138), .Z(n12539) );
  XOR U4528 ( .A(n13165), .B(n13780), .Z(n13169) );
  XOR U4529 ( .A(n11857), .B(n12498), .Z(n11861) );
  XOR U4530 ( .A(n15750), .B(n16263), .Z(n15754) );
  XOR U4531 ( .A(n17029), .B(n17464), .Z(n17033) );
  XOR U4532 ( .A(n15795), .B(n16254), .Z(n15799) );
  XOR U4533 ( .A(n14537), .B(n15020), .Z(n14541) );
  XOR U4534 ( .A(n17682), .B(n18051), .Z(n17686) );
  XOR U4535 ( .A(n16460), .B(n16853), .Z(n16464) );
  XNOR U4536 ( .A(n38187), .B(n37851), .Z(n37853) );
  XOR U4537 ( .A(n19013), .B(n19321), .Z(n19017) );
  XOR U4538 ( .A(n10532), .B(n11189), .Z(n10536) );
  XOR U4539 ( .A(n14497), .B(n15028), .Z(n14501) );
  XOR U4540 ( .A(n13215), .B(n13770), .Z(n13219) );
  XOR U4541 ( .A(n39761), .B(n40057), .Z(n39765) );
  XOR U4542 ( .A(n39149), .B(n39445), .Z(n39153) );
  XOR U4543 ( .A(n38513), .B(n38809), .Z(n38517) );
  XOR U4544 ( .A(n17712), .B(n18045), .Z(n17716) );
  XOR U4545 ( .A(n16490), .B(n16847), .Z(n16494) );
  XOR U4546 ( .A(n17059), .B(n17458), .Z(n17063) );
  XOR U4547 ( .A(n15825), .B(n16248), .Z(n15829) );
  XOR U4548 ( .A(n14567), .B(n15014), .Z(n14571) );
  XOR U4549 ( .A(n15154), .B(n15643), .Z(n15158) );
  XOR U4550 ( .A(n13884), .B(n14397), .Z(n13888) );
  XOR U4551 ( .A(n13839), .B(n14406), .Z(n13843) );
  XNOR U4552 ( .A(n38524), .B(n38194), .Z(n38196) );
  XNOR U4553 ( .A(n38197), .B(n37861), .Z(n37863) );
  XNOR U4554 ( .A(n37864), .B(n37522), .Z(n37524) );
  XNOR U4555 ( .A(n37525), .B(n37177), .Z(n37179) );
  XNOR U4556 ( .A(n37180), .B(n36826), .Z(n36828) );
  XNOR U4557 ( .A(n36829), .B(n36469), .Z(n36471) );
  XNOR U4558 ( .A(n36472), .B(n36106), .Z(n36108) );
  XNOR U4559 ( .A(n36109), .B(n35737), .Z(n35739) );
  XNOR U4560 ( .A(n35740), .B(n35362), .Z(n35364) );
  XNOR U4561 ( .A(n35365), .B(n34981), .Z(n34983) );
  XNOR U4562 ( .A(n34984), .B(n34594), .Z(n34596) );
  XNOR U4563 ( .A(n34597), .B(n34201), .Z(n34203) );
  XNOR U4564 ( .A(n34204), .B(n33802), .Z(n33804) );
  XNOR U4565 ( .A(n33805), .B(n33397), .Z(n33399) );
  XNOR U4566 ( .A(n33400), .B(n32986), .Z(n32988) );
  XNOR U4567 ( .A(n32989), .B(n32569), .Z(n32571) );
  XNOR U4568 ( .A(n32572), .B(n32146), .Z(n32148) );
  XNOR U4569 ( .A(n32149), .B(n31717), .Z(n31719) );
  XNOR U4570 ( .A(n31720), .B(n31282), .Z(n31284) );
  XNOR U4571 ( .A(n31285), .B(n30841), .Z(n30843) );
  XNOR U4572 ( .A(n30844), .B(n30394), .Z(n30396) );
  XNOR U4573 ( .A(n30397), .B(n29941), .Z(n29943) );
  XNOR U4574 ( .A(n29944), .B(n29482), .Z(n29484) );
  XNOR U4575 ( .A(n29485), .B(n29017), .Z(n29019) );
  XNOR U4576 ( .A(n29020), .B(n28546), .Z(n28548) );
  XNOR U4577 ( .A(n28549), .B(n28069), .Z(n28071) );
  XNOR U4578 ( .A(n28072), .B(n27586), .Z(n27588) );
  XNOR U4579 ( .A(n27589), .B(n27097), .Z(n27099) );
  XNOR U4580 ( .A(n27100), .B(n26600), .Z(n26602) );
  XNOR U4581 ( .A(n26603), .B(n26099), .Z(n26101) );
  XNOR U4582 ( .A(n26102), .B(n25591), .Z(n25593) );
  XNOR U4583 ( .A(n25594), .B(n25077), .Z(n25079) );
  XNOR U4584 ( .A(n25080), .B(n24554), .Z(n24556) );
  XNOR U4585 ( .A(n24557), .B(n24029), .Z(n24031) );
  XNOR U4586 ( .A(n24032), .B(n23498), .Z(n23500) );
  XNOR U4587 ( .A(n23501), .B(n22960), .Z(n22962) );
  XNOR U4588 ( .A(n22963), .B(n22416), .Z(n22418) );
  XNOR U4589 ( .A(n22419), .B(n21867), .Z(n21869) );
  XNOR U4590 ( .A(n21870), .B(n21312), .Z(n21314) );
  XNOR U4591 ( .A(n21315), .B(n20750), .Z(n20752) );
  XNOR U4592 ( .A(n20753), .B(n20183), .Z(n20185) );
  XNOR U4593 ( .A(n20186), .B(n19610), .Z(n19612) );
  XNOR U4594 ( .A(n19613), .B(n19031), .Z(n19033) );
  XOR U4595 ( .A(n18339), .B(n18683), .Z(n18343) );
  XOR U4596 ( .A(n11937), .B(n12482), .Z(n11941) );
  XOR U4597 ( .A(n12550), .B(n13135), .Z(n12554) );
  XOR U4598 ( .A(n11230), .B(n11839), .Z(n11234) );
  XOR U4599 ( .A(n11872), .B(n12495), .Z(n11876) );
  XOR U4600 ( .A(n15184), .B(n15637), .Z(n15188) );
  XOR U4601 ( .A(n13914), .B(n14391), .Z(n13918) );
  XOR U4602 ( .A(n17089), .B(n17452), .Z(n17093) );
  XOR U4603 ( .A(n15855), .B(n16242), .Z(n15859) );
  XOR U4604 ( .A(n14597), .B(n15008), .Z(n14601) );
  XOR U4605 ( .A(n16520), .B(n16841), .Z(n16524) );
  XNOR U4606 ( .A(n39165), .B(n38847), .Z(n38849) );
  XOR U4607 ( .A(n9893), .B(n10520), .Z(n9897) );
  XOR U4608 ( .A(n10547), .B(n11186), .Z(n10551) );
  XOR U4609 ( .A(n9193), .B(n9856), .Z(n9197) );
  XOR U4610 ( .A(n13230), .B(n13767), .Z(n13234) );
  XOR U4611 ( .A(n11922), .B(n12485), .Z(n11926) );
  XOR U4612 ( .A(n40649), .B(n40927), .Z(n40653) );
  XOR U4613 ( .A(n40073), .B(n40351), .Z(n40077) );
  XOR U4614 ( .A(n39473), .B(n39751), .Z(n39477) );
  XOR U4615 ( .A(n17119), .B(n17446), .Z(n17123) );
  XOR U4616 ( .A(n15885), .B(n16236), .Z(n15889) );
  XOR U4617 ( .A(n14627), .B(n15002), .Z(n14631) );
  XOR U4618 ( .A(n15214), .B(n15631), .Z(n15218) );
  XOR U4619 ( .A(n13944), .B(n14385), .Z(n13948) );
  XOR U4620 ( .A(n13255), .B(n13762), .Z(n13259) );
  XOR U4621 ( .A(n7820), .B(n8501), .Z(n7824) );
  XOR U4622 ( .A(n9923), .B(n10514), .Z(n9927) );
  XNOR U4623 ( .A(n39484), .B(n39172), .Z(n39174) );
  XNOR U4624 ( .A(n39175), .B(n38857), .Z(n38859) );
  XNOR U4625 ( .A(n38860), .B(n38536), .Z(n38538) );
  XNOR U4626 ( .A(n38539), .B(n38209), .Z(n38211) );
  XNOR U4627 ( .A(n38212), .B(n37876), .Z(n37878) );
  XNOR U4628 ( .A(n37879), .B(n37537), .Z(n37539) );
  XNOR U4629 ( .A(n37540), .B(n37192), .Z(n37194) );
  XNOR U4630 ( .A(n37195), .B(n36841), .Z(n36843) );
  XNOR U4631 ( .A(n36844), .B(n36484), .Z(n36486) );
  XNOR U4632 ( .A(n36487), .B(n36121), .Z(n36123) );
  XNOR U4633 ( .A(n36124), .B(n35752), .Z(n35754) );
  XNOR U4634 ( .A(n35755), .B(n35377), .Z(n35379) );
  XNOR U4635 ( .A(n35380), .B(n34996), .Z(n34998) );
  XNOR U4636 ( .A(n34999), .B(n34609), .Z(n34611) );
  XNOR U4637 ( .A(n34612), .B(n34216), .Z(n34218) );
  XNOR U4638 ( .A(n34219), .B(n33817), .Z(n33819) );
  XNOR U4639 ( .A(n33820), .B(n33412), .Z(n33414) );
  XNOR U4640 ( .A(n33415), .B(n33001), .Z(n33003) );
  XNOR U4641 ( .A(n33004), .B(n32584), .Z(n32586) );
  XNOR U4642 ( .A(n32587), .B(n32161), .Z(n32163) );
  XNOR U4643 ( .A(n32164), .B(n31732), .Z(n31734) );
  XNOR U4644 ( .A(n31735), .B(n31297), .Z(n31299) );
  XNOR U4645 ( .A(n31300), .B(n30856), .Z(n30858) );
  XNOR U4646 ( .A(n30859), .B(n30409), .Z(n30411) );
  XNOR U4647 ( .A(n30412), .B(n29956), .Z(n29958) );
  XNOR U4648 ( .A(n29959), .B(n29497), .Z(n29499) );
  XNOR U4649 ( .A(n29500), .B(n29032), .Z(n29034) );
  XNOR U4650 ( .A(n29035), .B(n28561), .Z(n28563) );
  XNOR U4651 ( .A(n28564), .B(n28084), .Z(n28086) );
  XNOR U4652 ( .A(n28087), .B(n27601), .Z(n27603) );
  XNOR U4653 ( .A(n27604), .B(n27112), .Z(n27114) );
  XNOR U4654 ( .A(n27115), .B(n26615), .Z(n26617) );
  XNOR U4655 ( .A(n26618), .B(n26114), .Z(n26116) );
  XNOR U4656 ( .A(n26117), .B(n25606), .Z(n25608) );
  XNOR U4657 ( .A(n25609), .B(n25092), .Z(n25094) );
  XNOR U4658 ( .A(n25095), .B(n24569), .Z(n24571) );
  XNOR U4659 ( .A(n24572), .B(n24044), .Z(n24046) );
  XNOR U4660 ( .A(n24047), .B(n23513), .Z(n23515) );
  XNOR U4661 ( .A(n23516), .B(n22975), .Z(n22977) );
  XNOR U4662 ( .A(n22978), .B(n22431), .Z(n22433) );
  XNOR U4663 ( .A(n22434), .B(n21882), .Z(n21884) );
  XNOR U4664 ( .A(n21885), .B(n21327), .Z(n21329) );
  XNOR U4665 ( .A(n21330), .B(n20765), .Z(n20767) );
  XNOR U4666 ( .A(n20768), .B(n20198), .Z(n20200) );
  XNOR U4667 ( .A(n20201), .B(n19625), .Z(n19627) );
  XNOR U4668 ( .A(n19628), .B(n19046), .Z(n19048) );
  XOR U4669 ( .A(n18354), .B(n18677), .Z(n18358) );
  XOR U4670 ( .A(n17164), .B(n17437), .Z(n17168) );
  XOR U4671 ( .A(n11290), .B(n11827), .Z(n11294) );
  XOR U4672 ( .A(n9948), .B(n10509), .Z(n9952) );
  XOR U4673 ( .A(n11245), .B(n11836), .Z(n11249) );
  XOR U4674 ( .A(n13285), .B(n13756), .Z(n13289) );
  XOR U4675 ( .A(n10647), .B(n11166), .Z(n10651) );
  XOR U4676 ( .A(n15244), .B(n15625), .Z(n15248) );
  XOR U4677 ( .A(n13974), .B(n14379), .Z(n13978) );
  XOR U4678 ( .A(n17149), .B(n17440), .Z(n17153) );
  XOR U4679 ( .A(n15915), .B(n16230), .Z(n15919) );
  XOR U4680 ( .A(n14657), .B(n14996), .Z(n14661) );
  XNOR U4681 ( .A(n40089), .B(n39789), .Z(n39791) );
  XOR U4682 ( .A(n9908), .B(n10517), .Z(n9912) );
  XOR U4683 ( .A(n8542), .B(n9175), .Z(n8546) );
  XOR U4684 ( .A(n9208), .B(n9853), .Z(n9212) );
  XOR U4685 ( .A(n10607), .B(n11174), .Z(n10611) );
  XOR U4686 ( .A(n11320), .B(n11821), .Z(n11324) );
  XOR U4687 ( .A(n41483), .B(n41743), .Z(n41487) );
  XOR U4688 ( .A(n40943), .B(n41203), .Z(n40947) );
  XOR U4689 ( .A(n40379), .B(n40639), .Z(n40383) );
  XOR U4690 ( .A(n15945), .B(n16224), .Z(n15949) );
  XOR U4691 ( .A(n14687), .B(n14990), .Z(n14691) );
  XOR U4692 ( .A(n15274), .B(n15619), .Z(n15278) );
  XOR U4693 ( .A(n14004), .B(n14373), .Z(n14008) );
  XOR U4694 ( .A(n13315), .B(n13750), .Z(n13319) );
  XOR U4695 ( .A(n10677), .B(n11160), .Z(n10681) );
  XOR U4696 ( .A(n11962), .B(n12477), .Z(n11966) );
  XOR U4697 ( .A(n7835), .B(n8498), .Z(n7839) );
  XOR U4698 ( .A(n6433), .B(n7120), .Z(n6437) );
  XOR U4699 ( .A(n9258), .B(n9843), .Z(n9262) );
  XNOR U4700 ( .A(n40390), .B(n40096), .Z(n40098) );
  XNOR U4701 ( .A(n40099), .B(n39799), .Z(n39801) );
  XNOR U4702 ( .A(n39802), .B(n39496), .Z(n39498) );
  XNOR U4703 ( .A(n39499), .B(n39187), .Z(n39189) );
  XNOR U4704 ( .A(n39190), .B(n38872), .Z(n38874) );
  XNOR U4705 ( .A(n38875), .B(n38551), .Z(n38553) );
  XNOR U4706 ( .A(n38554), .B(n38224), .Z(n38226) );
  XNOR U4707 ( .A(n38227), .B(n37891), .Z(n37893) );
  XNOR U4708 ( .A(n37894), .B(n37552), .Z(n37554) );
  XNOR U4709 ( .A(n37555), .B(n37207), .Z(n37209) );
  XNOR U4710 ( .A(n37210), .B(n36856), .Z(n36858) );
  XNOR U4711 ( .A(n36859), .B(n36499), .Z(n36501) );
  XNOR U4712 ( .A(n36502), .B(n36136), .Z(n36138) );
  XNOR U4713 ( .A(n36139), .B(n35767), .Z(n35769) );
  XNOR U4714 ( .A(n35770), .B(n35392), .Z(n35394) );
  XNOR U4715 ( .A(n35395), .B(n35011), .Z(n35013) );
  XNOR U4716 ( .A(n35014), .B(n34624), .Z(n34626) );
  XNOR U4717 ( .A(n34627), .B(n34231), .Z(n34233) );
  XNOR U4718 ( .A(n34234), .B(n33832), .Z(n33834) );
  XNOR U4719 ( .A(n33835), .B(n33427), .Z(n33429) );
  XNOR U4720 ( .A(n33430), .B(n33016), .Z(n33018) );
  XNOR U4721 ( .A(n33019), .B(n32599), .Z(n32601) );
  XNOR U4722 ( .A(n32602), .B(n32176), .Z(n32178) );
  XNOR U4723 ( .A(n32179), .B(n31747), .Z(n31749) );
  XNOR U4724 ( .A(n31750), .B(n31312), .Z(n31314) );
  XNOR U4725 ( .A(n31315), .B(n30871), .Z(n30873) );
  XNOR U4726 ( .A(n30874), .B(n30424), .Z(n30426) );
  XNOR U4727 ( .A(n30427), .B(n29971), .Z(n29973) );
  XNOR U4728 ( .A(n29974), .B(n29512), .Z(n29514) );
  XNOR U4729 ( .A(n29515), .B(n29047), .Z(n29049) );
  XNOR U4730 ( .A(n29050), .B(n28576), .Z(n28578) );
  XNOR U4731 ( .A(n28579), .B(n28099), .Z(n28101) );
  XNOR U4732 ( .A(n28102), .B(n27616), .Z(n27618) );
  XNOR U4733 ( .A(n27619), .B(n27127), .Z(n27129) );
  XNOR U4734 ( .A(n27130), .B(n26630), .Z(n26632) );
  XNOR U4735 ( .A(n26633), .B(n26129), .Z(n26131) );
  XNOR U4736 ( .A(n26132), .B(n25621), .Z(n25623) );
  XNOR U4737 ( .A(n25624), .B(n25107), .Z(n25109) );
  XNOR U4738 ( .A(n25110), .B(n24584), .Z(n24586) );
  XNOR U4739 ( .A(n24587), .B(n24059), .Z(n24061) );
  XNOR U4740 ( .A(n24062), .B(n23528), .Z(n23530) );
  XNOR U4741 ( .A(n23531), .B(n22990), .Z(n22992) );
  XNOR U4742 ( .A(n22993), .B(n22446), .Z(n22448) );
  XNOR U4743 ( .A(n22449), .B(n21897), .Z(n21899) );
  XNOR U4744 ( .A(n21900), .B(n21342), .Z(n21344) );
  XNOR U4745 ( .A(n21345), .B(n20780), .Z(n20782) );
  XNOR U4746 ( .A(n20783), .B(n20213), .Z(n20215) );
  XNOR U4747 ( .A(n20216), .B(n19640), .Z(n19642) );
  XNOR U4748 ( .A(n19643), .B(n19061), .Z(n19063) );
  XOR U4749 ( .A(n17777), .B(n18032), .Z(n17781) );
  XOR U4750 ( .A(n11350), .B(n11815), .Z(n11354) );
  XOR U4751 ( .A(n9283), .B(n9838), .Z(n9287) );
  XOR U4752 ( .A(n5010), .B(n5717), .Z(n5014) );
  XOR U4753 ( .A(n7187), .B(n7802), .Z(n7191) );
  XOR U4754 ( .A(n11992), .B(n12471), .Z(n11996) );
  XOR U4755 ( .A(n13345), .B(n13744), .Z(n13349) );
  XOR U4756 ( .A(n10707), .B(n11154), .Z(n10711) );
  XOR U4757 ( .A(n15304), .B(n15613), .Z(n15308) );
  XOR U4758 ( .A(n14034), .B(n14367), .Z(n14038) );
  XOR U4759 ( .A(n14717), .B(n14984), .Z(n14721) );
  XNOR U4760 ( .A(n40959), .B(n40677), .Z(n40679) );
  XOR U4761 ( .A(n9968), .B(n10505), .Z(n9972) );
  XOR U4762 ( .A(n8557), .B(n9172), .Z(n8561) );
  XOR U4763 ( .A(n5753), .B(n6416), .Z(n5757) );
  XOR U4764 ( .A(n9313), .B(n9832), .Z(n9317) );
  XOR U4765 ( .A(n11380), .B(n11809), .Z(n11384) );
  XOR U4766 ( .A(n42263), .B(n42505), .Z(n42267) );
  XOR U4767 ( .A(n41759), .B(n42001), .Z(n41763) );
  XOR U4768 ( .A(n41231), .B(n41473), .Z(n41235) );
  XOR U4769 ( .A(n15334), .B(n15607), .Z(n15338) );
  XOR U4770 ( .A(n14064), .B(n14361), .Z(n14068) );
  XOR U4771 ( .A(n13375), .B(n13738), .Z(n13379) );
  XOR U4772 ( .A(n10737), .B(n11148), .Z(n10741) );
  XOR U4773 ( .A(n12022), .B(n12465), .Z(n12026) );
  XOR U4774 ( .A(n7217), .B(n7796), .Z(n7221) );
  XOR U4775 ( .A(n6468), .B(n7113), .Z(n6472) );
  XOR U4776 ( .A(n6448), .B(n7117), .Z(n6452) );
  XOR U4777 ( .A(n8587), .B(n9166), .Z(n8591) );
  XOR U4778 ( .A(n9998), .B(n10499), .Z(n10002) );
  XNOR U4779 ( .A(n41242), .B(n40966), .Z(n40968) );
  XNOR U4780 ( .A(n40969), .B(n40687), .Z(n40689) );
  XNOR U4781 ( .A(n40690), .B(n40402), .Z(n40404) );
  XNOR U4782 ( .A(n40405), .B(n40111), .Z(n40113) );
  XNOR U4783 ( .A(n40114), .B(n39814), .Z(n39816) );
  XNOR U4784 ( .A(n39817), .B(n39511), .Z(n39513) );
  XNOR U4785 ( .A(n39514), .B(n39202), .Z(n39204) );
  XNOR U4786 ( .A(n39205), .B(n38887), .Z(n38889) );
  XNOR U4787 ( .A(n38890), .B(n38566), .Z(n38568) );
  XNOR U4788 ( .A(n38569), .B(n38239), .Z(n38241) );
  XNOR U4789 ( .A(n38242), .B(n37906), .Z(n37908) );
  XNOR U4790 ( .A(n37909), .B(n37567), .Z(n37569) );
  XNOR U4791 ( .A(n37570), .B(n37222), .Z(n37224) );
  XNOR U4792 ( .A(n37225), .B(n36871), .Z(n36873) );
  XNOR U4793 ( .A(n36874), .B(n36514), .Z(n36516) );
  XNOR U4794 ( .A(n36517), .B(n36151), .Z(n36153) );
  XNOR U4795 ( .A(n36154), .B(n35782), .Z(n35784) );
  XNOR U4796 ( .A(n35785), .B(n35407), .Z(n35409) );
  XNOR U4797 ( .A(n35410), .B(n35026), .Z(n35028) );
  XNOR U4798 ( .A(n35029), .B(n34639), .Z(n34641) );
  XNOR U4799 ( .A(n34642), .B(n34246), .Z(n34248) );
  XNOR U4800 ( .A(n34249), .B(n33847), .Z(n33849) );
  XNOR U4801 ( .A(n33850), .B(n33442), .Z(n33444) );
  XNOR U4802 ( .A(n33445), .B(n33031), .Z(n33033) );
  XNOR U4803 ( .A(n33034), .B(n32614), .Z(n32616) );
  XNOR U4804 ( .A(n32617), .B(n32191), .Z(n32193) );
  XNOR U4805 ( .A(n32194), .B(n31762), .Z(n31764) );
  XNOR U4806 ( .A(n31765), .B(n31327), .Z(n31329) );
  XNOR U4807 ( .A(n31330), .B(n30886), .Z(n30888) );
  XNOR U4808 ( .A(n30889), .B(n30439), .Z(n30441) );
  XNOR U4809 ( .A(n30442), .B(n29986), .Z(n29988) );
  XNOR U4810 ( .A(n29989), .B(n29527), .Z(n29529) );
  XNOR U4811 ( .A(n29530), .B(n29062), .Z(n29064) );
  XNOR U4812 ( .A(n29065), .B(n28591), .Z(n28593) );
  XNOR U4813 ( .A(n28594), .B(n28114), .Z(n28116) );
  XNOR U4814 ( .A(n28117), .B(n27631), .Z(n27633) );
  XNOR U4815 ( .A(n27634), .B(n27142), .Z(n27144) );
  XNOR U4816 ( .A(n27145), .B(n26645), .Z(n26647) );
  XNOR U4817 ( .A(n26648), .B(n26144), .Z(n26146) );
  XNOR U4818 ( .A(n26147), .B(n25636), .Z(n25638) );
  XNOR U4819 ( .A(n25639), .B(n25122), .Z(n25124) );
  XNOR U4820 ( .A(n25125), .B(n24599), .Z(n24601) );
  XNOR U4821 ( .A(n24602), .B(n24074), .Z(n24076) );
  XNOR U4822 ( .A(n24077), .B(n23543), .Z(n23545) );
  XNOR U4823 ( .A(n23546), .B(n23005), .Z(n23007) );
  XNOR U4824 ( .A(n23008), .B(n22461), .Z(n22463) );
  XNOR U4825 ( .A(n22464), .B(n21912), .Z(n21914) );
  XNOR U4826 ( .A(n21915), .B(n21357), .Z(n21359) );
  XNOR U4827 ( .A(n21360), .B(n20795), .Z(n20797) );
  XNOR U4828 ( .A(n20798), .B(n20228), .Z(n20230) );
  XNOR U4829 ( .A(n20231), .B(n19655), .Z(n19657) );
  XNOR U4830 ( .A(n19658), .B(n19076), .Z(n19078) );
  XOR U4831 ( .A(n17792), .B(n18029), .Z(n17796) );
  XOR U4832 ( .A(n16590), .B(n16827), .Z(n16594) );
  XOR U4833 ( .A(n14114), .B(n14351), .Z(n14118) );
  XOR U4834 ( .A(n11410), .B(n11803), .Z(n11414) );
  XOR U4835 ( .A(n9343), .B(n9826), .Z(n9347) );
  XOR U4836 ( .A(n5025), .B(n5714), .Z(n5029) );
  XOR U4837 ( .A(n3575), .B(n4286), .Z(n3579) );
  XOR U4838 ( .A(n7202), .B(n7799), .Z(n7206) );
  XOR U4839 ( .A(n7247), .B(n7790), .Z(n7251) );
  XOR U4840 ( .A(n12052), .B(n12459), .Z(n12056) );
  XOR U4841 ( .A(n13405), .B(n13732), .Z(n13409) );
  XOR U4842 ( .A(n10767), .B(n11142), .Z(n10771) );
  XOR U4843 ( .A(n15364), .B(n15601), .Z(n15368) );
  XOR U4844 ( .A(n14094), .B(n14355), .Z(n14098) );
  XNOR U4845 ( .A(n41775), .B(n41511), .Z(n41513) );
  XOR U4846 ( .A(n10028), .B(n10493), .Z(n10032) );
  XOR U4847 ( .A(n8617), .B(n9160), .Z(n8621) );
  XOR U4848 ( .A(n4328), .B(n4997), .Z(n4332) );
  XOR U4849 ( .A(n9373), .B(n9820), .Z(n9377) );
  XOR U4850 ( .A(n11440), .B(n11797), .Z(n11444) );
  XOR U4851 ( .A(n42989), .B(n43213), .Z(n42993) );
  XOR U4852 ( .A(n42521), .B(n42745), .Z(n42525) );
  XOR U4853 ( .A(n42029), .B(n42253), .Z(n42033) );
  XOR U4854 ( .A(n13435), .B(n13726), .Z(n13439) );
  XOR U4855 ( .A(n10797), .B(n11136), .Z(n10801) );
  XOR U4856 ( .A(n12082), .B(n12453), .Z(n12086) );
  XOR U4857 ( .A(n7277), .B(n7784), .Z(n7281) );
  XOR U4858 ( .A(n7232), .B(n7793), .Z(n7236) );
  XOR U4859 ( .A(n5773), .B(n6412), .Z(n5777) );
  XOR U4860 ( .A(n5080), .B(n5703), .Z(n5084) );
  XOR U4861 ( .A(n3630), .B(n4275), .Z(n3634) );
  XOR U4862 ( .A(n8647), .B(n9154), .Z(n8651) );
  XOR U4863 ( .A(n10058), .B(n10487), .Z(n10062) );
  XNOR U4864 ( .A(n42040), .B(n41782), .Z(n41784) );
  XNOR U4865 ( .A(n41785), .B(n41521), .Z(n41523) );
  XNOR U4866 ( .A(n41524), .B(n41254), .Z(n41256) );
  XNOR U4867 ( .A(n41257), .B(n40981), .Z(n40983) );
  XNOR U4868 ( .A(n40984), .B(n40702), .Z(n40704) );
  XNOR U4869 ( .A(n40705), .B(n40417), .Z(n40419) );
  XNOR U4870 ( .A(n40420), .B(n40126), .Z(n40128) );
  XNOR U4871 ( .A(n40129), .B(n39829), .Z(n39831) );
  XNOR U4872 ( .A(n39832), .B(n39526), .Z(n39528) );
  XNOR U4873 ( .A(n39529), .B(n39217), .Z(n39219) );
  XNOR U4874 ( .A(n39220), .B(n38902), .Z(n38904) );
  XNOR U4875 ( .A(n38905), .B(n38581), .Z(n38583) );
  XNOR U4876 ( .A(n38584), .B(n38254), .Z(n38256) );
  XNOR U4877 ( .A(n38257), .B(n37921), .Z(n37923) );
  XNOR U4878 ( .A(n37924), .B(n37582), .Z(n37584) );
  XNOR U4879 ( .A(n37585), .B(n37237), .Z(n37239) );
  XNOR U4880 ( .A(n37240), .B(n36886), .Z(n36888) );
  XNOR U4881 ( .A(n36889), .B(n36529), .Z(n36531) );
  XNOR U4882 ( .A(n36532), .B(n36166), .Z(n36168) );
  XNOR U4883 ( .A(n36169), .B(n35797), .Z(n35799) );
  XNOR U4884 ( .A(n35800), .B(n35422), .Z(n35424) );
  XNOR U4885 ( .A(n35425), .B(n35041), .Z(n35043) );
  XNOR U4886 ( .A(n35044), .B(n34654), .Z(n34656) );
  XNOR U4887 ( .A(n34657), .B(n34261), .Z(n34263) );
  XNOR U4888 ( .A(n34264), .B(n33862), .Z(n33864) );
  XNOR U4889 ( .A(n33865), .B(n33457), .Z(n33459) );
  XNOR U4890 ( .A(n33460), .B(n33046), .Z(n33048) );
  XNOR U4891 ( .A(n33049), .B(n32629), .Z(n32631) );
  XNOR U4892 ( .A(n32632), .B(n32206), .Z(n32208) );
  XNOR U4893 ( .A(n32209), .B(n31777), .Z(n31779) );
  XNOR U4894 ( .A(n31780), .B(n31342), .Z(n31344) );
  XNOR U4895 ( .A(n31345), .B(n30901), .Z(n30903) );
  XNOR U4896 ( .A(n30904), .B(n30454), .Z(n30456) );
  XNOR U4897 ( .A(n30457), .B(n30001), .Z(n30003) );
  XNOR U4898 ( .A(n30004), .B(n29542), .Z(n29544) );
  XNOR U4899 ( .A(n29545), .B(n29077), .Z(n29079) );
  XNOR U4900 ( .A(n29080), .B(n28606), .Z(n28608) );
  XNOR U4901 ( .A(n28609), .B(n28129), .Z(n28131) );
  XNOR U4902 ( .A(n28132), .B(n27646), .Z(n27648) );
  XNOR U4903 ( .A(n27649), .B(n27157), .Z(n27159) );
  XNOR U4904 ( .A(n27160), .B(n26660), .Z(n26662) );
  XNOR U4905 ( .A(n26663), .B(n26159), .Z(n26161) );
  XNOR U4906 ( .A(n26162), .B(n25651), .Z(n25653) );
  XNOR U4907 ( .A(n25654), .B(n25137), .Z(n25139) );
  XNOR U4908 ( .A(n25140), .B(n24614), .Z(n24616) );
  XNOR U4909 ( .A(n24617), .B(n24089), .Z(n24091) );
  XNOR U4910 ( .A(n24092), .B(n23558), .Z(n23560) );
  XNOR U4911 ( .A(n23561), .B(n23020), .Z(n23022) );
  XNOR U4912 ( .A(n23023), .B(n22476), .Z(n22478) );
  XNOR U4913 ( .A(n22479), .B(n21927), .Z(n21929) );
  XNOR U4914 ( .A(n21930), .B(n21372), .Z(n21374) );
  XNOR U4915 ( .A(n21375), .B(n20810), .Z(n20812) );
  XNOR U4916 ( .A(n20813), .B(n20243), .Z(n20245) );
  XNOR U4917 ( .A(n20246), .B(n19670), .Z(n19672) );
  XNOR U4918 ( .A(n19673), .B(n19091), .Z(n19093) );
  XOR U4919 ( .A(n17807), .B(n18026), .Z(n17811) );
  XOR U4920 ( .A(n16605), .B(n16824), .Z(n16609) );
  XOR U4921 ( .A(n15379), .B(n15598), .Z(n15383) );
  XOR U4922 ( .A(n11470), .B(n11791), .Z(n11474) );
  XOR U4923 ( .A(n9403), .B(n9814), .Z(n9407) );
  XOR U4924 ( .A(n1390), .B(n2095), .Z(n1394) );
  XOR U4925 ( .A(n3590), .B(n4283), .Z(n3594) );
  XOR U4926 ( .A(n5803), .B(n6406), .Z(n5807) );
  XOR U4927 ( .A(n7262), .B(n7787), .Z(n7266) );
  XOR U4928 ( .A(n7307), .B(n7778), .Z(n7311) );
  XOR U4929 ( .A(n12112), .B(n12447), .Z(n12116) );
  XOR U4930 ( .A(n13465), .B(n13720), .Z(n13469) );
  XOR U4931 ( .A(n10827), .B(n11130), .Z(n10831) );
  XNOR U4932 ( .A(n42537), .B(n42291), .Z(n42293) );
  XOR U4933 ( .A(n10088), .B(n10481), .Z(n10092) );
  XOR U4934 ( .A(n8677), .B(n9148), .Z(n8681) );
  XOR U4935 ( .A(n5110), .B(n5697), .Z(n5114) );
  XOR U4936 ( .A(n3660), .B(n4269), .Z(n3664) );
  XOR U4937 ( .A(n3615), .B(n4278), .Z(n3619) );
  XOR U4938 ( .A(n2141), .B(n2828), .Z(n2145) );
  XOR U4939 ( .A(n2121), .B(n2832), .Z(n2125) );
  XOR U4940 ( .A(n9433), .B(n9808), .Z(n9437) );
  XOR U4941 ( .A(n11500), .B(n11785), .Z(n11504) );
  XOR U4942 ( .A(n43661), .B(n43867), .Z(n43665) );
  XOR U4943 ( .A(n43229), .B(n43435), .Z(n43233) );
  XOR U4944 ( .A(n42773), .B(n42979), .Z(n42777) );
  XOR U4945 ( .A(n13495), .B(n13714), .Z(n13499) );
  XOR U4946 ( .A(n10857), .B(n11124), .Z(n10861) );
  XOR U4947 ( .A(n12142), .B(n12441), .Z(n12146) );
  XOR U4948 ( .A(n7337), .B(n7772), .Z(n7341) );
  XOR U4949 ( .A(n7292), .B(n7781), .Z(n7296) );
  XOR U4950 ( .A(n5833), .B(n6400), .Z(n5837) );
  XOR U4951 ( .A(n3645), .B(n4272), .Z(n3649) );
  XOR U4952 ( .A(n2171), .B(n2822), .Z(n2175) );
  XOR U4953 ( .A(n5140), .B(n5691), .Z(n5144) );
  XOR U4954 ( .A(n3690), .B(n4263), .Z(n3694) );
  XOR U4955 ( .A(n8707), .B(n9142), .Z(n8711) );
  XOR U4956 ( .A(n10118), .B(n10475), .Z(n10122) );
  XNOR U4957 ( .A(n42784), .B(n42544), .Z(n42546) );
  XNOR U4958 ( .A(n42547), .B(n42301), .Z(n42303) );
  XNOR U4959 ( .A(n42304), .B(n42052), .Z(n42054) );
  XNOR U4960 ( .A(n42055), .B(n41797), .Z(n41799) );
  XNOR U4961 ( .A(n41800), .B(n41536), .Z(n41538) );
  XNOR U4962 ( .A(n41539), .B(n41269), .Z(n41271) );
  XNOR U4963 ( .A(n41272), .B(n40996), .Z(n40998) );
  XNOR U4964 ( .A(n40999), .B(n40717), .Z(n40719) );
  XNOR U4965 ( .A(n40720), .B(n40432), .Z(n40434) );
  XNOR U4966 ( .A(n40435), .B(n40141), .Z(n40143) );
  XNOR U4967 ( .A(n40144), .B(n39844), .Z(n39846) );
  XNOR U4968 ( .A(n39847), .B(n39541), .Z(n39543) );
  XNOR U4969 ( .A(n39544), .B(n39232), .Z(n39234) );
  XNOR U4970 ( .A(n39235), .B(n38917), .Z(n38919) );
  XNOR U4971 ( .A(n38920), .B(n38596), .Z(n38598) );
  XNOR U4972 ( .A(n38599), .B(n38269), .Z(n38271) );
  XNOR U4973 ( .A(n38272), .B(n37936), .Z(n37938) );
  XNOR U4974 ( .A(n37939), .B(n37597), .Z(n37599) );
  XNOR U4975 ( .A(n37600), .B(n37252), .Z(n37254) );
  XNOR U4976 ( .A(n37255), .B(n36901), .Z(n36903) );
  XNOR U4977 ( .A(n36904), .B(n36544), .Z(n36546) );
  XNOR U4978 ( .A(n36547), .B(n36181), .Z(n36183) );
  XNOR U4979 ( .A(n36184), .B(n35812), .Z(n35814) );
  XNOR U4980 ( .A(n35815), .B(n35437), .Z(n35439) );
  XNOR U4981 ( .A(n35440), .B(n35056), .Z(n35058) );
  XNOR U4982 ( .A(n35059), .B(n34669), .Z(n34671) );
  XNOR U4983 ( .A(n34672), .B(n34276), .Z(n34278) );
  XNOR U4984 ( .A(n34279), .B(n33877), .Z(n33879) );
  XNOR U4985 ( .A(n33880), .B(n33472), .Z(n33474) );
  XNOR U4986 ( .A(n33475), .B(n33061), .Z(n33063) );
  XNOR U4987 ( .A(n33064), .B(n32644), .Z(n32646) );
  XNOR U4988 ( .A(n32647), .B(n32221), .Z(n32223) );
  XNOR U4989 ( .A(n32224), .B(n31792), .Z(n31794) );
  XNOR U4990 ( .A(n31795), .B(n31357), .Z(n31359) );
  XNOR U4991 ( .A(n31360), .B(n30916), .Z(n30918) );
  XNOR U4992 ( .A(n30919), .B(n30469), .Z(n30471) );
  XNOR U4993 ( .A(n30472), .B(n30016), .Z(n30018) );
  XNOR U4994 ( .A(n30019), .B(n29557), .Z(n29559) );
  XNOR U4995 ( .A(n29560), .B(n29092), .Z(n29094) );
  XNOR U4996 ( .A(n29095), .B(n28621), .Z(n28623) );
  XNOR U4997 ( .A(n28624), .B(n28144), .Z(n28146) );
  XNOR U4998 ( .A(n28147), .B(n27661), .Z(n27663) );
  XNOR U4999 ( .A(n27664), .B(n27172), .Z(n27174) );
  XNOR U5000 ( .A(n27175), .B(n26675), .Z(n26677) );
  XNOR U5001 ( .A(n26678), .B(n26174), .Z(n26176) );
  XNOR U5002 ( .A(n26177), .B(n25666), .Z(n25668) );
  XNOR U5003 ( .A(n25669), .B(n25152), .Z(n25154) );
  XNOR U5004 ( .A(n25155), .B(n24629), .Z(n24631) );
  XNOR U5005 ( .A(n24632), .B(n24104), .Z(n24106) );
  XNOR U5006 ( .A(n24107), .B(n23573), .Z(n23575) );
  XNOR U5007 ( .A(n23576), .B(n23035), .Z(n23037) );
  XNOR U5008 ( .A(n23038), .B(n22491), .Z(n22493) );
  XNOR U5009 ( .A(n22494), .B(n21942), .Z(n21944) );
  XNOR U5010 ( .A(n21945), .B(n21387), .Z(n21389) );
  XNOR U5011 ( .A(n21390), .B(n20825), .Z(n20827) );
  XNOR U5012 ( .A(n20828), .B(n20258), .Z(n20260) );
  XNOR U5013 ( .A(n20261), .B(n19685), .Z(n19687) );
  XNOR U5014 ( .A(n19688), .B(n19106), .Z(n19108) );
  XOR U5015 ( .A(n18414), .B(n18653), .Z(n18418) );
  XOR U5016 ( .A(n17224), .B(n17425), .Z(n17228) );
  XOR U5017 ( .A(n16010), .B(n16211), .Z(n16014) );
  XOR U5018 ( .A(n14772), .B(n14973), .Z(n14776) );
  XOR U5019 ( .A(n13510), .B(n13711), .Z(n13514) );
  XOR U5020 ( .A(n11530), .B(n11779), .Z(n11534) );
  XOR U5021 ( .A(n9463), .B(n9802), .Z(n9467) );
  XOR U5022 ( .A(n5863), .B(n6394), .Z(n5867) );
  XOR U5023 ( .A(n7322), .B(n7775), .Z(n7326) );
  XOR U5024 ( .A(n7367), .B(n7766), .Z(n7371) );
  XOR U5025 ( .A(n12172), .B(n12435), .Z(n12176) );
  XOR U5026 ( .A(n10887), .B(n11118), .Z(n10891) );
  XNOR U5027 ( .A(n43245), .B(n43017), .Z(n43019) );
  XOR U5028 ( .A(n10148), .B(n10469), .Z(n10152) );
  XOR U5029 ( .A(n8737), .B(n9136), .Z(n8741) );
  XOR U5030 ( .A(n5170), .B(n5685), .Z(n5174) );
  XOR U5031 ( .A(n3720), .B(n4257), .Z(n3724) );
  XOR U5032 ( .A(n3675), .B(n4266), .Z(n3679) );
  XOR U5033 ( .A(n2201), .B(n2816), .Z(n2205) );
  XOR U5034 ( .A(n2156), .B(n2825), .Z(n2160) );
  XOR U5035 ( .A(n9493), .B(n9796), .Z(n9497) );
  XOR U5036 ( .A(n11560), .B(n11773), .Z(n11564) );
  XOR U5037 ( .A(n44279), .B(n44467), .Z(n44283) );
  XOR U5038 ( .A(n43883), .B(n44071), .Z(n43887) );
  XOR U5039 ( .A(n43463), .B(n43651), .Z(n43467) );
  XOR U5040 ( .A(n12202), .B(n12429), .Z(n12206) );
  XOR U5041 ( .A(n7397), .B(n7760), .Z(n7401) );
  XOR U5042 ( .A(n7352), .B(n7769), .Z(n7356) );
  XOR U5043 ( .A(n5893), .B(n6388), .Z(n5897) );
  XOR U5044 ( .A(n2186), .B(n2819), .Z(n2190) );
  XOR U5045 ( .A(n3705), .B(n4260), .Z(n3709) );
  XOR U5046 ( .A(n2231), .B(n2810), .Z(n2235) );
  XOR U5047 ( .A(n5200), .B(n5679), .Z(n5204) );
  XOR U5048 ( .A(n3750), .B(n4251), .Z(n3754) );
  XOR U5049 ( .A(n8767), .B(n9130), .Z(n8771) );
  XOR U5050 ( .A(n10178), .B(n10463), .Z(n10182) );
  XNOR U5051 ( .A(n43474), .B(n43252), .Z(n43254) );
  XNOR U5052 ( .A(n43255), .B(n43027), .Z(n43029) );
  XNOR U5053 ( .A(n43030), .B(n42796), .Z(n42798) );
  XNOR U5054 ( .A(n42799), .B(n42559), .Z(n42561) );
  XNOR U5055 ( .A(n42562), .B(n42316), .Z(n42318) );
  XNOR U5056 ( .A(n42319), .B(n42067), .Z(n42069) );
  XNOR U5057 ( .A(n42070), .B(n41812), .Z(n41814) );
  XNOR U5058 ( .A(n41815), .B(n41551), .Z(n41553) );
  XNOR U5059 ( .A(n41554), .B(n41284), .Z(n41286) );
  XNOR U5060 ( .A(n41287), .B(n41011), .Z(n41013) );
  XNOR U5061 ( .A(n41014), .B(n40732), .Z(n40734) );
  XNOR U5062 ( .A(n40735), .B(n40447), .Z(n40449) );
  XNOR U5063 ( .A(n40450), .B(n40156), .Z(n40158) );
  XNOR U5064 ( .A(n40159), .B(n39859), .Z(n39861) );
  XNOR U5065 ( .A(n39862), .B(n39556), .Z(n39558) );
  XNOR U5066 ( .A(n39559), .B(n39247), .Z(n39249) );
  XNOR U5067 ( .A(n39250), .B(n38932), .Z(n38934) );
  XNOR U5068 ( .A(n38935), .B(n38611), .Z(n38613) );
  XNOR U5069 ( .A(n38614), .B(n38284), .Z(n38286) );
  XNOR U5070 ( .A(n38287), .B(n37951), .Z(n37953) );
  XNOR U5071 ( .A(n37954), .B(n37612), .Z(n37614) );
  XNOR U5072 ( .A(n37615), .B(n37267), .Z(n37269) );
  XNOR U5073 ( .A(n37270), .B(n36916), .Z(n36918) );
  XNOR U5074 ( .A(n36919), .B(n36559), .Z(n36561) );
  XNOR U5075 ( .A(n36562), .B(n36196), .Z(n36198) );
  XNOR U5076 ( .A(n36199), .B(n35827), .Z(n35829) );
  XNOR U5077 ( .A(n35830), .B(n35452), .Z(n35454) );
  XNOR U5078 ( .A(n35455), .B(n35071), .Z(n35073) );
  XNOR U5079 ( .A(n35074), .B(n34684), .Z(n34686) );
  XNOR U5080 ( .A(n34687), .B(n34291), .Z(n34293) );
  XNOR U5081 ( .A(n34294), .B(n33892), .Z(n33894) );
  XNOR U5082 ( .A(n33895), .B(n33487), .Z(n33489) );
  XNOR U5083 ( .A(n33490), .B(n33076), .Z(n33078) );
  XNOR U5084 ( .A(n33079), .B(n32659), .Z(n32661) );
  XNOR U5085 ( .A(n32662), .B(n32236), .Z(n32238) );
  XNOR U5086 ( .A(n32239), .B(n31807), .Z(n31809) );
  XNOR U5087 ( .A(n31810), .B(n31372), .Z(n31374) );
  XNOR U5088 ( .A(n31375), .B(n30931), .Z(n30933) );
  XNOR U5089 ( .A(n30934), .B(n30484), .Z(n30486) );
  XNOR U5090 ( .A(n30487), .B(n30031), .Z(n30033) );
  XNOR U5091 ( .A(n30034), .B(n29572), .Z(n29574) );
  XNOR U5092 ( .A(n29575), .B(n29107), .Z(n29109) );
  XNOR U5093 ( .A(n29110), .B(n28636), .Z(n28638) );
  XNOR U5094 ( .A(n28639), .B(n28159), .Z(n28161) );
  XNOR U5095 ( .A(n28162), .B(n27676), .Z(n27678) );
  XNOR U5096 ( .A(n27679), .B(n27187), .Z(n27189) );
  XNOR U5097 ( .A(n27190), .B(n26690), .Z(n26692) );
  XNOR U5098 ( .A(n26693), .B(n26189), .Z(n26191) );
  XNOR U5099 ( .A(n26192), .B(n25681), .Z(n25683) );
  XNOR U5100 ( .A(n25684), .B(n25167), .Z(n25169) );
  XNOR U5101 ( .A(n25170), .B(n24644), .Z(n24646) );
  XNOR U5102 ( .A(n24647), .B(n24119), .Z(n24121) );
  XNOR U5103 ( .A(n24122), .B(n23588), .Z(n23590) );
  XNOR U5104 ( .A(n23591), .B(n23050), .Z(n23052) );
  XNOR U5105 ( .A(n23053), .B(n22506), .Z(n22508) );
  XNOR U5106 ( .A(n22509), .B(n21957), .Z(n21959) );
  XNOR U5107 ( .A(n21960), .B(n21402), .Z(n21404) );
  XNOR U5108 ( .A(n21405), .B(n20840), .Z(n20842) );
  XNOR U5109 ( .A(n20843), .B(n20273), .Z(n20275) );
  XNOR U5110 ( .A(n20276), .B(n19700), .Z(n19702) );
  XNOR U5111 ( .A(n19703), .B(n19121), .Z(n19123) );
  XOR U5112 ( .A(n18429), .B(n18647), .Z(n18433) );
  XOR U5113 ( .A(n17239), .B(n17422), .Z(n17243) );
  XOR U5114 ( .A(n16025), .B(n16208), .Z(n16029) );
  XOR U5115 ( .A(n14787), .B(n14970), .Z(n14791) );
  XOR U5116 ( .A(n13525), .B(n13708), .Z(n13529) );
  XOR U5117 ( .A(n11585), .B(n11768), .Z(n11589) );
  XOR U5118 ( .A(n9523), .B(n9790), .Z(n9527) );
  XOR U5119 ( .A(n5923), .B(n6382), .Z(n5927) );
  XOR U5120 ( .A(n7382), .B(n7763), .Z(n7386) );
  XOR U5121 ( .A(n7427), .B(n7754), .Z(n7431) );
  XOR U5122 ( .A(n12232), .B(n12423), .Z(n12236) );
  XNOR U5123 ( .A(n43899), .B(n43689), .Z(n43691) );
  XOR U5124 ( .A(n10208), .B(n10457), .Z(n10212) );
  XOR U5125 ( .A(n8797), .B(n9124), .Z(n8801) );
  XOR U5126 ( .A(n5230), .B(n5673), .Z(n5234) );
  XOR U5127 ( .A(n3780), .B(n4245), .Z(n3784) );
  XOR U5128 ( .A(n3735), .B(n4254), .Z(n3739) );
  XOR U5129 ( .A(n2261), .B(n2804), .Z(n2265) );
  XOR U5130 ( .A(n2216), .B(n2813), .Z(n2220) );
  XOR U5131 ( .A(n9553), .B(n9784), .Z(n9557) );
  XOR U5132 ( .A(n44843), .B(n45013), .Z(n44847) );
  XOR U5133 ( .A(n44483), .B(n44653), .Z(n44487) );
  XOR U5134 ( .A(n44099), .B(n44269), .Z(n44103) );
  XOR U5135 ( .A(n7457), .B(n7748), .Z(n7461) );
  XOR U5136 ( .A(n7412), .B(n7757), .Z(n7416) );
  XOR U5137 ( .A(n5953), .B(n6376), .Z(n5957) );
  XOR U5138 ( .A(n2246), .B(n2807), .Z(n2250) );
  XOR U5139 ( .A(n3765), .B(n4248), .Z(n3769) );
  XOR U5140 ( .A(n2291), .B(n2798), .Z(n2295) );
  XOR U5141 ( .A(n5260), .B(n5667), .Z(n5264) );
  XOR U5142 ( .A(n3810), .B(n4239), .Z(n3814) );
  XOR U5143 ( .A(n8827), .B(n9118), .Z(n8831) );
  XOR U5144 ( .A(n10238), .B(n10451), .Z(n10242) );
  XNOR U5145 ( .A(n44110), .B(n43906), .Z(n43908) );
  XNOR U5146 ( .A(n43909), .B(n43699), .Z(n43701) );
  XNOR U5147 ( .A(n43702), .B(n43486), .Z(n43488) );
  XNOR U5148 ( .A(n43489), .B(n43267), .Z(n43269) );
  XNOR U5149 ( .A(n43270), .B(n43042), .Z(n43044) );
  XNOR U5150 ( .A(n43045), .B(n42811), .Z(n42813) );
  XNOR U5151 ( .A(n42814), .B(n42574), .Z(n42576) );
  XNOR U5152 ( .A(n42577), .B(n42331), .Z(n42333) );
  XNOR U5153 ( .A(n42334), .B(n42082), .Z(n42084) );
  XNOR U5154 ( .A(n42085), .B(n41827), .Z(n41829) );
  XNOR U5155 ( .A(n41830), .B(n41566), .Z(n41568) );
  XNOR U5156 ( .A(n41569), .B(n41299), .Z(n41301) );
  XNOR U5157 ( .A(n41302), .B(n41026), .Z(n41028) );
  XNOR U5158 ( .A(n41029), .B(n40747), .Z(n40749) );
  XNOR U5159 ( .A(n40750), .B(n40462), .Z(n40464) );
  XNOR U5160 ( .A(n40465), .B(n40171), .Z(n40173) );
  XNOR U5161 ( .A(n40174), .B(n39874), .Z(n39876) );
  XNOR U5162 ( .A(n39877), .B(n39571), .Z(n39573) );
  XNOR U5163 ( .A(n39574), .B(n39262), .Z(n39264) );
  XNOR U5164 ( .A(n39265), .B(n38947), .Z(n38949) );
  XNOR U5165 ( .A(n38950), .B(n38626), .Z(n38628) );
  XNOR U5166 ( .A(n38629), .B(n38299), .Z(n38301) );
  XNOR U5167 ( .A(n38302), .B(n37966), .Z(n37968) );
  XNOR U5168 ( .A(n37969), .B(n37627), .Z(n37629) );
  XNOR U5169 ( .A(n37630), .B(n37282), .Z(n37284) );
  XNOR U5170 ( .A(n37285), .B(n36931), .Z(n36933) );
  XNOR U5171 ( .A(n36934), .B(n36574), .Z(n36576) );
  XNOR U5172 ( .A(n36577), .B(n36211), .Z(n36213) );
  XNOR U5173 ( .A(n36214), .B(n35842), .Z(n35844) );
  XNOR U5174 ( .A(n35845), .B(n35467), .Z(n35469) );
  XNOR U5175 ( .A(n35470), .B(n35086), .Z(n35088) );
  XNOR U5176 ( .A(n35089), .B(n34699), .Z(n34701) );
  XNOR U5177 ( .A(n34702), .B(n34306), .Z(n34308) );
  XNOR U5178 ( .A(n34309), .B(n33907), .Z(n33909) );
  XNOR U5179 ( .A(n33910), .B(n33502), .Z(n33504) );
  XNOR U5180 ( .A(n33505), .B(n33091), .Z(n33093) );
  XNOR U5181 ( .A(n33094), .B(n32674), .Z(n32676) );
  XNOR U5182 ( .A(n32677), .B(n32251), .Z(n32253) );
  XNOR U5183 ( .A(n32254), .B(n31822), .Z(n31824) );
  XNOR U5184 ( .A(n31825), .B(n31387), .Z(n31389) );
  XNOR U5185 ( .A(n31390), .B(n30946), .Z(n30948) );
  XNOR U5186 ( .A(n30949), .B(n30499), .Z(n30501) );
  XNOR U5187 ( .A(n30502), .B(n30046), .Z(n30048) );
  XNOR U5188 ( .A(n30049), .B(n29587), .Z(n29589) );
  XNOR U5189 ( .A(n29590), .B(n29122), .Z(n29124) );
  XNOR U5190 ( .A(n29125), .B(n28651), .Z(n28653) );
  XNOR U5191 ( .A(n28654), .B(n28174), .Z(n28176) );
  XNOR U5192 ( .A(n28177), .B(n27691), .Z(n27693) );
  XNOR U5193 ( .A(n27694), .B(n27202), .Z(n27204) );
  XNOR U5194 ( .A(n27205), .B(n26705), .Z(n26707) );
  XNOR U5195 ( .A(n26708), .B(n26204), .Z(n26206) );
  XNOR U5196 ( .A(n26207), .B(n25696), .Z(n25698) );
  XNOR U5197 ( .A(n25699), .B(n25182), .Z(n25184) );
  XNOR U5198 ( .A(n25185), .B(n24659), .Z(n24661) );
  XNOR U5199 ( .A(n24662), .B(n24134), .Z(n24136) );
  XNOR U5200 ( .A(n24137), .B(n23603), .Z(n23605) );
  XNOR U5201 ( .A(n23606), .B(n23065), .Z(n23067) );
  XNOR U5202 ( .A(n23068), .B(n22521), .Z(n22523) );
  XNOR U5203 ( .A(n22524), .B(n21972), .Z(n21974) );
  XNOR U5204 ( .A(n21975), .B(n21417), .Z(n21419) );
  XNOR U5205 ( .A(n21420), .B(n20855), .Z(n20857) );
  XNOR U5206 ( .A(n20858), .B(n20288), .Z(n20290) );
  XNOR U5207 ( .A(n20291), .B(n19715), .Z(n19717) );
  XNOR U5208 ( .A(n19718), .B(n19136), .Z(n19138) );
  XOR U5209 ( .A(n18444), .B(n18641), .Z(n18448) );
  XOR U5210 ( .A(n17254), .B(n17419), .Z(n17258) );
  XOR U5211 ( .A(n16040), .B(n16205), .Z(n16044) );
  XOR U5212 ( .A(n14802), .B(n14967), .Z(n14806) );
  XOR U5213 ( .A(n13540), .B(n13705), .Z(n13544) );
  XOR U5214 ( .A(n12252), .B(n12419), .Z(n12256) );
  XOR U5215 ( .A(n9583), .B(n9778), .Z(n9587) );
  XOR U5216 ( .A(n5983), .B(n6370), .Z(n5987) );
  XOR U5217 ( .A(n7442), .B(n7751), .Z(n7446) );
  XOR U5218 ( .A(n7487), .B(n7742), .Z(n7491) );
  XNOR U5219 ( .A(n44499), .B(n44307), .Z(n44309) );
  XOR U5220 ( .A(n10268), .B(n10445), .Z(n10272) );
  XOR U5221 ( .A(n8857), .B(n9112), .Z(n8861) );
  XOR U5222 ( .A(n5290), .B(n5661), .Z(n5294) );
  XOR U5223 ( .A(n3840), .B(n4233), .Z(n3844) );
  XOR U5224 ( .A(n3795), .B(n4242), .Z(n3799) );
  XOR U5225 ( .A(n2321), .B(n2792), .Z(n2325) );
  XOR U5226 ( .A(n2276), .B(n2801), .Z(n2280) );
  XOR U5227 ( .A(n9613), .B(n9772), .Z(n9617) );
  XOR U5228 ( .A(n45353), .B(n45505), .Z(n45357) );
  XOR U5229 ( .A(n45029), .B(n45181), .Z(n45033) );
  XOR U5230 ( .A(n44681), .B(n44833), .Z(n44685) );
  XOR U5231 ( .A(n7517), .B(n7736), .Z(n7521) );
  XOR U5232 ( .A(n7472), .B(n7745), .Z(n7476) );
  XOR U5233 ( .A(n6013), .B(n6364), .Z(n6017) );
  XOR U5234 ( .A(n2306), .B(n2795), .Z(n2310) );
  XOR U5235 ( .A(n3825), .B(n4236), .Z(n3829) );
  XOR U5236 ( .A(n2351), .B(n2786), .Z(n2355) );
  XOR U5237 ( .A(n5320), .B(n5655), .Z(n5324) );
  XOR U5238 ( .A(n3870), .B(n4227), .Z(n3874) );
  XOR U5239 ( .A(n8887), .B(n9106), .Z(n8891) );
  XNOR U5240 ( .A(n44692), .B(n44506), .Z(n44508) );
  XNOR U5241 ( .A(n44509), .B(n44317), .Z(n44319) );
  XNOR U5242 ( .A(n44320), .B(n44122), .Z(n44124) );
  XNOR U5243 ( .A(n44125), .B(n43921), .Z(n43923) );
  XNOR U5244 ( .A(n43924), .B(n43714), .Z(n43716) );
  XNOR U5245 ( .A(n43717), .B(n43501), .Z(n43503) );
  XNOR U5246 ( .A(n43504), .B(n43282), .Z(n43284) );
  XNOR U5247 ( .A(n43285), .B(n43057), .Z(n43059) );
  XNOR U5248 ( .A(n43060), .B(n42826), .Z(n42828) );
  XNOR U5249 ( .A(n42829), .B(n42589), .Z(n42591) );
  XNOR U5250 ( .A(n42592), .B(n42346), .Z(n42348) );
  XNOR U5251 ( .A(n42349), .B(n42097), .Z(n42099) );
  XNOR U5252 ( .A(n42100), .B(n41842), .Z(n41844) );
  XNOR U5253 ( .A(n41845), .B(n41581), .Z(n41583) );
  XNOR U5254 ( .A(n41584), .B(n41314), .Z(n41316) );
  XNOR U5255 ( .A(n41317), .B(n41041), .Z(n41043) );
  XNOR U5256 ( .A(n41044), .B(n40762), .Z(n40764) );
  XNOR U5257 ( .A(n40765), .B(n40477), .Z(n40479) );
  XNOR U5258 ( .A(n40480), .B(n40186), .Z(n40188) );
  XNOR U5259 ( .A(n40189), .B(n39889), .Z(n39891) );
  XNOR U5260 ( .A(n39892), .B(n39586), .Z(n39588) );
  XNOR U5261 ( .A(n39589), .B(n39277), .Z(n39279) );
  XNOR U5262 ( .A(n39280), .B(n38962), .Z(n38964) );
  XNOR U5263 ( .A(n38965), .B(n38641), .Z(n38643) );
  XNOR U5264 ( .A(n38644), .B(n38314), .Z(n38316) );
  XNOR U5265 ( .A(n38317), .B(n37981), .Z(n37983) );
  XNOR U5266 ( .A(n37984), .B(n37642), .Z(n37644) );
  XNOR U5267 ( .A(n37645), .B(n37297), .Z(n37299) );
  XNOR U5268 ( .A(n37300), .B(n36946), .Z(n36948) );
  XNOR U5269 ( .A(n36949), .B(n36589), .Z(n36591) );
  XNOR U5270 ( .A(n36592), .B(n36226), .Z(n36228) );
  XNOR U5271 ( .A(n36229), .B(n35857), .Z(n35859) );
  XNOR U5272 ( .A(n35860), .B(n35482), .Z(n35484) );
  XNOR U5273 ( .A(n35485), .B(n35101), .Z(n35103) );
  XNOR U5274 ( .A(n35104), .B(n34714), .Z(n34716) );
  XNOR U5275 ( .A(n34717), .B(n34321), .Z(n34323) );
  XNOR U5276 ( .A(n34324), .B(n33922), .Z(n33924) );
  XNOR U5277 ( .A(n33925), .B(n33517), .Z(n33519) );
  XNOR U5278 ( .A(n33520), .B(n33106), .Z(n33108) );
  XNOR U5279 ( .A(n33109), .B(n32689), .Z(n32691) );
  XNOR U5280 ( .A(n32692), .B(n32266), .Z(n32268) );
  XNOR U5281 ( .A(n32269), .B(n31837), .Z(n31839) );
  XNOR U5282 ( .A(n31840), .B(n31402), .Z(n31404) );
  XNOR U5283 ( .A(n31405), .B(n30961), .Z(n30963) );
  XNOR U5284 ( .A(n30964), .B(n30514), .Z(n30516) );
  XNOR U5285 ( .A(n30517), .B(n30061), .Z(n30063) );
  XNOR U5286 ( .A(n30064), .B(n29602), .Z(n29604) );
  XNOR U5287 ( .A(n29605), .B(n29137), .Z(n29139) );
  XNOR U5288 ( .A(n29140), .B(n28666), .Z(n28668) );
  XNOR U5289 ( .A(n28669), .B(n28189), .Z(n28191) );
  XNOR U5290 ( .A(n28192), .B(n27706), .Z(n27708) );
  XNOR U5291 ( .A(n27709), .B(n27217), .Z(n27219) );
  XNOR U5292 ( .A(n27220), .B(n26720), .Z(n26722) );
  XNOR U5293 ( .A(n26723), .B(n26219), .Z(n26221) );
  XNOR U5294 ( .A(n26222), .B(n25711), .Z(n25713) );
  XNOR U5295 ( .A(n25714), .B(n25197), .Z(n25199) );
  XNOR U5296 ( .A(n25200), .B(n24674), .Z(n24676) );
  XNOR U5297 ( .A(n24677), .B(n24149), .Z(n24151) );
  XNOR U5298 ( .A(n24152), .B(n23618), .Z(n23620) );
  XNOR U5299 ( .A(n23621), .B(n23080), .Z(n23082) );
  XNOR U5300 ( .A(n23083), .B(n22536), .Z(n22538) );
  XNOR U5301 ( .A(n22539), .B(n21987), .Z(n21989) );
  XNOR U5302 ( .A(n21990), .B(n21432), .Z(n21434) );
  XNOR U5303 ( .A(n21435), .B(n20870), .Z(n20872) );
  XNOR U5304 ( .A(n20873), .B(n20303), .Z(n20305) );
  XNOR U5305 ( .A(n20306), .B(n19730), .Z(n19732) );
  XNOR U5306 ( .A(n19733), .B(n19151), .Z(n19153) );
  XOR U5307 ( .A(n18459), .B(n18635), .Z(n18463) );
  XOR U5308 ( .A(n17269), .B(n17416), .Z(n17273) );
  XOR U5309 ( .A(n16055), .B(n16202), .Z(n16059) );
  XOR U5310 ( .A(n14817), .B(n14964), .Z(n14821) );
  XOR U5311 ( .A(n13555), .B(n13702), .Z(n13559) );
  XOR U5312 ( .A(n12267), .B(n12416), .Z(n12271) );
  XOR U5313 ( .A(n6043), .B(n6358), .Z(n6047) );
  XOR U5314 ( .A(n7502), .B(n7739), .Z(n7506) );
  XOR U5315 ( .A(n7547), .B(n7730), .Z(n7551) );
  XNOR U5316 ( .A(n45045), .B(n44871), .Z(n44873) );
  XOR U5317 ( .A(n10298), .B(n10439), .Z(n10302) );
  XOR U5318 ( .A(n8917), .B(n9100), .Z(n8921) );
  XOR U5319 ( .A(n5350), .B(n5649), .Z(n5354) );
  XOR U5320 ( .A(n3900), .B(n4221), .Z(n3904) );
  XOR U5321 ( .A(n3855), .B(n4230), .Z(n3859) );
  XOR U5322 ( .A(n2381), .B(n2780), .Z(n2385) );
  XOR U5323 ( .A(n2336), .B(n2789), .Z(n2340) );
  XOR U5324 ( .A(n45809), .B(n45943), .Z(n45813) );
  XOR U5325 ( .A(n45521), .B(n45655), .Z(n45525) );
  XOR U5326 ( .A(n45209), .B(n45343), .Z(n45213) );
  XOR U5327 ( .A(n11625), .B(n11760), .Z(n11629) );
  XOR U5328 ( .A(n7577), .B(n7724), .Z(n7581) );
  XOR U5329 ( .A(n7532), .B(n7733), .Z(n7536) );
  XOR U5330 ( .A(n6073), .B(n6352), .Z(n6077) );
  XOR U5331 ( .A(n2366), .B(n2783), .Z(n2370) );
  XOR U5332 ( .A(n3885), .B(n4224), .Z(n3889) );
  XOR U5333 ( .A(n2411), .B(n2774), .Z(n2415) );
  XOR U5334 ( .A(n5380), .B(n5643), .Z(n5384) );
  XOR U5335 ( .A(n3930), .B(n4215), .Z(n3934) );
  XOR U5336 ( .A(n8947), .B(n9094), .Z(n8951) );
  XNOR U5337 ( .A(n45220), .B(n45052), .Z(n45054) );
  XNOR U5338 ( .A(n45055), .B(n44881), .Z(n44883) );
  XNOR U5339 ( .A(n44884), .B(n44704), .Z(n44706) );
  XNOR U5340 ( .A(n44707), .B(n44521), .Z(n44523) );
  XNOR U5341 ( .A(n44524), .B(n44332), .Z(n44334) );
  XNOR U5342 ( .A(n44335), .B(n44137), .Z(n44139) );
  XNOR U5343 ( .A(n44140), .B(n43936), .Z(n43938) );
  XNOR U5344 ( .A(n43939), .B(n43729), .Z(n43731) );
  XNOR U5345 ( .A(n43732), .B(n43516), .Z(n43518) );
  XNOR U5346 ( .A(n43519), .B(n43297), .Z(n43299) );
  XNOR U5347 ( .A(n43300), .B(n43072), .Z(n43074) );
  XNOR U5348 ( .A(n43075), .B(n42841), .Z(n42843) );
  XNOR U5349 ( .A(n42844), .B(n42604), .Z(n42606) );
  XNOR U5350 ( .A(n42607), .B(n42361), .Z(n42363) );
  XNOR U5351 ( .A(n42364), .B(n42112), .Z(n42114) );
  XNOR U5352 ( .A(n42115), .B(n41857), .Z(n41859) );
  XNOR U5353 ( .A(n41860), .B(n41596), .Z(n41598) );
  XNOR U5354 ( .A(n41599), .B(n41329), .Z(n41331) );
  XNOR U5355 ( .A(n41332), .B(n41056), .Z(n41058) );
  XNOR U5356 ( .A(n41059), .B(n40777), .Z(n40779) );
  XNOR U5357 ( .A(n40780), .B(n40492), .Z(n40494) );
  XNOR U5358 ( .A(n40495), .B(n40201), .Z(n40203) );
  XNOR U5359 ( .A(n40204), .B(n39904), .Z(n39906) );
  XNOR U5360 ( .A(n39907), .B(n39601), .Z(n39603) );
  XNOR U5361 ( .A(n39604), .B(n39292), .Z(n39294) );
  XNOR U5362 ( .A(n39295), .B(n38977), .Z(n38979) );
  XNOR U5363 ( .A(n38980), .B(n38656), .Z(n38658) );
  XNOR U5364 ( .A(n38659), .B(n38329), .Z(n38331) );
  XNOR U5365 ( .A(n38332), .B(n37996), .Z(n37998) );
  XNOR U5366 ( .A(n37999), .B(n37657), .Z(n37659) );
  XNOR U5367 ( .A(n37660), .B(n37312), .Z(n37314) );
  XNOR U5368 ( .A(n37315), .B(n36961), .Z(n36963) );
  XNOR U5369 ( .A(n36964), .B(n36604), .Z(n36606) );
  XNOR U5370 ( .A(n36607), .B(n36241), .Z(n36243) );
  XNOR U5371 ( .A(n36244), .B(n35872), .Z(n35874) );
  XNOR U5372 ( .A(n35875), .B(n35497), .Z(n35499) );
  XNOR U5373 ( .A(n35500), .B(n35116), .Z(n35118) );
  XNOR U5374 ( .A(n35119), .B(n34729), .Z(n34731) );
  XNOR U5375 ( .A(n34732), .B(n34336), .Z(n34338) );
  XNOR U5376 ( .A(n34339), .B(n33937), .Z(n33939) );
  XNOR U5377 ( .A(n33940), .B(n33532), .Z(n33534) );
  XNOR U5378 ( .A(n33535), .B(n33121), .Z(n33123) );
  XNOR U5379 ( .A(n33124), .B(n32704), .Z(n32706) );
  XNOR U5380 ( .A(n32707), .B(n32281), .Z(n32283) );
  XNOR U5381 ( .A(n32284), .B(n31852), .Z(n31854) );
  XNOR U5382 ( .A(n31855), .B(n31417), .Z(n31419) );
  XNOR U5383 ( .A(n31420), .B(n30976), .Z(n30978) );
  XNOR U5384 ( .A(n30979), .B(n30529), .Z(n30531) );
  XNOR U5385 ( .A(n30532), .B(n30076), .Z(n30078) );
  XNOR U5386 ( .A(n30079), .B(n29617), .Z(n29619) );
  XNOR U5387 ( .A(n29620), .B(n29152), .Z(n29154) );
  XNOR U5388 ( .A(n29155), .B(n28681), .Z(n28683) );
  XNOR U5389 ( .A(n28684), .B(n28204), .Z(n28206) );
  XNOR U5390 ( .A(n28207), .B(n27721), .Z(n27723) );
  XNOR U5391 ( .A(n27724), .B(n27232), .Z(n27234) );
  XNOR U5392 ( .A(n27235), .B(n26735), .Z(n26737) );
  XNOR U5393 ( .A(n26738), .B(n26234), .Z(n26236) );
  XNOR U5394 ( .A(n26237), .B(n25726), .Z(n25728) );
  XNOR U5395 ( .A(n25729), .B(n25212), .Z(n25214) );
  XNOR U5396 ( .A(n25215), .B(n24689), .Z(n24691) );
  XNOR U5397 ( .A(n24692), .B(n24164), .Z(n24166) );
  XNOR U5398 ( .A(n24167), .B(n23633), .Z(n23635) );
  XNOR U5399 ( .A(n23636), .B(n23095), .Z(n23097) );
  XNOR U5400 ( .A(n23098), .B(n22551), .Z(n22553) );
  XNOR U5401 ( .A(n22554), .B(n22002), .Z(n22004) );
  XNOR U5402 ( .A(n22005), .B(n21447), .Z(n21449) );
  XNOR U5403 ( .A(n21450), .B(n20885), .Z(n20887) );
  XNOR U5404 ( .A(n20888), .B(n20318), .Z(n20320) );
  XNOR U5405 ( .A(n20321), .B(n19745), .Z(n19747) );
  XNOR U5406 ( .A(n19748), .B(n19166), .Z(n19168) );
  XOR U5407 ( .A(n18474), .B(n18629), .Z(n18478) );
  XOR U5408 ( .A(n17284), .B(n17413), .Z(n17288) );
  XOR U5409 ( .A(n16070), .B(n16199), .Z(n16074) );
  XOR U5410 ( .A(n14832), .B(n14961), .Z(n14836) );
  XOR U5411 ( .A(n13570), .B(n13699), .Z(n13574) );
  XOR U5412 ( .A(n6103), .B(n6346), .Z(n6107) );
  XOR U5413 ( .A(n7562), .B(n7727), .Z(n7566) );
  XNOR U5414 ( .A(n45537), .B(n45381), .Z(n45383) );
  XOR U5415 ( .A(n10977), .B(n11100), .Z(n10981) );
  XOR U5416 ( .A(n5410), .B(n5637), .Z(n5414) );
  XOR U5417 ( .A(n3960), .B(n4209), .Z(n3964) );
  XOR U5418 ( .A(n3915), .B(n4218), .Z(n3919) );
  XOR U5419 ( .A(n2441), .B(n2768), .Z(n2445) );
  XOR U5420 ( .A(n2396), .B(n2777), .Z(n2400) );
  XOR U5421 ( .A(n46211), .B(n46327), .Z(n46215) );
  XOR U5422 ( .A(n45959), .B(n46075), .Z(n45963) );
  XOR U5423 ( .A(n45683), .B(n45799), .Z(n45687) );
  XOR U5424 ( .A(n12940), .B(n13057), .Z(n12944) );
  XOR U5425 ( .A(n10318), .B(n10435), .Z(n10322) );
  XOR U5426 ( .A(n6908), .B(n7025), .Z(n6912) );
  XOR U5427 ( .A(n7592), .B(n7721), .Z(n7596) );
  XOR U5428 ( .A(n6133), .B(n6340), .Z(n6137) );
  XOR U5429 ( .A(n2426), .B(n2771), .Z(n2430) );
  XOR U5430 ( .A(n3945), .B(n4212), .Z(n3949) );
  XOR U5431 ( .A(n2471), .B(n2762), .Z(n2475) );
  XOR U5432 ( .A(n5440), .B(n5631), .Z(n5444) );
  XOR U5433 ( .A(n3990), .B(n4203), .Z(n3994) );
  XNOR U5434 ( .A(n45694), .B(n45544), .Z(n45546) );
  XNOR U5435 ( .A(n45547), .B(n45391), .Z(n45393) );
  XNOR U5436 ( .A(n45394), .B(n45232), .Z(n45234) );
  XNOR U5437 ( .A(n45235), .B(n45067), .Z(n45069) );
  XNOR U5438 ( .A(n45070), .B(n44896), .Z(n44898) );
  XNOR U5439 ( .A(n44899), .B(n44719), .Z(n44721) );
  XNOR U5440 ( .A(n44722), .B(n44536), .Z(n44538) );
  XNOR U5441 ( .A(n44539), .B(n44347), .Z(n44349) );
  XNOR U5442 ( .A(n44350), .B(n44152), .Z(n44154) );
  XNOR U5443 ( .A(n44155), .B(n43951), .Z(n43953) );
  XNOR U5444 ( .A(n43954), .B(n43744), .Z(n43746) );
  XNOR U5445 ( .A(n43747), .B(n43531), .Z(n43533) );
  XNOR U5446 ( .A(n43534), .B(n43312), .Z(n43314) );
  XNOR U5447 ( .A(n43315), .B(n43087), .Z(n43089) );
  XNOR U5448 ( .A(n43090), .B(n42856), .Z(n42858) );
  XNOR U5449 ( .A(n42859), .B(n42619), .Z(n42621) );
  XNOR U5450 ( .A(n42622), .B(n42376), .Z(n42378) );
  XNOR U5451 ( .A(n42379), .B(n42127), .Z(n42129) );
  XNOR U5452 ( .A(n42130), .B(n41872), .Z(n41874) );
  XNOR U5453 ( .A(n41875), .B(n41611), .Z(n41613) );
  XNOR U5454 ( .A(n41614), .B(n41344), .Z(n41346) );
  XNOR U5455 ( .A(n41347), .B(n41071), .Z(n41073) );
  XNOR U5456 ( .A(n41074), .B(n40792), .Z(n40794) );
  XNOR U5457 ( .A(n40795), .B(n40507), .Z(n40509) );
  XNOR U5458 ( .A(n40510), .B(n40216), .Z(n40218) );
  XNOR U5459 ( .A(n40219), .B(n39919), .Z(n39921) );
  XNOR U5460 ( .A(n39922), .B(n39616), .Z(n39618) );
  XNOR U5461 ( .A(n39619), .B(n39307), .Z(n39309) );
  XNOR U5462 ( .A(n39310), .B(n38992), .Z(n38994) );
  XNOR U5463 ( .A(n38995), .B(n38671), .Z(n38673) );
  XNOR U5464 ( .A(n38674), .B(n38344), .Z(n38346) );
  XNOR U5465 ( .A(n38347), .B(n38011), .Z(n38013) );
  XNOR U5466 ( .A(n38014), .B(n37672), .Z(n37674) );
  XNOR U5467 ( .A(n37675), .B(n37327), .Z(n37329) );
  XNOR U5468 ( .A(n37330), .B(n36976), .Z(n36978) );
  XNOR U5469 ( .A(n36979), .B(n36619), .Z(n36621) );
  XNOR U5470 ( .A(n36622), .B(n36256), .Z(n36258) );
  XNOR U5471 ( .A(n36259), .B(n35887), .Z(n35889) );
  XNOR U5472 ( .A(n35890), .B(n35512), .Z(n35514) );
  XNOR U5473 ( .A(n35515), .B(n35131), .Z(n35133) );
  XNOR U5474 ( .A(n35134), .B(n34744), .Z(n34746) );
  XNOR U5475 ( .A(n34747), .B(n34351), .Z(n34353) );
  XNOR U5476 ( .A(n34354), .B(n33952), .Z(n33954) );
  XNOR U5477 ( .A(n33955), .B(n33547), .Z(n33549) );
  XNOR U5478 ( .A(n33550), .B(n33136), .Z(n33138) );
  XNOR U5479 ( .A(n33139), .B(n32719), .Z(n32721) );
  XNOR U5480 ( .A(n32722), .B(n32296), .Z(n32298) );
  XNOR U5481 ( .A(n32299), .B(n31867), .Z(n31869) );
  XNOR U5482 ( .A(n31870), .B(n31432), .Z(n31434) );
  XNOR U5483 ( .A(n31435), .B(n30991), .Z(n30993) );
  XNOR U5484 ( .A(n30994), .B(n30544), .Z(n30546) );
  XNOR U5485 ( .A(n30547), .B(n30091), .Z(n30093) );
  XNOR U5486 ( .A(n30094), .B(n29632), .Z(n29634) );
  XNOR U5487 ( .A(n29635), .B(n29167), .Z(n29169) );
  XNOR U5488 ( .A(n29170), .B(n28696), .Z(n28698) );
  XNOR U5489 ( .A(n28699), .B(n28219), .Z(n28221) );
  XNOR U5490 ( .A(n28222), .B(n27736), .Z(n27738) );
  XNOR U5491 ( .A(n27739), .B(n27247), .Z(n27249) );
  XNOR U5492 ( .A(n27250), .B(n26750), .Z(n26752) );
  XNOR U5493 ( .A(n26753), .B(n26249), .Z(n26251) );
  XNOR U5494 ( .A(n26252), .B(n25741), .Z(n25743) );
  XNOR U5495 ( .A(n25744), .B(n25227), .Z(n25229) );
  XNOR U5496 ( .A(n25230), .B(n24704), .Z(n24706) );
  XNOR U5497 ( .A(n24707), .B(n24179), .Z(n24181) );
  XNOR U5498 ( .A(n24182), .B(n23648), .Z(n23650) );
  XNOR U5499 ( .A(n23651), .B(n23110), .Z(n23112) );
  XNOR U5500 ( .A(n23113), .B(n22566), .Z(n22568) );
  XNOR U5501 ( .A(n22569), .B(n22017), .Z(n22019) );
  XNOR U5502 ( .A(n22020), .B(n21462), .Z(n21464) );
  XNOR U5503 ( .A(n21465), .B(n20900), .Z(n20902) );
  XNOR U5504 ( .A(n20903), .B(n20333), .Z(n20335) );
  XNOR U5505 ( .A(n20336), .B(n19760), .Z(n19762) );
  XNOR U5506 ( .A(n19763), .B(n19181), .Z(n19183) );
  XOR U5507 ( .A(n17897), .B(n18008), .Z(n17901) );
  XOR U5508 ( .A(n16695), .B(n16806), .Z(n16699) );
  XOR U5509 ( .A(n15469), .B(n15580), .Z(n15473) );
  XOR U5510 ( .A(n14219), .B(n14330), .Z(n14223) );
  XOR U5511 ( .A(n9653), .B(n9764), .Z(n9657) );
  XOR U5512 ( .A(n8295), .B(n8406), .Z(n8299) );
  XOR U5513 ( .A(n6163), .B(n6334), .Z(n6167) );
  XNOR U5514 ( .A(n45975), .B(n45837), .Z(n45839) );
  XOR U5515 ( .A(n12302), .B(n12409), .Z(n12306) );
  XOR U5516 ( .A(n5470), .B(n5625), .Z(n5474) );
  XOR U5517 ( .A(n4020), .B(n4197), .Z(n4024) );
  XOR U5518 ( .A(n3975), .B(n4206), .Z(n3979) );
  XOR U5519 ( .A(n2501), .B(n2756), .Z(n2505) );
  XOR U5520 ( .A(n2456), .B(n2765), .Z(n2460) );
  XOR U5521 ( .A(n46559), .B(n46657), .Z(n46563) );
  XOR U5522 ( .A(n46343), .B(n46441), .Z(n46347) );
  XOR U5523 ( .A(n46103), .B(n46201), .Z(n46107) );
  XOR U5524 ( .A(n11655), .B(n11754), .Z(n11659) );
  XOR U5525 ( .A(n6193), .B(n6328), .Z(n6197) );
  XOR U5526 ( .A(n2486), .B(n2759), .Z(n2490) );
  XOR U5527 ( .A(n4005), .B(n4200), .Z(n4009) );
  XOR U5528 ( .A(n2531), .B(n2750), .Z(n2535) );
  XOR U5529 ( .A(n5500), .B(n5619), .Z(n5504) );
  XOR U5530 ( .A(n4050), .B(n4191), .Z(n4054) );
  XNOR U5531 ( .A(n46114), .B(n45982), .Z(n45984) );
  XNOR U5532 ( .A(n45985), .B(n45847), .Z(n45849) );
  XNOR U5533 ( .A(n45850), .B(n45706), .Z(n45708) );
  XNOR U5534 ( .A(n45709), .B(n45559), .Z(n45561) );
  XNOR U5535 ( .A(n45562), .B(n45406), .Z(n45408) );
  XNOR U5536 ( .A(n45409), .B(n45247), .Z(n45249) );
  XNOR U5537 ( .A(n45250), .B(n45082), .Z(n45084) );
  XNOR U5538 ( .A(n45085), .B(n44911), .Z(n44913) );
  XNOR U5539 ( .A(n44914), .B(n44734), .Z(n44736) );
  XNOR U5540 ( .A(n44737), .B(n44551), .Z(n44553) );
  XNOR U5541 ( .A(n44554), .B(n44362), .Z(n44364) );
  XNOR U5542 ( .A(n44365), .B(n44167), .Z(n44169) );
  XNOR U5543 ( .A(n44170), .B(n43966), .Z(n43968) );
  XNOR U5544 ( .A(n43969), .B(n43759), .Z(n43761) );
  XNOR U5545 ( .A(n43762), .B(n43546), .Z(n43548) );
  XNOR U5546 ( .A(n43549), .B(n43327), .Z(n43329) );
  XNOR U5547 ( .A(n43330), .B(n43102), .Z(n43104) );
  XNOR U5548 ( .A(n43105), .B(n42871), .Z(n42873) );
  XNOR U5549 ( .A(n42874), .B(n42634), .Z(n42636) );
  XNOR U5550 ( .A(n42637), .B(n42391), .Z(n42393) );
  XNOR U5551 ( .A(n42394), .B(n42142), .Z(n42144) );
  XNOR U5552 ( .A(n42145), .B(n41887), .Z(n41889) );
  XNOR U5553 ( .A(n41890), .B(n41626), .Z(n41628) );
  XNOR U5554 ( .A(n41629), .B(n41359), .Z(n41361) );
  XNOR U5555 ( .A(n41362), .B(n41086), .Z(n41088) );
  XNOR U5556 ( .A(n41089), .B(n40807), .Z(n40809) );
  XNOR U5557 ( .A(n40810), .B(n40522), .Z(n40524) );
  XNOR U5558 ( .A(n40525), .B(n40231), .Z(n40233) );
  XNOR U5559 ( .A(n40234), .B(n39934), .Z(n39936) );
  XNOR U5560 ( .A(n39937), .B(n39631), .Z(n39633) );
  XNOR U5561 ( .A(n39634), .B(n39322), .Z(n39324) );
  XNOR U5562 ( .A(n39325), .B(n39007), .Z(n39009) );
  XNOR U5563 ( .A(n39010), .B(n38686), .Z(n38688) );
  XNOR U5564 ( .A(n38689), .B(n38359), .Z(n38361) );
  XNOR U5565 ( .A(n38362), .B(n38026), .Z(n38028) );
  XNOR U5566 ( .A(n38029), .B(n37687), .Z(n37689) );
  XNOR U5567 ( .A(n37690), .B(n37342), .Z(n37344) );
  XNOR U5568 ( .A(n37345), .B(n36991), .Z(n36993) );
  XNOR U5569 ( .A(n36994), .B(n36634), .Z(n36636) );
  XNOR U5570 ( .A(n36637), .B(n36271), .Z(n36273) );
  XNOR U5571 ( .A(n36274), .B(n35902), .Z(n35904) );
  XNOR U5572 ( .A(n35905), .B(n35527), .Z(n35529) );
  XNOR U5573 ( .A(n35530), .B(n35146), .Z(n35148) );
  XNOR U5574 ( .A(n35149), .B(n34759), .Z(n34761) );
  XNOR U5575 ( .A(n34762), .B(n34366), .Z(n34368) );
  XNOR U5576 ( .A(n34369), .B(n33967), .Z(n33969) );
  XNOR U5577 ( .A(n33970), .B(n33562), .Z(n33564) );
  XNOR U5578 ( .A(n33565), .B(n33151), .Z(n33153) );
  XNOR U5579 ( .A(n33154), .B(n32734), .Z(n32736) );
  XNOR U5580 ( .A(n32737), .B(n32311), .Z(n32313) );
  XNOR U5581 ( .A(n32314), .B(n31882), .Z(n31884) );
  XNOR U5582 ( .A(n31885), .B(n31447), .Z(n31449) );
  XNOR U5583 ( .A(n31450), .B(n31006), .Z(n31008) );
  XNOR U5584 ( .A(n31009), .B(n30559), .Z(n30561) );
  XNOR U5585 ( .A(n30562), .B(n30106), .Z(n30108) );
  XNOR U5586 ( .A(n30109), .B(n29647), .Z(n29649) );
  XNOR U5587 ( .A(n29650), .B(n29182), .Z(n29184) );
  XNOR U5588 ( .A(n29185), .B(n28711), .Z(n28713) );
  XNOR U5589 ( .A(n28714), .B(n28234), .Z(n28236) );
  XNOR U5590 ( .A(n28237), .B(n27751), .Z(n27753) );
  XNOR U5591 ( .A(n27754), .B(n27262), .Z(n27264) );
  XNOR U5592 ( .A(n27265), .B(n26765), .Z(n26767) );
  XNOR U5593 ( .A(n26768), .B(n26264), .Z(n26266) );
  XNOR U5594 ( .A(n26267), .B(n25756), .Z(n25758) );
  XNOR U5595 ( .A(n25759), .B(n25242), .Z(n25244) );
  XNOR U5596 ( .A(n25245), .B(n24719), .Z(n24721) );
  XNOR U5597 ( .A(n24722), .B(n24194), .Z(n24196) );
  XNOR U5598 ( .A(n24197), .B(n23663), .Z(n23665) );
  XNOR U5599 ( .A(n23666), .B(n23125), .Z(n23127) );
  XNOR U5600 ( .A(n23128), .B(n22581), .Z(n22583) );
  XNOR U5601 ( .A(n22584), .B(n22032), .Z(n22034) );
  XNOR U5602 ( .A(n22035), .B(n21477), .Z(n21479) );
  XNOR U5603 ( .A(n21480), .B(n20915), .Z(n20917) );
  XNOR U5604 ( .A(n20918), .B(n20348), .Z(n20350) );
  XNOR U5605 ( .A(n20351), .B(n19775), .Z(n19777) );
  XNOR U5606 ( .A(n19778), .B(n19196), .Z(n19198) );
  XOR U5607 ( .A(n18504), .B(n18617), .Z(n18508) );
  XOR U5608 ( .A(n17314), .B(n17407), .Z(n17318) );
  XOR U5609 ( .A(n16100), .B(n16193), .Z(n16104) );
  XOR U5610 ( .A(n14862), .B(n14955), .Z(n14866) );
  XOR U5611 ( .A(n11002), .B(n11095), .Z(n11006) );
  XOR U5612 ( .A(n9668), .B(n9761), .Z(n9672) );
  XOR U5613 ( .A(n8310), .B(n8403), .Z(n8314) );
  XOR U5614 ( .A(n6223), .B(n6322), .Z(n6227) );
  XNOR U5615 ( .A(n46359), .B(n46239), .Z(n46241) );
  XOR U5616 ( .A(n13605), .B(n13692), .Z(n13609) );
  XOR U5617 ( .A(n4080), .B(n4185), .Z(n4084) );
  XOR U5618 ( .A(n4035), .B(n4194), .Z(n4039) );
  XOR U5619 ( .A(n2561), .B(n2744), .Z(n2565) );
  XOR U5620 ( .A(n2516), .B(n2753), .Z(n2520) );
  XOR U5621 ( .A(n46853), .B(n46933), .Z(n46857) );
  XOR U5622 ( .A(n46673), .B(n46753), .Z(n46677) );
  XOR U5623 ( .A(n46469), .B(n46549), .Z(n46473) );
  XOR U5624 ( .A(n2546), .B(n2747), .Z(n2550) );
  XOR U5625 ( .A(n4065), .B(n4188), .Z(n4069) );
  XOR U5626 ( .A(n2591), .B(n2738), .Z(n2595) );
  XNOR U5627 ( .A(n46480), .B(n46366), .Z(n46368) );
  XNOR U5628 ( .A(n46369), .B(n46249), .Z(n46251) );
  XNOR U5629 ( .A(n46252), .B(n46126), .Z(n46128) );
  XNOR U5630 ( .A(n46129), .B(n45997), .Z(n45999) );
  XNOR U5631 ( .A(n46000), .B(n45862), .Z(n45864) );
  XNOR U5632 ( .A(n45865), .B(n45721), .Z(n45723) );
  XNOR U5633 ( .A(n45724), .B(n45574), .Z(n45576) );
  XNOR U5634 ( .A(n45577), .B(n45421), .Z(n45423) );
  XNOR U5635 ( .A(n45424), .B(n45262), .Z(n45264) );
  XNOR U5636 ( .A(n45265), .B(n45097), .Z(n45099) );
  XNOR U5637 ( .A(n45100), .B(n44926), .Z(n44928) );
  XNOR U5638 ( .A(n44929), .B(n44749), .Z(n44751) );
  XNOR U5639 ( .A(n44752), .B(n44566), .Z(n44568) );
  XNOR U5640 ( .A(n44569), .B(n44377), .Z(n44379) );
  XNOR U5641 ( .A(n44380), .B(n44182), .Z(n44184) );
  XNOR U5642 ( .A(n44185), .B(n43981), .Z(n43983) );
  XNOR U5643 ( .A(n43984), .B(n43774), .Z(n43776) );
  XNOR U5644 ( .A(n43777), .B(n43561), .Z(n43563) );
  XNOR U5645 ( .A(n43564), .B(n43342), .Z(n43344) );
  XNOR U5646 ( .A(n43345), .B(n43117), .Z(n43119) );
  XNOR U5647 ( .A(n43120), .B(n42886), .Z(n42888) );
  XNOR U5648 ( .A(n42889), .B(n42649), .Z(n42651) );
  XNOR U5649 ( .A(n42652), .B(n42406), .Z(n42408) );
  XNOR U5650 ( .A(n42409), .B(n42157), .Z(n42159) );
  XNOR U5651 ( .A(n42160), .B(n41902), .Z(n41904) );
  XNOR U5652 ( .A(n41905), .B(n41641), .Z(n41643) );
  XNOR U5653 ( .A(n41644), .B(n41374), .Z(n41376) );
  XNOR U5654 ( .A(n41377), .B(n41101), .Z(n41103) );
  XNOR U5655 ( .A(n41104), .B(n40822), .Z(n40824) );
  XNOR U5656 ( .A(n40825), .B(n40537), .Z(n40539) );
  XNOR U5657 ( .A(n40540), .B(n40246), .Z(n40248) );
  XNOR U5658 ( .A(n40249), .B(n39949), .Z(n39951) );
  XNOR U5659 ( .A(n39952), .B(n39646), .Z(n39648) );
  XNOR U5660 ( .A(n39649), .B(n39337), .Z(n39339) );
  XNOR U5661 ( .A(n39340), .B(n39022), .Z(n39024) );
  XNOR U5662 ( .A(n39025), .B(n38701), .Z(n38703) );
  XNOR U5663 ( .A(n38704), .B(n38374), .Z(n38376) );
  XNOR U5664 ( .A(n38377), .B(n38041), .Z(n38043) );
  XNOR U5665 ( .A(n38044), .B(n37702), .Z(n37704) );
  XNOR U5666 ( .A(n37705), .B(n37357), .Z(n37359) );
  XNOR U5667 ( .A(n37360), .B(n37006), .Z(n37008) );
  XNOR U5668 ( .A(n37009), .B(n36649), .Z(n36651) );
  XNOR U5669 ( .A(n36652), .B(n36286), .Z(n36288) );
  XNOR U5670 ( .A(n36289), .B(n35917), .Z(n35919) );
  XNOR U5671 ( .A(n35920), .B(n35542), .Z(n35544) );
  XNOR U5672 ( .A(n35545), .B(n35161), .Z(n35163) );
  XNOR U5673 ( .A(n35164), .B(n34774), .Z(n34776) );
  XNOR U5674 ( .A(n34777), .B(n34381), .Z(n34383) );
  XNOR U5675 ( .A(n34384), .B(n33982), .Z(n33984) );
  XNOR U5676 ( .A(n33985), .B(n33577), .Z(n33579) );
  XNOR U5677 ( .A(n33580), .B(n33166), .Z(n33168) );
  XNOR U5678 ( .A(n33169), .B(n32749), .Z(n32751) );
  XNOR U5679 ( .A(n32752), .B(n32326), .Z(n32328) );
  XNOR U5680 ( .A(n32329), .B(n31897), .Z(n31899) );
  XNOR U5681 ( .A(n31900), .B(n31462), .Z(n31464) );
  XNOR U5682 ( .A(n31465), .B(n31021), .Z(n31023) );
  XNOR U5683 ( .A(n31024), .B(n30574), .Z(n30576) );
  XNOR U5684 ( .A(n30577), .B(n30121), .Z(n30123) );
  XNOR U5685 ( .A(n30124), .B(n29662), .Z(n29664) );
  XNOR U5686 ( .A(n29665), .B(n29197), .Z(n29199) );
  XNOR U5687 ( .A(n29200), .B(n28726), .Z(n28728) );
  XNOR U5688 ( .A(n28729), .B(n28249), .Z(n28251) );
  XNOR U5689 ( .A(n28252), .B(n27766), .Z(n27768) );
  XNOR U5690 ( .A(n27769), .B(n27277), .Z(n27279) );
  XNOR U5691 ( .A(n27280), .B(n26780), .Z(n26782) );
  XNOR U5692 ( .A(n26783), .B(n26279), .Z(n26281) );
  XNOR U5693 ( .A(n26282), .B(n25771), .Z(n25773) );
  XNOR U5694 ( .A(n25774), .B(n25257), .Z(n25259) );
  XNOR U5695 ( .A(n25260), .B(n24734), .Z(n24736) );
  XNOR U5696 ( .A(n24737), .B(n24209), .Z(n24211) );
  XNOR U5697 ( .A(n24212), .B(n23678), .Z(n23680) );
  XNOR U5698 ( .A(n23681), .B(n23140), .Z(n23142) );
  XNOR U5699 ( .A(n23143), .B(n22596), .Z(n22598) );
  XNOR U5700 ( .A(n22599), .B(n22047), .Z(n22049) );
  XNOR U5701 ( .A(n22050), .B(n21492), .Z(n21494) );
  XNOR U5702 ( .A(n21495), .B(n20930), .Z(n20932) );
  XNOR U5703 ( .A(n20933), .B(n20363), .Z(n20365) );
  XNOR U5704 ( .A(n20366), .B(n19790), .Z(n19792) );
  XNOR U5705 ( .A(n19793), .B(n19211), .Z(n19213) );
  XOR U5706 ( .A(n17927), .B(n18002), .Z(n17931) );
  XOR U5707 ( .A(n16725), .B(n16800), .Z(n16729) );
  XOR U5708 ( .A(n15499), .B(n15574), .Z(n15503) );
  XOR U5709 ( .A(n12975), .B(n13050), .Z(n12979) );
  XOR U5710 ( .A(n11675), .B(n11750), .Z(n11679) );
  XOR U5711 ( .A(n10353), .B(n10428), .Z(n10357) );
  XOR U5712 ( .A(n9007), .B(n9082), .Z(n9011) );
  XOR U5713 ( .A(n7637), .B(n7712), .Z(n7641) );
  XOR U5714 ( .A(n6243), .B(n6318), .Z(n6247) );
  XOR U5715 ( .A(n3381), .B(n3456), .Z(n3385) );
  XNOR U5716 ( .A(n46689), .B(n46587), .Z(n46589) );
  XOR U5717 ( .A(n14882), .B(n14951), .Z(n14886) );
  XOR U5718 ( .A(n4095), .B(n4182), .Z(n4099) );
  XOR U5719 ( .A(n2621), .B(n2732), .Z(n2625) );
  XOR U5720 ( .A(n2576), .B(n2741), .Z(n2580) );
  XOR U5721 ( .A(n47093), .B(n47155), .Z(n47097) );
  XOR U5722 ( .A(n46949), .B(n47011), .Z(n46953) );
  XOR U5723 ( .A(n46781), .B(n46843), .Z(n46785) );
  XOR U5724 ( .A(n1925), .B(n1988), .Z(n1929) );
  XOR U5725 ( .A(n2606), .B(n2735), .Z(n2610) );
  XNOR U5726 ( .A(n46792), .B(n46696), .Z(n46698) );
  XNOR U5727 ( .A(n46699), .B(n46597), .Z(n46599) );
  XNOR U5728 ( .A(n46600), .B(n46492), .Z(n46494) );
  XNOR U5729 ( .A(n46495), .B(n46381), .Z(n46383) );
  XNOR U5730 ( .A(n46384), .B(n46264), .Z(n46266) );
  XNOR U5731 ( .A(n46267), .B(n46141), .Z(n46143) );
  XNOR U5732 ( .A(n46144), .B(n46012), .Z(n46014) );
  XNOR U5733 ( .A(n46015), .B(n45877), .Z(n45879) );
  XNOR U5734 ( .A(n45880), .B(n45736), .Z(n45738) );
  XNOR U5735 ( .A(n45739), .B(n45589), .Z(n45591) );
  XNOR U5736 ( .A(n45592), .B(n45436), .Z(n45438) );
  XNOR U5737 ( .A(n45439), .B(n45277), .Z(n45279) );
  XNOR U5738 ( .A(n45280), .B(n45112), .Z(n45114) );
  XNOR U5739 ( .A(n45115), .B(n44941), .Z(n44943) );
  XNOR U5740 ( .A(n44944), .B(n44764), .Z(n44766) );
  XNOR U5741 ( .A(n44767), .B(n44581), .Z(n44583) );
  XNOR U5742 ( .A(n44584), .B(n44392), .Z(n44394) );
  XNOR U5743 ( .A(n44395), .B(n44197), .Z(n44199) );
  XNOR U5744 ( .A(n44200), .B(n43996), .Z(n43998) );
  XNOR U5745 ( .A(n43999), .B(n43789), .Z(n43791) );
  XNOR U5746 ( .A(n43792), .B(n43576), .Z(n43578) );
  XNOR U5747 ( .A(n43579), .B(n43357), .Z(n43359) );
  XNOR U5748 ( .A(n43360), .B(n43132), .Z(n43134) );
  XNOR U5749 ( .A(n43135), .B(n42901), .Z(n42903) );
  XNOR U5750 ( .A(n42904), .B(n42664), .Z(n42666) );
  XNOR U5751 ( .A(n42667), .B(n42421), .Z(n42423) );
  XNOR U5752 ( .A(n42424), .B(n42172), .Z(n42174) );
  XNOR U5753 ( .A(n42175), .B(n41917), .Z(n41919) );
  XNOR U5754 ( .A(n41920), .B(n41656), .Z(n41658) );
  XNOR U5755 ( .A(n41659), .B(n41389), .Z(n41391) );
  XNOR U5756 ( .A(n41392), .B(n41116), .Z(n41118) );
  XNOR U5757 ( .A(n41119), .B(n40837), .Z(n40839) );
  XNOR U5758 ( .A(n40840), .B(n40552), .Z(n40554) );
  XNOR U5759 ( .A(n40555), .B(n40261), .Z(n40263) );
  XNOR U5760 ( .A(n40264), .B(n39964), .Z(n39966) );
  XNOR U5761 ( .A(n39967), .B(n39661), .Z(n39663) );
  XNOR U5762 ( .A(n39664), .B(n39352), .Z(n39354) );
  XNOR U5763 ( .A(n39355), .B(n39037), .Z(n39039) );
  XNOR U5764 ( .A(n39040), .B(n38716), .Z(n38718) );
  XNOR U5765 ( .A(n38719), .B(n38389), .Z(n38391) );
  XNOR U5766 ( .A(n38392), .B(n38056), .Z(n38058) );
  XNOR U5767 ( .A(n38059), .B(n37717), .Z(n37719) );
  XNOR U5768 ( .A(n37720), .B(n37372), .Z(n37374) );
  XNOR U5769 ( .A(n37375), .B(n37021), .Z(n37023) );
  XNOR U5770 ( .A(n37024), .B(n36664), .Z(n36666) );
  XNOR U5771 ( .A(n36667), .B(n36301), .Z(n36303) );
  XNOR U5772 ( .A(n36304), .B(n35932), .Z(n35934) );
  XNOR U5773 ( .A(n35935), .B(n35557), .Z(n35559) );
  XNOR U5774 ( .A(n35560), .B(n35176), .Z(n35178) );
  XNOR U5775 ( .A(n35179), .B(n34789), .Z(n34791) );
  XNOR U5776 ( .A(n34792), .B(n34396), .Z(n34398) );
  XNOR U5777 ( .A(n34399), .B(n33997), .Z(n33999) );
  XNOR U5778 ( .A(n34000), .B(n33592), .Z(n33594) );
  XNOR U5779 ( .A(n33595), .B(n33181), .Z(n33183) );
  XNOR U5780 ( .A(n33184), .B(n32764), .Z(n32766) );
  XNOR U5781 ( .A(n32767), .B(n32341), .Z(n32343) );
  XNOR U5782 ( .A(n32344), .B(n31912), .Z(n31914) );
  XNOR U5783 ( .A(n31915), .B(n31477), .Z(n31479) );
  XNOR U5784 ( .A(n31480), .B(n31036), .Z(n31038) );
  XNOR U5785 ( .A(n31039), .B(n30589), .Z(n30591) );
  XNOR U5786 ( .A(n30592), .B(n30136), .Z(n30138) );
  XNOR U5787 ( .A(n30139), .B(n29677), .Z(n29679) );
  XNOR U5788 ( .A(n29680), .B(n29212), .Z(n29214) );
  XNOR U5789 ( .A(n29215), .B(n28741), .Z(n28743) );
  XNOR U5790 ( .A(n28744), .B(n28264), .Z(n28266) );
  XNOR U5791 ( .A(n28267), .B(n27781), .Z(n27783) );
  XNOR U5792 ( .A(n27784), .B(n27292), .Z(n27294) );
  XNOR U5793 ( .A(n27295), .B(n26795), .Z(n26797) );
  XNOR U5794 ( .A(n26798), .B(n26294), .Z(n26296) );
  XNOR U5795 ( .A(n26297), .B(n25786), .Z(n25788) );
  XNOR U5796 ( .A(n25789), .B(n25272), .Z(n25274) );
  XNOR U5797 ( .A(n25275), .B(n24749), .Z(n24751) );
  XNOR U5798 ( .A(n24752), .B(n24224), .Z(n24226) );
  XNOR U5799 ( .A(n24227), .B(n23693), .Z(n23695) );
  XNOR U5800 ( .A(n23696), .B(n23155), .Z(n23157) );
  XNOR U5801 ( .A(n23158), .B(n22611), .Z(n22613) );
  XNOR U5802 ( .A(n22614), .B(n22062), .Z(n22064) );
  XNOR U5803 ( .A(n22065), .B(n21507), .Z(n21509) );
  XNOR U5804 ( .A(n21510), .B(n20945), .Z(n20947) );
  XNOR U5805 ( .A(n20948), .B(n20378), .Z(n20380) );
  XNOR U5806 ( .A(n20381), .B(n19805), .Z(n19807) );
  XNOR U5807 ( .A(n19808), .B(n19226), .Z(n19228) );
  XOR U5808 ( .A(n18534), .B(n18605), .Z(n18538) );
  XOR U5809 ( .A(n17344), .B(n17401), .Z(n17348) );
  XOR U5810 ( .A(n14264), .B(n14321), .Z(n14268) );
  XOR U5811 ( .A(n12990), .B(n13047), .Z(n12994) );
  XOR U5812 ( .A(n11690), .B(n11747), .Z(n11694) );
  XOR U5813 ( .A(n10368), .B(n10425), .Z(n10372) );
  XOR U5814 ( .A(n9022), .B(n9079), .Z(n9026) );
  XOR U5815 ( .A(n7652), .B(n7709), .Z(n7656) );
  XOR U5816 ( .A(n6258), .B(n6315), .Z(n6262) );
  XOR U5817 ( .A(n4838), .B(n4895), .Z(n4842) );
  XOR U5818 ( .A(n2656), .B(n2725), .Z(n2660) );
  XNOR U5819 ( .A(n46965), .B(n46881), .Z(n46883) );
  XOR U5820 ( .A(n16745), .B(n16796), .Z(n16749) );
  XOR U5821 ( .A(n2636), .B(n2729), .Z(n2640) );
  XOR U5822 ( .A(n47171), .B(n47214), .Z(n47175) );
  XOR U5823 ( .A(n47039), .B(n47083), .Z(n47043) );
  XNOR U5824 ( .A(n47373), .B(n47331), .Z(n47333) );
  XNOR U5825 ( .A(n47334), .B(n47286), .Z(n47288) );
  XNOR U5826 ( .A(n47050), .B(n46972), .Z(n46974) );
  XNOR U5827 ( .A(n46975), .B(n46891), .Z(n46893) );
  XNOR U5828 ( .A(n46894), .B(n46804), .Z(n46806) );
  XNOR U5829 ( .A(n46807), .B(n46711), .Z(n46713) );
  XNOR U5830 ( .A(n46714), .B(n46612), .Z(n46614) );
  XNOR U5831 ( .A(n46615), .B(n46507), .Z(n46509) );
  XNOR U5832 ( .A(n46510), .B(n46396), .Z(n46398) );
  XNOR U5833 ( .A(n46399), .B(n46279), .Z(n46281) );
  XNOR U5834 ( .A(n46282), .B(n46156), .Z(n46158) );
  XNOR U5835 ( .A(n46159), .B(n46027), .Z(n46029) );
  XNOR U5836 ( .A(n46030), .B(n45892), .Z(n45894) );
  XNOR U5837 ( .A(n45895), .B(n45751), .Z(n45753) );
  XNOR U5838 ( .A(n45754), .B(n45604), .Z(n45606) );
  XNOR U5839 ( .A(n45607), .B(n45451), .Z(n45453) );
  XNOR U5840 ( .A(n45454), .B(n45292), .Z(n45294) );
  XNOR U5841 ( .A(n45295), .B(n45127), .Z(n45129) );
  XNOR U5842 ( .A(n45130), .B(n44956), .Z(n44958) );
  XNOR U5843 ( .A(n44959), .B(n44779), .Z(n44781) );
  XNOR U5844 ( .A(n44782), .B(n44596), .Z(n44598) );
  XNOR U5845 ( .A(n44599), .B(n44407), .Z(n44409) );
  XNOR U5846 ( .A(n44410), .B(n44212), .Z(n44214) );
  XNOR U5847 ( .A(n44215), .B(n44011), .Z(n44013) );
  XNOR U5848 ( .A(n44014), .B(n43804), .Z(n43806) );
  XNOR U5849 ( .A(n43807), .B(n43591), .Z(n43593) );
  XNOR U5850 ( .A(n43594), .B(n43372), .Z(n43374) );
  XNOR U5851 ( .A(n43375), .B(n43147), .Z(n43149) );
  XNOR U5852 ( .A(n43150), .B(n42916), .Z(n42918) );
  XNOR U5853 ( .A(n42919), .B(n42679), .Z(n42681) );
  XNOR U5854 ( .A(n42682), .B(n42436), .Z(n42438) );
  XNOR U5855 ( .A(n42439), .B(n42187), .Z(n42189) );
  XNOR U5856 ( .A(n42190), .B(n41932), .Z(n41934) );
  XNOR U5857 ( .A(n41935), .B(n41671), .Z(n41673) );
  XNOR U5858 ( .A(n41674), .B(n41404), .Z(n41406) );
  XNOR U5859 ( .A(n41407), .B(n41131), .Z(n41133) );
  XNOR U5860 ( .A(n41134), .B(n40852), .Z(n40854) );
  XNOR U5861 ( .A(n40855), .B(n40567), .Z(n40569) );
  XNOR U5862 ( .A(n40570), .B(n40276), .Z(n40278) );
  XNOR U5863 ( .A(n40279), .B(n39979), .Z(n39981) );
  XNOR U5864 ( .A(n39982), .B(n39676), .Z(n39678) );
  XNOR U5865 ( .A(n39679), .B(n39367), .Z(n39369) );
  XNOR U5866 ( .A(n39370), .B(n39052), .Z(n39054) );
  XNOR U5867 ( .A(n39055), .B(n38731), .Z(n38733) );
  XNOR U5868 ( .A(n38734), .B(n38404), .Z(n38406) );
  XNOR U5869 ( .A(n38407), .B(n38071), .Z(n38073) );
  XNOR U5870 ( .A(n38074), .B(n37732), .Z(n37734) );
  XNOR U5871 ( .A(n37735), .B(n37387), .Z(n37389) );
  XNOR U5872 ( .A(n37390), .B(n37036), .Z(n37038) );
  XNOR U5873 ( .A(n37039), .B(n36679), .Z(n36681) );
  XNOR U5874 ( .A(n36682), .B(n36316), .Z(n36318) );
  XNOR U5875 ( .A(n36319), .B(n35947), .Z(n35949) );
  XNOR U5876 ( .A(n35950), .B(n35572), .Z(n35574) );
  XNOR U5877 ( .A(n35575), .B(n35191), .Z(n35193) );
  XNOR U5878 ( .A(n35194), .B(n34804), .Z(n34806) );
  XNOR U5879 ( .A(n34807), .B(n34411), .Z(n34413) );
  XNOR U5880 ( .A(n34414), .B(n34012), .Z(n34014) );
  XNOR U5881 ( .A(n34015), .B(n33607), .Z(n33609) );
  XNOR U5882 ( .A(n33610), .B(n33196), .Z(n33198) );
  XNOR U5883 ( .A(n33199), .B(n32779), .Z(n32781) );
  XNOR U5884 ( .A(n32782), .B(n32356), .Z(n32358) );
  XNOR U5885 ( .A(n32359), .B(n31927), .Z(n31929) );
  XNOR U5886 ( .A(n31930), .B(n31492), .Z(n31494) );
  XNOR U5887 ( .A(n31495), .B(n31051), .Z(n31053) );
  XNOR U5888 ( .A(n31054), .B(n30604), .Z(n30606) );
  XNOR U5889 ( .A(n30607), .B(n30151), .Z(n30153) );
  XNOR U5890 ( .A(n30154), .B(n29692), .Z(n29694) );
  XNOR U5891 ( .A(n29695), .B(n29227), .Z(n29229) );
  XNOR U5892 ( .A(n29230), .B(n28756), .Z(n28758) );
  XNOR U5893 ( .A(n28759), .B(n28279), .Z(n28281) );
  XNOR U5894 ( .A(n28282), .B(n27796), .Z(n27798) );
  XNOR U5895 ( .A(n27799), .B(n27307), .Z(n27309) );
  XNOR U5896 ( .A(n27310), .B(n26810), .Z(n26812) );
  XNOR U5897 ( .A(n26813), .B(n26309), .Z(n26311) );
  XNOR U5898 ( .A(n26312), .B(n25801), .Z(n25803) );
  XNOR U5899 ( .A(n25804), .B(n25287), .Z(n25289) );
  XNOR U5900 ( .A(n25290), .B(n24764), .Z(n24766) );
  XNOR U5901 ( .A(n24767), .B(n24239), .Z(n24241) );
  XNOR U5902 ( .A(n24242), .B(n23708), .Z(n23710) );
  XNOR U5903 ( .A(n23711), .B(n23170), .Z(n23172) );
  XNOR U5904 ( .A(n23173), .B(n22626), .Z(n22628) );
  XNOR U5905 ( .A(n22629), .B(n22077), .Z(n22079) );
  XNOR U5906 ( .A(n22080), .B(n21522), .Z(n21524) );
  XNOR U5907 ( .A(n21525), .B(n20960), .Z(n20962) );
  XNOR U5908 ( .A(n20963), .B(n20393), .Z(n20395) );
  XNOR U5909 ( .A(n20396), .B(n19820), .Z(n19822) );
  XNOR U5910 ( .A(n19823), .B(n19241), .Z(n19243) );
  XOR U5911 ( .A(n18549), .B(n18599), .Z(n18553) );
  XOR U5912 ( .A(n16145), .B(n16184), .Z(n16149) );
  XOR U5913 ( .A(n14907), .B(n14946), .Z(n14911) );
  XOR U5914 ( .A(n13645), .B(n13684), .Z(n13649) );
  XOR U5915 ( .A(n12357), .B(n12398), .Z(n12361) );
  XOR U5916 ( .A(n11047), .B(n11086), .Z(n11051) );
  XOR U5917 ( .A(n9713), .B(n9752), .Z(n9717) );
  XOR U5918 ( .A(n8355), .B(n8394), .Z(n8359) );
  XOR U5919 ( .A(n6973), .B(n7012), .Z(n6977) );
  XOR U5920 ( .A(n5565), .B(n5606), .Z(n5569) );
  XOR U5921 ( .A(n4135), .B(n4174), .Z(n4139) );
  XOR U5922 ( .A(n2681), .B(n2720), .Z(n2685) );
  XNOR U5923 ( .A(n47187), .B(n47121), .Z(n47123) );
  XOR U5924 ( .A(n17962), .B(n17995), .Z(n17966) );
  XOR U5925 ( .A(n47242), .B(n47268), .Z(n47246) );
  XNOR U5926 ( .A(n47469), .B(n47445), .Z(n47447) );
  XNOR U5927 ( .A(n47448), .B(n47418), .Z(n47420) );
  XNOR U5928 ( .A(n47421), .B(n47385), .Z(n47387) );
  XNOR U5929 ( .A(n47388), .B(n47346), .Z(n47348) );
  XNOR U5930 ( .A(n47197), .B(n47131), .Z(n47133) );
  XNOR U5931 ( .A(n47134), .B(n47062), .Z(n47064) );
  XNOR U5932 ( .A(n47065), .B(n46987), .Z(n46989) );
  XNOR U5933 ( .A(n46990), .B(n46906), .Z(n46908) );
  XNOR U5934 ( .A(n46909), .B(n46819), .Z(n46821) );
  XNOR U5935 ( .A(n46822), .B(n46726), .Z(n46728) );
  XNOR U5936 ( .A(n46729), .B(n46627), .Z(n46629) );
  XNOR U5937 ( .A(n46630), .B(n46522), .Z(n46524) );
  XNOR U5938 ( .A(n46525), .B(n46411), .Z(n46413) );
  XNOR U5939 ( .A(n46414), .B(n46294), .Z(n46296) );
  XNOR U5940 ( .A(n46297), .B(n46171), .Z(n46173) );
  XNOR U5941 ( .A(n46174), .B(n46042), .Z(n46044) );
  XNOR U5942 ( .A(n46045), .B(n45907), .Z(n45909) );
  XNOR U5943 ( .A(n45910), .B(n45766), .Z(n45768) );
  XNOR U5944 ( .A(n45769), .B(n45619), .Z(n45621) );
  XNOR U5945 ( .A(n45622), .B(n45466), .Z(n45468) );
  XNOR U5946 ( .A(n45469), .B(n45307), .Z(n45309) );
  XNOR U5947 ( .A(n45310), .B(n45142), .Z(n45144) );
  XNOR U5948 ( .A(n45145), .B(n44971), .Z(n44973) );
  XNOR U5949 ( .A(n44974), .B(n44794), .Z(n44796) );
  XNOR U5950 ( .A(n44797), .B(n44611), .Z(n44613) );
  XNOR U5951 ( .A(n44614), .B(n44422), .Z(n44424) );
  XNOR U5952 ( .A(n44425), .B(n44227), .Z(n44229) );
  XNOR U5953 ( .A(n44230), .B(n44026), .Z(n44028) );
  XNOR U5954 ( .A(n44029), .B(n43819), .Z(n43821) );
  XNOR U5955 ( .A(n43822), .B(n43606), .Z(n43608) );
  XNOR U5956 ( .A(n43609), .B(n43387), .Z(n43389) );
  XNOR U5957 ( .A(n43390), .B(n43162), .Z(n43164) );
  XNOR U5958 ( .A(n43165), .B(n42931), .Z(n42933) );
  XNOR U5959 ( .A(n42934), .B(n42694), .Z(n42696) );
  XNOR U5960 ( .A(n42697), .B(n42451), .Z(n42453) );
  XNOR U5961 ( .A(n42454), .B(n42202), .Z(n42204) );
  XNOR U5962 ( .A(n42205), .B(n41947), .Z(n41949) );
  XNOR U5963 ( .A(n41950), .B(n41686), .Z(n41688) );
  XNOR U5964 ( .A(n41689), .B(n41419), .Z(n41421) );
  XNOR U5965 ( .A(n41422), .B(n41146), .Z(n41148) );
  XNOR U5966 ( .A(n41149), .B(n40867), .Z(n40869) );
  XNOR U5967 ( .A(n40870), .B(n40582), .Z(n40584) );
  XNOR U5968 ( .A(n40585), .B(n40291), .Z(n40293) );
  XNOR U5969 ( .A(n40294), .B(n39994), .Z(n39996) );
  XNOR U5970 ( .A(n39997), .B(n39691), .Z(n39693) );
  XNOR U5971 ( .A(n39694), .B(n39382), .Z(n39384) );
  XNOR U5972 ( .A(n39385), .B(n39067), .Z(n39069) );
  XNOR U5973 ( .A(n39070), .B(n38746), .Z(n38748) );
  XNOR U5974 ( .A(n38749), .B(n38419), .Z(n38421) );
  XNOR U5975 ( .A(n38422), .B(n38086), .Z(n38088) );
  XNOR U5976 ( .A(n38089), .B(n37747), .Z(n37749) );
  XNOR U5977 ( .A(n37750), .B(n37402), .Z(n37404) );
  XNOR U5978 ( .A(n37405), .B(n37051), .Z(n37053) );
  XNOR U5979 ( .A(n37054), .B(n36694), .Z(n36696) );
  XNOR U5980 ( .A(n36697), .B(n36331), .Z(n36333) );
  XNOR U5981 ( .A(n36334), .B(n35962), .Z(n35964) );
  XNOR U5982 ( .A(n35965), .B(n35587), .Z(n35589) );
  XNOR U5983 ( .A(n35590), .B(n35206), .Z(n35208) );
  XNOR U5984 ( .A(n35209), .B(n34819), .Z(n34821) );
  XNOR U5985 ( .A(n34822), .B(n34426), .Z(n34428) );
  XNOR U5986 ( .A(n34429), .B(n34027), .Z(n34029) );
  XNOR U5987 ( .A(n34030), .B(n33622), .Z(n33624) );
  XNOR U5988 ( .A(n33625), .B(n33211), .Z(n33213) );
  XNOR U5989 ( .A(n33214), .B(n32794), .Z(n32796) );
  XNOR U5990 ( .A(n32797), .B(n32371), .Z(n32373) );
  XNOR U5991 ( .A(n32374), .B(n31942), .Z(n31944) );
  XNOR U5992 ( .A(n31945), .B(n31507), .Z(n31509) );
  XNOR U5993 ( .A(n31510), .B(n31066), .Z(n31068) );
  XNOR U5994 ( .A(n31069), .B(n30619), .Z(n30621) );
  XNOR U5995 ( .A(n30622), .B(n30166), .Z(n30168) );
  XNOR U5996 ( .A(n30169), .B(n29707), .Z(n29709) );
  XNOR U5997 ( .A(n29710), .B(n29242), .Z(n29244) );
  XNOR U5998 ( .A(n29245), .B(n28771), .Z(n28773) );
  XNOR U5999 ( .A(n28774), .B(n28294), .Z(n28296) );
  XNOR U6000 ( .A(n28297), .B(n27811), .Z(n27813) );
  XNOR U6001 ( .A(n27814), .B(n27322), .Z(n27324) );
  XNOR U6002 ( .A(n27325), .B(n26825), .Z(n26827) );
  XNOR U6003 ( .A(n26828), .B(n26324), .Z(n26326) );
  XNOR U6004 ( .A(n26327), .B(n25816), .Z(n25818) );
  XNOR U6005 ( .A(n25819), .B(n25302), .Z(n25304) );
  XNOR U6006 ( .A(n25305), .B(n24779), .Z(n24781) );
  XNOR U6007 ( .A(n24782), .B(n24254), .Z(n24256) );
  XNOR U6008 ( .A(n24257), .B(n23723), .Z(n23725) );
  XNOR U6009 ( .A(n23726), .B(n23185), .Z(n23187) );
  XNOR U6010 ( .A(n23188), .B(n22641), .Z(n22643) );
  XNOR U6011 ( .A(n22644), .B(n22092), .Z(n22094) );
  XNOR U6012 ( .A(n22095), .B(n21537), .Z(n21539) );
  XNOR U6013 ( .A(n21540), .B(n20975), .Z(n20977) );
  XNOR U6014 ( .A(n20978), .B(n20408), .Z(n20410) );
  XNOR U6015 ( .A(n20411), .B(n19835), .Z(n19837) );
  XOR U6016 ( .A(n17374), .B(n17395), .Z(n17378) );
  XOR U6017 ( .A(n16160), .B(n16181), .Z(n16164) );
  XOR U6018 ( .A(n14922), .B(n14943), .Z(n14926) );
  XOR U6019 ( .A(n13660), .B(n13681), .Z(n13664) );
  XOR U6020 ( .A(n12372), .B(n12395), .Z(n12376) );
  XOR U6021 ( .A(n11062), .B(n11083), .Z(n11066) );
  XOR U6022 ( .A(n9728), .B(n9749), .Z(n9732) );
  XOR U6023 ( .A(n8370), .B(n8391), .Z(n8374) );
  XOR U6024 ( .A(n6988), .B(n7009), .Z(n6992) );
  XOR U6025 ( .A(n5580), .B(n5603), .Z(n5584) );
  XOR U6026 ( .A(n4150), .B(n4171), .Z(n4154) );
  XOR U6027 ( .A(n2696), .B(n2717), .Z(n2700) );
  XOR U6028 ( .A(n47303), .B(n47308), .Z(n47263) );
  XNOR U6029 ( .A(n47256), .B(n47255), .Z(n47206) );
  XOR U6030 ( .A(n19258), .B(n19263), .Z(n18588) );
  XOR U6031 ( .A(n18569), .B(n18583), .Z(n18574) );
  XOR U6032 ( .A(n26929), .B(n27417), .Z(n26933) );
  XOR U6033 ( .A(n28869), .B(n29333), .Z(n28873) );
  XOR U6034 ( .A(n28398), .B(n28862), .Z(n28402) );
  XOR U6035 ( .A(n27921), .B(n28385), .Z(n27925) );
  XNOR U6036 ( .A(n26955), .B(n26455), .Z(n26457) );
  XNOR U6037 ( .A(n27927), .B(n27441), .Z(n27443) );
  XNOR U6038 ( .A(n26935), .B(n26435), .Z(n26437) );
  XNOR U6039 ( .A(n26940), .B(n26440), .Z(n26442) );
  XOR U6040 ( .A(n25408), .B(n25915), .Z(n25412) );
  XNOR U6041 ( .A(n26458), .B(n25954), .Z(n25956) );
  XOR U6042 ( .A(n30261), .B(n30707), .Z(n30265) );
  XOR U6043 ( .A(n29808), .B(n30254), .Z(n29812) );
  XOR U6044 ( .A(n29349), .B(n29795), .Z(n29353) );
  XOR U6045 ( .A(n28884), .B(n29330), .Z(n28888) );
  XOR U6046 ( .A(n28413), .B(n28859), .Z(n28417) );
  XOR U6047 ( .A(n27453), .B(n27899), .Z(n27457) );
  XNOR U6048 ( .A(n27459), .B(n26967), .Z(n26969) );
  XNOR U6049 ( .A(n25434), .B(n24916), .Z(n24918) );
  XNOR U6050 ( .A(n26950), .B(n26450), .Z(n26452) );
  XNOR U6051 ( .A(n26443), .B(n25939), .Z(n25941) );
  XNOR U6052 ( .A(n25414), .B(n24896), .Z(n24898) );
  XNOR U6053 ( .A(n26468), .B(n25964), .Z(n25966) );
  XNOR U6054 ( .A(n25957), .B(n25446), .Z(n25448) );
  XNOR U6055 ( .A(n25419), .B(n24901), .Z(n24903) );
  XOR U6056 ( .A(n23831), .B(n24355), .Z(n23835) );
  XNOR U6057 ( .A(n25464), .B(n24946), .Z(n24948) );
  XNOR U6058 ( .A(n24919), .B(n24394), .Z(n24396) );
  XNOR U6059 ( .A(n25469), .B(n24951), .Z(n24953) );
  XOR U6060 ( .A(n31599), .B(n32027), .Z(n31603) );
  XOR U6061 ( .A(n31164), .B(n31592), .Z(n31168) );
  XOR U6062 ( .A(n30723), .B(n31151), .Z(n30727) );
  XOR U6063 ( .A(n30276), .B(n30704), .Z(n30280) );
  XOR U6064 ( .A(n29823), .B(n30251), .Z(n29827) );
  XOR U6065 ( .A(n28899), .B(n29327), .Z(n28903) );
  XOR U6066 ( .A(n28428), .B(n28856), .Z(n28432) );
  XOR U6067 ( .A(n27951), .B(n28379), .Z(n27955) );
  XOR U6068 ( .A(n27468), .B(n27896), .Z(n27472) );
  XOR U6069 ( .A(n26482), .B(n26910), .Z(n26486) );
  XNOR U6070 ( .A(n26478), .B(n25974), .Z(n25976) );
  XNOR U6071 ( .A(n23857), .B(n23323), .Z(n23325) );
  XNOR U6072 ( .A(n25429), .B(n24911), .Z(n24913) );
  XNOR U6073 ( .A(n24904), .B(n24379), .Z(n24381) );
  XNOR U6074 ( .A(n23837), .B(n23303), .Z(n23305) );
  XNOR U6075 ( .A(n25474), .B(n24956), .Z(n24958) );
  XOR U6076 ( .A(n24933), .B(n25393), .Z(n24937) );
  XNOR U6077 ( .A(n24929), .B(n24404), .Z(n24406) );
  XNOR U6078 ( .A(n24397), .B(n23869), .Z(n23871) );
  XNOR U6079 ( .A(n23842), .B(n23308), .Z(n23310) );
  XOR U6080 ( .A(n22203), .B(n22746), .Z(n22207) );
  XNOR U6081 ( .A(n23326), .B(n22785), .Z(n22787) );
  XOR U6082 ( .A(n23355), .B(n23813), .Z(n23359) );
  XOR U6083 ( .A(n32883), .B(n33293), .Z(n32887) );
  XOR U6084 ( .A(n32466), .B(n32876), .Z(n32470) );
  XOR U6085 ( .A(n32043), .B(n32453), .Z(n32047) );
  XOR U6086 ( .A(n31614), .B(n32024), .Z(n31618) );
  XOR U6087 ( .A(n31179), .B(n31589), .Z(n31183) );
  XOR U6088 ( .A(n30291), .B(n30701), .Z(n30295) );
  XOR U6089 ( .A(n29838), .B(n30248), .Z(n29842) );
  XOR U6090 ( .A(n29379), .B(n29789), .Z(n29383) );
  XOR U6091 ( .A(n28914), .B(n29324), .Z(n28918) );
  XOR U6092 ( .A(n28443), .B(n28853), .Z(n28447) );
  XOR U6093 ( .A(n27966), .B(n28376), .Z(n27970) );
  XOR U6094 ( .A(n27483), .B(n27893), .Z(n27487) );
  XOR U6095 ( .A(n26994), .B(n27404), .Z(n26998) );
  XOR U6096 ( .A(n26497), .B(n26907), .Z(n26501) );
  XOR U6097 ( .A(n25996), .B(n26406), .Z(n26000) );
  XOR U6098 ( .A(n24973), .B(n25384), .Z(n24977) );
  XNOR U6099 ( .A(n24939), .B(n24414), .Z(n24416) );
  XNOR U6100 ( .A(n22229), .B(n21677), .Z(n21679) );
  XNOR U6101 ( .A(n23852), .B(n23318), .Z(n23320) );
  XNOR U6102 ( .A(n23311), .B(n22770), .Z(n22772) );
  XNOR U6103 ( .A(n22209), .B(n21657), .Z(n21659) );
  XOR U6104 ( .A(n23901), .B(n24341), .Z(n23905) );
  XOR U6105 ( .A(n23385), .B(n23807), .Z(n23389) );
  XOR U6106 ( .A(n23340), .B(n23816), .Z(n23344) );
  XNOR U6107 ( .A(n23336), .B(n22795), .Z(n22797) );
  XNOR U6108 ( .A(n22788), .B(n22241), .Z(n22243) );
  XNOR U6109 ( .A(n22214), .B(n21662), .Z(n21664) );
  XOR U6110 ( .A(n20522), .B(n21083), .Z(n20526) );
  XOR U6111 ( .A(n24441), .B(n24866), .Z(n24445) );
  XNOR U6112 ( .A(n21680), .B(n21122), .Z(n21124) );
  XOR U6113 ( .A(n23370), .B(n23810), .Z(n23374) );
  XOR U6114 ( .A(n21709), .B(n22185), .Z(n21713) );
  XOR U6115 ( .A(n34113), .B(n34505), .Z(n34117) );
  XOR U6116 ( .A(n33714), .B(n34106), .Z(n33718) );
  XOR U6117 ( .A(n33309), .B(n33701), .Z(n33313) );
  XOR U6118 ( .A(n32898), .B(n33290), .Z(n32902) );
  XOR U6119 ( .A(n32481), .B(n32873), .Z(n32485) );
  XOR U6120 ( .A(n31629), .B(n32021), .Z(n31633) );
  XOR U6121 ( .A(n31194), .B(n31586), .Z(n31198) );
  XOR U6122 ( .A(n30753), .B(n31145), .Z(n30757) );
  XOR U6123 ( .A(n30306), .B(n30698), .Z(n30310) );
  XOR U6124 ( .A(n29853), .B(n30245), .Z(n29857) );
  XOR U6125 ( .A(n29394), .B(n29786), .Z(n29398) );
  XOR U6126 ( .A(n28929), .B(n29321), .Z(n28933) );
  XOR U6127 ( .A(n28458), .B(n28850), .Z(n28462) );
  XOR U6128 ( .A(n27981), .B(n28373), .Z(n27985) );
  XOR U6129 ( .A(n27498), .B(n27890), .Z(n27502) );
  XOR U6130 ( .A(n27009), .B(n27401), .Z(n27013) );
  XOR U6131 ( .A(n26512), .B(n26904), .Z(n26516) );
  XOR U6132 ( .A(n26011), .B(n26403), .Z(n26015) );
  XOR U6133 ( .A(n25503), .B(n25895), .Z(n25507) );
  XOR U6134 ( .A(n24988), .B(n25381), .Z(n24993) );
  XNOR U6135 ( .A(n23346), .B(n22805), .Z(n22807) );
  XNOR U6136 ( .A(n20548), .B(n19978), .Z(n19980) );
  XNOR U6137 ( .A(n22224), .B(n21672), .Z(n21674) );
  XNOR U6138 ( .A(n21665), .B(n21107), .Z(n21109) );
  XNOR U6139 ( .A(n20528), .B(n19958), .Z(n19960) );
  XOR U6140 ( .A(n22273), .B(n22732), .Z(n22277) );
  XOR U6141 ( .A(n23400), .B(n23804), .Z(n23404) );
  XOR U6142 ( .A(n22852), .B(n23269), .Z(n22856) );
  XOR U6143 ( .A(n21739), .B(n22179), .Z(n21743) );
  XOR U6144 ( .A(n21694), .B(n22188), .Z(n21698) );
  XNOR U6145 ( .A(n21690), .B(n21132), .Z(n21134) );
  XNOR U6146 ( .A(n21125), .B(n20560), .Z(n20562) );
  XNOR U6147 ( .A(n20533), .B(n19963), .Z(n19965) );
  XOR U6148 ( .A(n18788), .B(n19366), .Z(n18792) );
  XOR U6149 ( .A(n22832), .B(n23273), .Z(n22836) );
  XNOR U6150 ( .A(n22319), .B(n21767), .Z(n21769) );
  XOR U6151 ( .A(n21724), .B(n22182), .Z(n21728) );
  XOR U6152 ( .A(n20010), .B(n20504), .Z(n20014) );
  XOR U6153 ( .A(n19427), .B(n19933), .Z(n19431) );
  XOR U6154 ( .A(n22328), .B(n22721), .Z(n22332) );
  XOR U6155 ( .A(n35289), .B(n35663), .Z(n35293) );
  XOR U6156 ( .A(n34908), .B(n35282), .Z(n34912) );
  XOR U6157 ( .A(n34521), .B(n34895), .Z(n34525) );
  XOR U6158 ( .A(n34128), .B(n34502), .Z(n34132) );
  XOR U6159 ( .A(n33729), .B(n34103), .Z(n33733) );
  XOR U6160 ( .A(n32913), .B(n33287), .Z(n32917) );
  XOR U6161 ( .A(n32496), .B(n32870), .Z(n32500) );
  XOR U6162 ( .A(n32073), .B(n32447), .Z(n32077) );
  XOR U6163 ( .A(n31644), .B(n32018), .Z(n31648) );
  XOR U6164 ( .A(n31209), .B(n31583), .Z(n31213) );
  XOR U6165 ( .A(n30768), .B(n31142), .Z(n30772) );
  XOR U6166 ( .A(n30321), .B(n30695), .Z(n30325) );
  XOR U6167 ( .A(n29868), .B(n30242), .Z(n29872) );
  XOR U6168 ( .A(n29409), .B(n29783), .Z(n29413) );
  XOR U6169 ( .A(n28944), .B(n29318), .Z(n28948) );
  XOR U6170 ( .A(n28473), .B(n28847), .Z(n28477) );
  XOR U6171 ( .A(n27996), .B(n28370), .Z(n28000) );
  XOR U6172 ( .A(n27513), .B(n27887), .Z(n27517) );
  XOR U6173 ( .A(n27024), .B(n27398), .Z(n27028) );
  XOR U6174 ( .A(n26527), .B(n26901), .Z(n26531) );
  XOR U6175 ( .A(n26026), .B(n26400), .Z(n26030) );
  XOR U6176 ( .A(n25518), .B(n25892), .Z(n25522) );
  XOR U6177 ( .A(n25004), .B(n25378), .Z(n25008) );
  XOR U6178 ( .A(n24481), .B(n24855), .Z(n24485) );
  XOR U6179 ( .A(n23956), .B(n24330), .Z(n23960) );
  XOR U6180 ( .A(n23425), .B(n23799), .Z(n23429) );
  XNOR U6181 ( .A(n22349), .B(n21797), .Z(n21799) );
  XNOR U6182 ( .A(n23406), .B(n22865), .Z(n22867) );
  XNOR U6183 ( .A(n21700), .B(n21142), .Z(n21144) );
  XOR U6184 ( .A(n18818), .B(n19360), .Z(n18822) );
  XNOR U6185 ( .A(n20543), .B(n19973), .Z(n19975) );
  XOR U6186 ( .A(n20592), .B(n21069), .Z(n20596) );
  XOR U6187 ( .A(n21754), .B(n22176), .Z(n21758) );
  XOR U6188 ( .A(n21189), .B(n21623), .Z(n21193) );
  XOR U6189 ( .A(n20040), .B(n20498), .Z(n20044) );
  XOR U6190 ( .A(n19995), .B(n20507), .Z(n19999) );
  XNOR U6191 ( .A(n19991), .B(n19415), .Z(n19417) );
  XNOR U6192 ( .A(n19408), .B(n18826), .Z(n18828) );
  XOR U6193 ( .A(n18099), .B(n18779), .Z(n18103) );
  XOR U6194 ( .A(n18803), .B(n19363), .Z(n18807) );
  XOR U6195 ( .A(n21169), .B(n21627), .Z(n21173) );
  XOR U6196 ( .A(n21779), .B(n22171), .Z(n21783) );
  XOR U6197 ( .A(n16894), .B(n17491), .Z(n16898) );
  XOR U6198 ( .A(n20025), .B(n20501), .Z(n20029) );
  XNOR U6199 ( .A(n22339), .B(n21787), .Z(n21789) );
  XOR U6200 ( .A(n20647), .B(n21058), .Z(n20651) );
  XOR U6201 ( .A(n19487), .B(n19921), .Z(n19491) );
  XOR U6202 ( .A(n36411), .B(n36767), .Z(n36415) );
  XOR U6203 ( .A(n36048), .B(n36404), .Z(n36052) );
  XOR U6204 ( .A(n35679), .B(n36035), .Z(n35683) );
  XOR U6205 ( .A(n35304), .B(n35660), .Z(n35308) );
  XOR U6206 ( .A(n34923), .B(n35279), .Z(n34927) );
  XOR U6207 ( .A(n34143), .B(n34499), .Z(n34147) );
  XOR U6208 ( .A(n33744), .B(n34100), .Z(n33748) );
  XOR U6209 ( .A(n33339), .B(n33695), .Z(n33343) );
  XOR U6210 ( .A(n32928), .B(n33284), .Z(n32932) );
  XOR U6211 ( .A(n32511), .B(n32867), .Z(n32515) );
  XOR U6212 ( .A(n32088), .B(n32444), .Z(n32092) );
  XOR U6213 ( .A(n31659), .B(n32015), .Z(n31663) );
  XOR U6214 ( .A(n31224), .B(n31580), .Z(n31228) );
  XOR U6215 ( .A(n30783), .B(n31139), .Z(n30787) );
  XOR U6216 ( .A(n30336), .B(n30692), .Z(n30340) );
  XOR U6217 ( .A(n29883), .B(n30239), .Z(n29887) );
  XOR U6218 ( .A(n29424), .B(n29780), .Z(n29428) );
  XOR U6219 ( .A(n28959), .B(n29315), .Z(n28963) );
  XOR U6220 ( .A(n28488), .B(n28844), .Z(n28492) );
  XOR U6221 ( .A(n28011), .B(n28367), .Z(n28015) );
  XOR U6222 ( .A(n27528), .B(n27884), .Z(n27532) );
  XOR U6223 ( .A(n27039), .B(n27395), .Z(n27043) );
  XOR U6224 ( .A(n26542), .B(n26898), .Z(n26546) );
  XOR U6225 ( .A(n26041), .B(n26397), .Z(n26045) );
  XOR U6226 ( .A(n25533), .B(n25889), .Z(n25537) );
  XOR U6227 ( .A(n25019), .B(n25375), .Z(n25023) );
  XOR U6228 ( .A(n24496), .B(n24852), .Z(n24500) );
  XOR U6229 ( .A(n23971), .B(n24327), .Z(n23975) );
  XOR U6230 ( .A(n23440), .B(n23796), .Z(n23444) );
  XOR U6231 ( .A(n22902), .B(n23258), .Z(n22906) );
  XNOR U6232 ( .A(n22908), .B(n22361), .Z(n22363) );
  XOR U6233 ( .A(n21809), .B(n22165), .Z(n21813) );
  XNOR U6234 ( .A(n21760), .B(n21202), .Z(n21204) );
  XOR U6235 ( .A(n18154), .B(n18757), .Z(n18158) );
  XOR U6236 ( .A(n18858), .B(n19352), .Z(n18862) );
  XOR U6237 ( .A(n20677), .B(n21052), .Z(n20681) );
  XOR U6238 ( .A(n19517), .B(n19915), .Z(n19521) );
  XOR U6239 ( .A(n20055), .B(n20495), .Z(n20059) );
  XOR U6240 ( .A(n19472), .B(n19924), .Z(n19476) );
  XOR U6241 ( .A(n18883), .B(n19347), .Z(n18887) );
  XOR U6242 ( .A(n18838), .B(n19356), .Z(n18842) );
  XOR U6243 ( .A(n17532), .B(n18081), .Z(n17536) );
  XOR U6244 ( .A(n18114), .B(n18773), .Z(n18118) );
  XNOR U6245 ( .A(n20031), .B(n19455), .Z(n19457) );
  XNOR U6246 ( .A(n21790), .B(n21232), .Z(n21234) );
  XOR U6247 ( .A(n20080), .B(n20490), .Z(n20084) );
  XNOR U6248 ( .A(n21270), .B(n20705), .Z(n20707) );
  XOR U6249 ( .A(n16315), .B(n16882), .Z(n16319) );
  XOR U6250 ( .A(n16909), .B(n17488), .Z(n16913) );
  XOR U6251 ( .A(n15675), .B(n16278), .Z(n15679) );
  XNOR U6252 ( .A(n20658), .B(n20088), .Z(n20090) );
  XOR U6253 ( .A(n18913), .B(n19341), .Z(n18917) );
  XOR U6254 ( .A(n19547), .B(n19909), .Z(n19551) );
  XOR U6255 ( .A(n37479), .B(n37817), .Z(n37483) );
  XOR U6256 ( .A(n37134), .B(n37472), .Z(n37138) );
  XOR U6257 ( .A(n36783), .B(n37121), .Z(n36787) );
  XOR U6258 ( .A(n36426), .B(n36764), .Z(n36430) );
  XOR U6259 ( .A(n36063), .B(n36401), .Z(n36067) );
  XOR U6260 ( .A(n35319), .B(n35657), .Z(n35323) );
  XOR U6261 ( .A(n34938), .B(n35276), .Z(n34942) );
  XOR U6262 ( .A(n34551), .B(n34889), .Z(n34555) );
  XOR U6263 ( .A(n34158), .B(n34496), .Z(n34162) );
  XOR U6264 ( .A(n33759), .B(n34097), .Z(n33763) );
  XOR U6265 ( .A(n33354), .B(n33692), .Z(n33358) );
  XOR U6266 ( .A(n32943), .B(n33281), .Z(n32947) );
  XOR U6267 ( .A(n32526), .B(n32864), .Z(n32530) );
  XOR U6268 ( .A(n32103), .B(n32441), .Z(n32107) );
  XOR U6269 ( .A(n31674), .B(n32012), .Z(n31678) );
  XOR U6270 ( .A(n31239), .B(n31577), .Z(n31243) );
  XOR U6271 ( .A(n30798), .B(n31136), .Z(n30802) );
  XOR U6272 ( .A(n30351), .B(n30689), .Z(n30355) );
  XOR U6273 ( .A(n29898), .B(n30236), .Z(n29902) );
  XOR U6274 ( .A(n29439), .B(n29777), .Z(n29443) );
  XOR U6275 ( .A(n28974), .B(n29312), .Z(n28978) );
  XOR U6276 ( .A(n28503), .B(n28841), .Z(n28507) );
  XOR U6277 ( .A(n28026), .B(n28364), .Z(n28030) );
  XOR U6278 ( .A(n27543), .B(n27881), .Z(n27547) );
  XOR U6279 ( .A(n27054), .B(n27392), .Z(n27058) );
  XOR U6280 ( .A(n26557), .B(n26895), .Z(n26561) );
  XOR U6281 ( .A(n26056), .B(n26394), .Z(n26060) );
  XOR U6282 ( .A(n25548), .B(n25886), .Z(n25552) );
  XOR U6283 ( .A(n25034), .B(n25372), .Z(n25038) );
  XOR U6284 ( .A(n24511), .B(n24849), .Z(n24515) );
  XOR U6285 ( .A(n23986), .B(n24324), .Z(n23990) );
  XOR U6286 ( .A(n23455), .B(n23793), .Z(n23459) );
  XOR U6287 ( .A(n22917), .B(n23255), .Z(n22921) );
  XOR U6288 ( .A(n21824), .B(n22162), .Z(n21828) );
  XNOR U6289 ( .A(n21275), .B(n20710), .Z(n20712) );
  XNOR U6290 ( .A(n21820), .B(n21262), .Z(n21264) );
  XOR U6291 ( .A(n20110), .B(n20484), .Z(n20114) );
  XOR U6292 ( .A(n14422), .B(n15043), .Z(n14426) );
  XOR U6293 ( .A(n18169), .B(n18751), .Z(n18173) );
  XOR U6294 ( .A(n16959), .B(n17478), .Z(n16963) );
  XNOR U6295 ( .A(n20688), .B(n20118), .Z(n20120) );
  XOR U6296 ( .A(n18943), .B(n19335), .Z(n18947) );
  XOR U6297 ( .A(n18898), .B(n19344), .Z(n18902) );
  XOR U6298 ( .A(n17592), .B(n18069), .Z(n17596) );
  XOR U6299 ( .A(n17547), .B(n18078), .Z(n17551) );
  XOR U6300 ( .A(n15730), .B(n16267), .Z(n15734) );
  XOR U6301 ( .A(n20140), .B(n20478), .Z(n20144) );
  XOR U6302 ( .A(n16330), .B(n16879), .Z(n16334) );
  XOR U6303 ( .A(n15084), .B(n15657), .Z(n15088) );
  XOR U6304 ( .A(n15690), .B(n16275), .Z(n15694) );
  XOR U6305 ( .A(n18928), .B(n19338), .Z(n18932) );
  XOR U6306 ( .A(n18224), .B(n18729), .Z(n18228) );
  XOR U6307 ( .A(n17014), .B(n17467), .Z(n17018) );
  XOR U6308 ( .A(n18973), .B(n19329), .Z(n18977) );
  XOR U6309 ( .A(n38493), .B(n38813), .Z(n38497) );
  XOR U6310 ( .A(n38166), .B(n38486), .Z(n38170) );
  XOR U6311 ( .A(n37833), .B(n38153), .Z(n37837) );
  XOR U6312 ( .A(n37494), .B(n37814), .Z(n37498) );
  XOR U6313 ( .A(n37149), .B(n37469), .Z(n37153) );
  XOR U6314 ( .A(n36441), .B(n36761), .Z(n36445) );
  XOR U6315 ( .A(n36078), .B(n36398), .Z(n36082) );
  XOR U6316 ( .A(n35709), .B(n36029), .Z(n35713) );
  XOR U6317 ( .A(n35334), .B(n35654), .Z(n35338) );
  XOR U6318 ( .A(n34953), .B(n35273), .Z(n34957) );
  XOR U6319 ( .A(n34566), .B(n34886), .Z(n34570) );
  XOR U6320 ( .A(n34173), .B(n34493), .Z(n34177) );
  XOR U6321 ( .A(n33774), .B(n34094), .Z(n33778) );
  XOR U6322 ( .A(n33369), .B(n33689), .Z(n33373) );
  XOR U6323 ( .A(n32958), .B(n33278), .Z(n32962) );
  XOR U6324 ( .A(n32541), .B(n32861), .Z(n32545) );
  XOR U6325 ( .A(n32118), .B(n32438), .Z(n32122) );
  XOR U6326 ( .A(n31689), .B(n32009), .Z(n31693) );
  XOR U6327 ( .A(n31254), .B(n31574), .Z(n31258) );
  XOR U6328 ( .A(n30813), .B(n31133), .Z(n30817) );
  XOR U6329 ( .A(n30366), .B(n30686), .Z(n30370) );
  XOR U6330 ( .A(n29913), .B(n30233), .Z(n29917) );
  XOR U6331 ( .A(n29454), .B(n29774), .Z(n29458) );
  XOR U6332 ( .A(n28989), .B(n29309), .Z(n28993) );
  XOR U6333 ( .A(n28518), .B(n28838), .Z(n28522) );
  XOR U6334 ( .A(n28041), .B(n28361), .Z(n28045) );
  XOR U6335 ( .A(n27558), .B(n27878), .Z(n27562) );
  XOR U6336 ( .A(n27069), .B(n27389), .Z(n27073) );
  XOR U6337 ( .A(n26572), .B(n26892), .Z(n26576) );
  XOR U6338 ( .A(n26071), .B(n26391), .Z(n26075) );
  XOR U6339 ( .A(n25563), .B(n25883), .Z(n25567) );
  XOR U6340 ( .A(n25049), .B(n25369), .Z(n25053) );
  XOR U6341 ( .A(n24526), .B(n24846), .Z(n24530) );
  XOR U6342 ( .A(n24001), .B(n24321), .Z(n24005) );
  XOR U6343 ( .A(n23470), .B(n23790), .Z(n23474) );
  XOR U6344 ( .A(n22932), .B(n23252), .Z(n22936) );
  XOR U6345 ( .A(n22388), .B(n22708), .Z(n22392) );
  XOR U6346 ( .A(n21839), .B(n22159), .Z(n21843) );
  XOR U6347 ( .A(n21284), .B(n21604), .Z(n21288) );
  XOR U6348 ( .A(n20155), .B(n20475), .Z(n20159) );
  XNOR U6349 ( .A(n19583), .B(n19001), .Z(n19003) );
  XOR U6350 ( .A(n13819), .B(n14410), .Z(n13823) );
  XOR U6351 ( .A(n14437), .B(n15040), .Z(n14441) );
  XOR U6352 ( .A(n13155), .B(n13782), .Z(n13159) );
  XOR U6353 ( .A(n16974), .B(n17475), .Z(n16978) );
  XOR U6354 ( .A(n18958), .B(n19332), .Z(n18962) );
  XOR U6355 ( .A(n18254), .B(n18717), .Z(n18258) );
  XOR U6356 ( .A(n17044), .B(n17461), .Z(n17048) );
  XOR U6357 ( .A(n17607), .B(n18066), .Z(n17611) );
  XOR U6358 ( .A(n16385), .B(n16868), .Z(n16389) );
  XOR U6359 ( .A(n15139), .B(n15646), .Z(n15143) );
  XOR U6360 ( .A(n11852), .B(n12499), .Z(n11856) );
  XOR U6361 ( .A(n15745), .B(n16264), .Z(n15749) );
  XOR U6362 ( .A(n14487), .B(n15030), .Z(n14491) );
  XOR U6363 ( .A(n15099), .B(n15654), .Z(n15103) );
  XOR U6364 ( .A(n13210), .B(n13771), .Z(n13214) );
  XOR U6365 ( .A(n17637), .B(n18060), .Z(n17641) );
  XOR U6366 ( .A(n16415), .B(n16862), .Z(n16419) );
  XOR U6367 ( .A(n15169), .B(n15640), .Z(n15173) );
  XOR U6368 ( .A(n18988), .B(n19326), .Z(n18992) );
  XOR U6369 ( .A(n18284), .B(n18705), .Z(n18288) );
  XOR U6370 ( .A(n17074), .B(n17455), .Z(n17078) );
  XOR U6371 ( .A(n39453), .B(n39755), .Z(n39457) );
  XOR U6372 ( .A(n39144), .B(n39446), .Z(n39148) );
  XOR U6373 ( .A(n38829), .B(n39131), .Z(n38833) );
  XOR U6374 ( .A(n38508), .B(n38810), .Z(n38512) );
  XOR U6375 ( .A(n38181), .B(n38483), .Z(n38185) );
  XOR U6376 ( .A(n37509), .B(n37811), .Z(n37513) );
  XOR U6377 ( .A(n37164), .B(n37466), .Z(n37168) );
  XOR U6378 ( .A(n36813), .B(n37115), .Z(n36817) );
  XOR U6379 ( .A(n36456), .B(n36758), .Z(n36460) );
  XOR U6380 ( .A(n36093), .B(n36395), .Z(n36097) );
  XOR U6381 ( .A(n35724), .B(n36026), .Z(n35728) );
  XOR U6382 ( .A(n35349), .B(n35651), .Z(n35353) );
  XOR U6383 ( .A(n34968), .B(n35270), .Z(n34972) );
  XOR U6384 ( .A(n34581), .B(n34883), .Z(n34585) );
  XOR U6385 ( .A(n34188), .B(n34490), .Z(n34192) );
  XOR U6386 ( .A(n33789), .B(n34091), .Z(n33793) );
  XOR U6387 ( .A(n33384), .B(n33686), .Z(n33388) );
  XOR U6388 ( .A(n32973), .B(n33275), .Z(n32977) );
  XOR U6389 ( .A(n32556), .B(n32858), .Z(n32560) );
  XOR U6390 ( .A(n32133), .B(n32435), .Z(n32137) );
  XOR U6391 ( .A(n31704), .B(n32006), .Z(n31708) );
  XOR U6392 ( .A(n31269), .B(n31571), .Z(n31273) );
  XOR U6393 ( .A(n30828), .B(n31130), .Z(n30832) );
  XOR U6394 ( .A(n30381), .B(n30683), .Z(n30385) );
  XOR U6395 ( .A(n29928), .B(n30230), .Z(n29932) );
  XOR U6396 ( .A(n29469), .B(n29771), .Z(n29473) );
  XOR U6397 ( .A(n29004), .B(n29306), .Z(n29008) );
  XOR U6398 ( .A(n28533), .B(n28835), .Z(n28537) );
  XOR U6399 ( .A(n28056), .B(n28358), .Z(n28060) );
  XOR U6400 ( .A(n27573), .B(n27875), .Z(n27577) );
  XOR U6401 ( .A(n27084), .B(n27386), .Z(n27088) );
  XOR U6402 ( .A(n26587), .B(n26889), .Z(n26591) );
  XOR U6403 ( .A(n26086), .B(n26388), .Z(n26090) );
  XOR U6404 ( .A(n25578), .B(n25880), .Z(n25582) );
  XOR U6405 ( .A(n25064), .B(n25366), .Z(n25068) );
  XOR U6406 ( .A(n24541), .B(n24843), .Z(n24545) );
  XOR U6407 ( .A(n24016), .B(n24318), .Z(n24020) );
  XOR U6408 ( .A(n23485), .B(n23787), .Z(n23489) );
  XOR U6409 ( .A(n22947), .B(n23249), .Z(n22951) );
  XOR U6410 ( .A(n22403), .B(n22705), .Z(n22407) );
  XOR U6411 ( .A(n21854), .B(n22156), .Z(n21858) );
  XOR U6412 ( .A(n21299), .B(n21601), .Z(n21303) );
  XOR U6413 ( .A(n20737), .B(n21039), .Z(n20741) );
  XOR U6414 ( .A(n20170), .B(n20472), .Z(n20174) );
  XOR U6415 ( .A(n13834), .B(n14407), .Z(n13838) );
  XOR U6416 ( .A(n12540), .B(n13137), .Z(n12544) );
  XOR U6417 ( .A(n13170), .B(n13779), .Z(n13174) );
  XOR U6418 ( .A(n19018), .B(n19320), .Z(n19022) );
  XOR U6419 ( .A(n18314), .B(n18693), .Z(n18318) );
  XOR U6420 ( .A(n17104), .B(n17449), .Z(n17108) );
  XOR U6421 ( .A(n17667), .B(n18054), .Z(n17671) );
  XOR U6422 ( .A(n16445), .B(n16856), .Z(n16449) );
  XOR U6423 ( .A(n15199), .B(n15634), .Z(n15203) );
  XOR U6424 ( .A(n15780), .B(n16257), .Z(n15784) );
  XOR U6425 ( .A(n14522), .B(n15023), .Z(n14526) );
  XOR U6426 ( .A(n13240), .B(n13765), .Z(n13244) );
  XOR U6427 ( .A(n11225), .B(n11840), .Z(n11229) );
  XOR U6428 ( .A(n11867), .B(n12496), .Z(n11871) );
  XOR U6429 ( .A(n10537), .B(n11188), .Z(n10541) );
  XOR U6430 ( .A(n14502), .B(n15027), .Z(n14506) );
  XOR U6431 ( .A(n9188), .B(n9857), .Z(n9192) );
  XOR U6432 ( .A(n12575), .B(n13130), .Z(n12579) );
  XOR U6433 ( .A(n11255), .B(n11834), .Z(n11259) );
  XOR U6434 ( .A(n15810), .B(n16251), .Z(n15814) );
  XOR U6435 ( .A(n14552), .B(n15017), .Z(n14556) );
  XOR U6436 ( .A(n13270), .B(n13759), .Z(n13274) );
  XOR U6437 ( .A(n17697), .B(n18048), .Z(n17701) );
  XOR U6438 ( .A(n16475), .B(n16850), .Z(n16479) );
  XOR U6439 ( .A(n15229), .B(n15628), .Z(n15233) );
  XOR U6440 ( .A(n17134), .B(n17443), .Z(n17138) );
  XOR U6441 ( .A(n40359), .B(n40643), .Z(n40363) );
  XOR U6442 ( .A(n40068), .B(n40352), .Z(n40072) );
  XOR U6443 ( .A(n39771), .B(n40055), .Z(n39775) );
  XOR U6444 ( .A(n39468), .B(n39752), .Z(n39472) );
  XOR U6445 ( .A(n39159), .B(n39443), .Z(n39163) );
  XOR U6446 ( .A(n38523), .B(n38807), .Z(n38527) );
  XOR U6447 ( .A(n38196), .B(n38480), .Z(n38200) );
  XOR U6448 ( .A(n37863), .B(n38147), .Z(n37867) );
  XOR U6449 ( .A(n37524), .B(n37808), .Z(n37528) );
  XOR U6450 ( .A(n37179), .B(n37463), .Z(n37183) );
  XOR U6451 ( .A(n36828), .B(n37112), .Z(n36832) );
  XOR U6452 ( .A(n36471), .B(n36755), .Z(n36475) );
  XOR U6453 ( .A(n36108), .B(n36392), .Z(n36112) );
  XOR U6454 ( .A(n35739), .B(n36023), .Z(n35743) );
  XOR U6455 ( .A(n35364), .B(n35648), .Z(n35368) );
  XOR U6456 ( .A(n34983), .B(n35267), .Z(n34987) );
  XOR U6457 ( .A(n34596), .B(n34880), .Z(n34600) );
  XOR U6458 ( .A(n34203), .B(n34487), .Z(n34207) );
  XOR U6459 ( .A(n33804), .B(n34088), .Z(n33808) );
  XOR U6460 ( .A(n33399), .B(n33683), .Z(n33403) );
  XOR U6461 ( .A(n32988), .B(n33272), .Z(n32992) );
  XOR U6462 ( .A(n32571), .B(n32855), .Z(n32575) );
  XOR U6463 ( .A(n32148), .B(n32432), .Z(n32152) );
  XOR U6464 ( .A(n31719), .B(n32003), .Z(n31723) );
  XOR U6465 ( .A(n31284), .B(n31568), .Z(n31288) );
  XOR U6466 ( .A(n30843), .B(n31127), .Z(n30847) );
  XOR U6467 ( .A(n30396), .B(n30680), .Z(n30400) );
  XOR U6468 ( .A(n29943), .B(n30227), .Z(n29947) );
  XOR U6469 ( .A(n29484), .B(n29768), .Z(n29488) );
  XOR U6470 ( .A(n29019), .B(n29303), .Z(n29023) );
  XOR U6471 ( .A(n28548), .B(n28832), .Z(n28552) );
  XOR U6472 ( .A(n28071), .B(n28355), .Z(n28075) );
  XOR U6473 ( .A(n27588), .B(n27872), .Z(n27592) );
  XOR U6474 ( .A(n27099), .B(n27383), .Z(n27103) );
  XOR U6475 ( .A(n26602), .B(n26886), .Z(n26606) );
  XOR U6476 ( .A(n26101), .B(n26385), .Z(n26105) );
  XOR U6477 ( .A(n25593), .B(n25877), .Z(n25597) );
  XOR U6478 ( .A(n25079), .B(n25363), .Z(n25083) );
  XOR U6479 ( .A(n24556), .B(n24840), .Z(n24560) );
  XOR U6480 ( .A(n24031), .B(n24315), .Z(n24035) );
  XOR U6481 ( .A(n23500), .B(n23784), .Z(n23504) );
  XOR U6482 ( .A(n22962), .B(n23246), .Z(n22966) );
  XOR U6483 ( .A(n22418), .B(n22702), .Z(n22422) );
  XOR U6484 ( .A(n21869), .B(n22153), .Z(n21873) );
  XOR U6485 ( .A(n21314), .B(n21598), .Z(n21318) );
  XOR U6486 ( .A(n20752), .B(n21036), .Z(n20756) );
  XOR U6487 ( .A(n20185), .B(n20469), .Z(n20189) );
  XOR U6488 ( .A(n19612), .B(n19896), .Z(n19616) );
  XOR U6489 ( .A(n19033), .B(n19317), .Z(n19037) );
  XOR U6490 ( .A(n12555), .B(n13134), .Z(n12559) );
  XOR U6491 ( .A(n11967), .B(n12476), .Z(n11971) );
  XOR U6492 ( .A(n17727), .B(n18042), .Z(n17731) );
  XOR U6493 ( .A(n16505), .B(n16844), .Z(n16509) );
  XOR U6494 ( .A(n15259), .B(n15622), .Z(n15263) );
  XOR U6495 ( .A(n15840), .B(n16245), .Z(n15844) );
  XOR U6496 ( .A(n14582), .B(n15011), .Z(n14586) );
  XOR U6497 ( .A(n13300), .B(n13753), .Z(n13304) );
  XOR U6498 ( .A(n13899), .B(n14394), .Z(n13903) );
  XOR U6499 ( .A(n12605), .B(n13124), .Z(n12609) );
  XOR U6500 ( .A(n11240), .B(n11837), .Z(n11244) );
  XOR U6501 ( .A(n9898), .B(n10519), .Z(n9902) );
  XOR U6502 ( .A(n10552), .B(n11185), .Z(n10556) );
  XOR U6503 ( .A(n17752), .B(n18037), .Z(n17756) );
  XOR U6504 ( .A(n11997), .B(n12470), .Z(n12001) );
  XOR U6505 ( .A(n9203), .B(n9854), .Z(n9207) );
  XOR U6506 ( .A(n7825), .B(n8500), .Z(n7829) );
  XOR U6507 ( .A(n11932), .B(n12483), .Z(n11936) );
  XOR U6508 ( .A(n10602), .B(n11175), .Z(n10606) );
  XOR U6509 ( .A(n13929), .B(n14388), .Z(n13933) );
  XOR U6510 ( .A(n12635), .B(n13118), .Z(n12639) );
  XOR U6511 ( .A(n15870), .B(n16239), .Z(n15874) );
  XOR U6512 ( .A(n14612), .B(n15005), .Z(n14616) );
  XOR U6513 ( .A(n13330), .B(n13747), .Z(n13334) );
  XOR U6514 ( .A(n16535), .B(n16838), .Z(n16539) );
  XOR U6515 ( .A(n15289), .B(n15616), .Z(n15293) );
  XOR U6516 ( .A(n41211), .B(n41477), .Z(n41215) );
  XOR U6517 ( .A(n40938), .B(n41204), .Z(n40942) );
  XOR U6518 ( .A(n40659), .B(n40925), .Z(n40663) );
  XOR U6519 ( .A(n40374), .B(n40640), .Z(n40378) );
  XOR U6520 ( .A(n40083), .B(n40349), .Z(n40087) );
  XOR U6521 ( .A(n39483), .B(n39749), .Z(n39487) );
  XOR U6522 ( .A(n39174), .B(n39440), .Z(n39178) );
  XOR U6523 ( .A(n38859), .B(n39125), .Z(n38863) );
  XOR U6524 ( .A(n38538), .B(n38804), .Z(n38542) );
  XOR U6525 ( .A(n38211), .B(n38477), .Z(n38215) );
  XOR U6526 ( .A(n37878), .B(n38144), .Z(n37882) );
  XOR U6527 ( .A(n37539), .B(n37805), .Z(n37543) );
  XOR U6528 ( .A(n37194), .B(n37460), .Z(n37198) );
  XOR U6529 ( .A(n36843), .B(n37109), .Z(n36847) );
  XOR U6530 ( .A(n36486), .B(n36752), .Z(n36490) );
  XOR U6531 ( .A(n36123), .B(n36389), .Z(n36127) );
  XOR U6532 ( .A(n35754), .B(n36020), .Z(n35758) );
  XOR U6533 ( .A(n35379), .B(n35645), .Z(n35383) );
  XOR U6534 ( .A(n34998), .B(n35264), .Z(n35002) );
  XOR U6535 ( .A(n34611), .B(n34877), .Z(n34615) );
  XOR U6536 ( .A(n34218), .B(n34484), .Z(n34222) );
  XOR U6537 ( .A(n33819), .B(n34085), .Z(n33823) );
  XOR U6538 ( .A(n33414), .B(n33680), .Z(n33418) );
  XOR U6539 ( .A(n33003), .B(n33269), .Z(n33007) );
  XOR U6540 ( .A(n32586), .B(n32852), .Z(n32590) );
  XOR U6541 ( .A(n32163), .B(n32429), .Z(n32167) );
  XOR U6542 ( .A(n31734), .B(n32000), .Z(n31738) );
  XOR U6543 ( .A(n31299), .B(n31565), .Z(n31303) );
  XOR U6544 ( .A(n30858), .B(n31124), .Z(n30862) );
  XOR U6545 ( .A(n30411), .B(n30677), .Z(n30415) );
  XOR U6546 ( .A(n29958), .B(n30224), .Z(n29962) );
  XOR U6547 ( .A(n29499), .B(n29765), .Z(n29503) );
  XOR U6548 ( .A(n29034), .B(n29300), .Z(n29038) );
  XOR U6549 ( .A(n28563), .B(n28829), .Z(n28567) );
  XOR U6550 ( .A(n28086), .B(n28352), .Z(n28090) );
  XOR U6551 ( .A(n27603), .B(n27869), .Z(n27607) );
  XOR U6552 ( .A(n27114), .B(n27380), .Z(n27118) );
  XOR U6553 ( .A(n26617), .B(n26883), .Z(n26621) );
  XOR U6554 ( .A(n26116), .B(n26382), .Z(n26120) );
  XOR U6555 ( .A(n25608), .B(n25874), .Z(n25612) );
  XOR U6556 ( .A(n25094), .B(n25360), .Z(n25098) );
  XOR U6557 ( .A(n24571), .B(n24837), .Z(n24575) );
  XOR U6558 ( .A(n24046), .B(n24312), .Z(n24050) );
  XOR U6559 ( .A(n23515), .B(n23781), .Z(n23519) );
  XOR U6560 ( .A(n22977), .B(n23243), .Z(n22981) );
  XOR U6561 ( .A(n22433), .B(n22699), .Z(n22437) );
  XOR U6562 ( .A(n21884), .B(n22150), .Z(n21888) );
  XOR U6563 ( .A(n21329), .B(n21595), .Z(n21333) );
  XOR U6564 ( .A(n20767), .B(n21033), .Z(n20771) );
  XOR U6565 ( .A(n20200), .B(n20466), .Z(n20204) );
  XOR U6566 ( .A(n19627), .B(n19893), .Z(n19631) );
  XOR U6567 ( .A(n19048), .B(n19314), .Z(n19052) );
  XOR U6568 ( .A(n17767), .B(n18034), .Z(n17771) );
  XOR U6569 ( .A(n16560), .B(n16833), .Z(n16564) );
  XOR U6570 ( .A(n10627), .B(n11170), .Z(n10631) );
  XOR U6571 ( .A(n6428), .B(n7121), .Z(n6432) );
  XOR U6572 ( .A(n12027), .B(n12464), .Z(n12031) );
  XOR U6573 ( .A(n15319), .B(n15610), .Z(n15323) );
  XOR U6574 ( .A(n15900), .B(n16233), .Z(n15904) );
  XOR U6575 ( .A(n14642), .B(n14999), .Z(n14646) );
  XOR U6576 ( .A(n13360), .B(n13741), .Z(n13364) );
  XOR U6577 ( .A(n13959), .B(n14382), .Z(n13963) );
  XOR U6578 ( .A(n12665), .B(n13112), .Z(n12669) );
  XOR U6579 ( .A(n11300), .B(n11825), .Z(n11304) );
  XOR U6580 ( .A(n9913), .B(n10516), .Z(n9917) );
  XOR U6581 ( .A(n7157), .B(n7808), .Z(n7161) );
  XOR U6582 ( .A(n8572), .B(n9169), .Z(n8576) );
  XOR U6583 ( .A(n10657), .B(n11164), .Z(n10661) );
  XOR U6584 ( .A(n17179), .B(n17434), .Z(n17183) );
  XOR U6585 ( .A(n12057), .B(n12458), .Z(n12061) );
  XOR U6586 ( .A(n7860), .B(n8493), .Z(n7864) );
  XOR U6587 ( .A(n7840), .B(n8497), .Z(n7844) );
  XOR U6588 ( .A(n9943), .B(n10510), .Z(n9947) );
  XOR U6589 ( .A(n11330), .B(n11819), .Z(n11334) );
  XOR U6590 ( .A(n13989), .B(n14376), .Z(n13993) );
  XOR U6591 ( .A(n12695), .B(n13106), .Z(n12699) );
  XOR U6592 ( .A(n15930), .B(n16227), .Z(n15934) );
  XOR U6593 ( .A(n14672), .B(n14993), .Z(n14676) );
  XOR U6594 ( .A(n13390), .B(n13735), .Z(n13394) );
  XOR U6595 ( .A(n15349), .B(n15604), .Z(n15353) );
  XOR U6596 ( .A(n42009), .B(n42257), .Z(n42013) );
  XOR U6597 ( .A(n41754), .B(n42002), .Z(n41758) );
  XOR U6598 ( .A(n41493), .B(n41741), .Z(n41497) );
  XOR U6599 ( .A(n41226), .B(n41474), .Z(n41230) );
  XOR U6600 ( .A(n40953), .B(n41201), .Z(n40957) );
  XOR U6601 ( .A(n40389), .B(n40637), .Z(n40393) );
  XOR U6602 ( .A(n40098), .B(n40346), .Z(n40102) );
  XOR U6603 ( .A(n39801), .B(n40049), .Z(n39805) );
  XOR U6604 ( .A(n39498), .B(n39746), .Z(n39502) );
  XOR U6605 ( .A(n39189), .B(n39437), .Z(n39193) );
  XOR U6606 ( .A(n38874), .B(n39122), .Z(n38878) );
  XOR U6607 ( .A(n38553), .B(n38801), .Z(n38557) );
  XOR U6608 ( .A(n38226), .B(n38474), .Z(n38230) );
  XOR U6609 ( .A(n37893), .B(n38141), .Z(n37897) );
  XOR U6610 ( .A(n37554), .B(n37802), .Z(n37558) );
  XOR U6611 ( .A(n37209), .B(n37457), .Z(n37213) );
  XOR U6612 ( .A(n36858), .B(n37106), .Z(n36862) );
  XOR U6613 ( .A(n36501), .B(n36749), .Z(n36505) );
  XOR U6614 ( .A(n36138), .B(n36386), .Z(n36142) );
  XOR U6615 ( .A(n35769), .B(n36017), .Z(n35773) );
  XOR U6616 ( .A(n35394), .B(n35642), .Z(n35398) );
  XOR U6617 ( .A(n35013), .B(n35261), .Z(n35017) );
  XOR U6618 ( .A(n34626), .B(n34874), .Z(n34630) );
  XOR U6619 ( .A(n34233), .B(n34481), .Z(n34237) );
  XOR U6620 ( .A(n33834), .B(n34082), .Z(n33838) );
  XOR U6621 ( .A(n33429), .B(n33677), .Z(n33433) );
  XOR U6622 ( .A(n33018), .B(n33266), .Z(n33022) );
  XOR U6623 ( .A(n32601), .B(n32849), .Z(n32605) );
  XOR U6624 ( .A(n32178), .B(n32426), .Z(n32182) );
  XOR U6625 ( .A(n31749), .B(n31997), .Z(n31753) );
  XOR U6626 ( .A(n31314), .B(n31562), .Z(n31318) );
  XOR U6627 ( .A(n30873), .B(n31121), .Z(n30877) );
  XOR U6628 ( .A(n30426), .B(n30674), .Z(n30430) );
  XOR U6629 ( .A(n29973), .B(n30221), .Z(n29977) );
  XOR U6630 ( .A(n29514), .B(n29762), .Z(n29518) );
  XOR U6631 ( .A(n29049), .B(n29297), .Z(n29053) );
  XOR U6632 ( .A(n28578), .B(n28826), .Z(n28582) );
  XOR U6633 ( .A(n28101), .B(n28349), .Z(n28105) );
  XOR U6634 ( .A(n27618), .B(n27866), .Z(n27622) );
  XOR U6635 ( .A(n27129), .B(n27377), .Z(n27133) );
  XOR U6636 ( .A(n26632), .B(n26880), .Z(n26636) );
  XOR U6637 ( .A(n26131), .B(n26379), .Z(n26135) );
  XOR U6638 ( .A(n25623), .B(n25871), .Z(n25627) );
  XOR U6639 ( .A(n25109), .B(n25357), .Z(n25113) );
  XOR U6640 ( .A(n24586), .B(n24834), .Z(n24590) );
  XOR U6641 ( .A(n24061), .B(n24309), .Z(n24065) );
  XOR U6642 ( .A(n23530), .B(n23778), .Z(n23534) );
  XOR U6643 ( .A(n22992), .B(n23240), .Z(n22996) );
  XOR U6644 ( .A(n22448), .B(n22696), .Z(n22452) );
  XOR U6645 ( .A(n21899), .B(n22147), .Z(n21903) );
  XOR U6646 ( .A(n21344), .B(n21592), .Z(n21348) );
  XOR U6647 ( .A(n20782), .B(n21030), .Z(n20786) );
  XOR U6648 ( .A(n20215), .B(n20463), .Z(n20219) );
  XOR U6649 ( .A(n19642), .B(n19890), .Z(n19646) );
  XOR U6650 ( .A(n19063), .B(n19311), .Z(n19067) );
  XOR U6651 ( .A(n18374), .B(n18669), .Z(n18378) );
  XOR U6652 ( .A(n10687), .B(n11158), .Z(n10691) );
  XOR U6653 ( .A(n9288), .B(n9837), .Z(n9292) );
  XOR U6654 ( .A(n7910), .B(n8483), .Z(n7914) );
  XOR U6655 ( .A(n6443), .B(n7118), .Z(n6447) );
  XOR U6656 ( .A(n5015), .B(n5716), .Z(n5019) );
  XOR U6657 ( .A(n12087), .B(n12452), .Z(n12091) );
  XOR U6658 ( .A(n15960), .B(n16221), .Z(n15964) );
  XOR U6659 ( .A(n14702), .B(n14987), .Z(n14706) );
  XOR U6660 ( .A(n13420), .B(n13729), .Z(n13424) );
  XOR U6661 ( .A(n14019), .B(n14370), .Z(n14023) );
  XOR U6662 ( .A(n12725), .B(n13100), .Z(n12729) );
  XOR U6663 ( .A(n11360), .B(n11813), .Z(n11364) );
  XOR U6664 ( .A(n9973), .B(n10504), .Z(n9977) );
  XOR U6665 ( .A(n5758), .B(n6415), .Z(n5762) );
  XOR U6666 ( .A(n7895), .B(n8486), .Z(n7899) );
  XOR U6667 ( .A(n6493), .B(n7108), .Z(n6497) );
  XOR U6668 ( .A(n9318), .B(n9831), .Z(n9322) );
  XOR U6669 ( .A(n7940), .B(n8477), .Z(n7944) );
  XOR U6670 ( .A(n10717), .B(n11152), .Z(n10721) );
  XOR U6671 ( .A(n12117), .B(n12446), .Z(n12121) );
  XOR U6672 ( .A(n7177), .B(n7804), .Z(n7181) );
  XOR U6673 ( .A(n5070), .B(n5705), .Z(n5074) );
  XOR U6674 ( .A(n10003), .B(n10498), .Z(n10007) );
  XOR U6675 ( .A(n11390), .B(n11807), .Z(n11394) );
  XOR U6676 ( .A(n14049), .B(n14364), .Z(n14053) );
  XOR U6677 ( .A(n12755), .B(n13094), .Z(n12759) );
  XOR U6678 ( .A(n14732), .B(n14981), .Z(n14736) );
  XOR U6679 ( .A(n13450), .B(n13723), .Z(n13454) );
  XOR U6680 ( .A(n42753), .B(n42983), .Z(n42757) );
  XOR U6681 ( .A(n42516), .B(n42746), .Z(n42520) );
  XOR U6682 ( .A(n42273), .B(n42503), .Z(n42277) );
  XOR U6683 ( .A(n42024), .B(n42254), .Z(n42028) );
  XOR U6684 ( .A(n41769), .B(n41999), .Z(n41773) );
  XOR U6685 ( .A(n41241), .B(n41471), .Z(n41245) );
  XOR U6686 ( .A(n40968), .B(n41198), .Z(n40972) );
  XOR U6687 ( .A(n40689), .B(n40919), .Z(n40693) );
  XOR U6688 ( .A(n40404), .B(n40634), .Z(n40408) );
  XOR U6689 ( .A(n40113), .B(n40343), .Z(n40117) );
  XOR U6690 ( .A(n39816), .B(n40046), .Z(n39820) );
  XOR U6691 ( .A(n39513), .B(n39743), .Z(n39517) );
  XOR U6692 ( .A(n39204), .B(n39434), .Z(n39208) );
  XOR U6693 ( .A(n38889), .B(n39119), .Z(n38893) );
  XOR U6694 ( .A(n38568), .B(n38798), .Z(n38572) );
  XOR U6695 ( .A(n38241), .B(n38471), .Z(n38245) );
  XOR U6696 ( .A(n37908), .B(n38138), .Z(n37912) );
  XOR U6697 ( .A(n37569), .B(n37799), .Z(n37573) );
  XOR U6698 ( .A(n37224), .B(n37454), .Z(n37228) );
  XOR U6699 ( .A(n36873), .B(n37103), .Z(n36877) );
  XOR U6700 ( .A(n36516), .B(n36746), .Z(n36520) );
  XOR U6701 ( .A(n36153), .B(n36383), .Z(n36157) );
  XOR U6702 ( .A(n35784), .B(n36014), .Z(n35788) );
  XOR U6703 ( .A(n35409), .B(n35639), .Z(n35413) );
  XOR U6704 ( .A(n35028), .B(n35258), .Z(n35032) );
  XOR U6705 ( .A(n34641), .B(n34871), .Z(n34645) );
  XOR U6706 ( .A(n34248), .B(n34478), .Z(n34252) );
  XOR U6707 ( .A(n33849), .B(n34079), .Z(n33853) );
  XOR U6708 ( .A(n33444), .B(n33674), .Z(n33448) );
  XOR U6709 ( .A(n33033), .B(n33263), .Z(n33037) );
  XOR U6710 ( .A(n32616), .B(n32846), .Z(n32620) );
  XOR U6711 ( .A(n32193), .B(n32423), .Z(n32197) );
  XOR U6712 ( .A(n31764), .B(n31994), .Z(n31768) );
  XOR U6713 ( .A(n31329), .B(n31559), .Z(n31333) );
  XOR U6714 ( .A(n30888), .B(n31118), .Z(n30892) );
  XOR U6715 ( .A(n30441), .B(n30671), .Z(n30445) );
  XOR U6716 ( .A(n29988), .B(n30218), .Z(n29992) );
  XOR U6717 ( .A(n29529), .B(n29759), .Z(n29533) );
  XOR U6718 ( .A(n29064), .B(n29294), .Z(n29068) );
  XOR U6719 ( .A(n28593), .B(n28823), .Z(n28597) );
  XOR U6720 ( .A(n28116), .B(n28346), .Z(n28120) );
  XOR U6721 ( .A(n27633), .B(n27863), .Z(n27637) );
  XOR U6722 ( .A(n27144), .B(n27374), .Z(n27148) );
  XOR U6723 ( .A(n26647), .B(n26877), .Z(n26651) );
  XOR U6724 ( .A(n26146), .B(n26376), .Z(n26150) );
  XOR U6725 ( .A(n25638), .B(n25868), .Z(n25642) );
  XOR U6726 ( .A(n25124), .B(n25354), .Z(n25128) );
  XOR U6727 ( .A(n24601), .B(n24831), .Z(n24605) );
  XOR U6728 ( .A(n24076), .B(n24306), .Z(n24080) );
  XOR U6729 ( .A(n23545), .B(n23775), .Z(n23549) );
  XOR U6730 ( .A(n23007), .B(n23237), .Z(n23011) );
  XOR U6731 ( .A(n22463), .B(n22693), .Z(n22467) );
  XOR U6732 ( .A(n21914), .B(n22144), .Z(n21918) );
  XOR U6733 ( .A(n21359), .B(n21589), .Z(n21363) );
  XOR U6734 ( .A(n20797), .B(n21027), .Z(n20801) );
  XOR U6735 ( .A(n20230), .B(n20460), .Z(n20234) );
  XOR U6736 ( .A(n19657), .B(n19887), .Z(n19661) );
  XOR U6737 ( .A(n19078), .B(n19308), .Z(n19082) );
  XOR U6738 ( .A(n17797), .B(n18028), .Z(n17801) );
  XOR U6739 ( .A(n16595), .B(n16826), .Z(n16599) );
  XOR U6740 ( .A(n10747), .B(n11146), .Z(n10751) );
  XOR U6741 ( .A(n9348), .B(n9825), .Z(n9352) );
  XOR U6742 ( .A(n7970), .B(n8471), .Z(n7974) );
  XOR U6743 ( .A(n7925), .B(n8480), .Z(n7929) );
  XOR U6744 ( .A(n6523), .B(n7102), .Z(n6527) );
  XOR U6745 ( .A(n3600), .B(n4281), .Z(n3604) );
  XOR U6746 ( .A(n5030), .B(n5713), .Z(n5034) );
  XOR U6747 ( .A(n2106), .B(n2835), .Z(n2110) );
  XOR U6748 ( .A(n12147), .B(n12440), .Z(n12151) );
  XOR U6749 ( .A(n13480), .B(n13717), .Z(n13484) );
  XOR U6750 ( .A(n14079), .B(n14358), .Z(n14083) );
  XOR U6751 ( .A(n12785), .B(n13088), .Z(n12789) );
  XOR U6752 ( .A(n11420), .B(n11801), .Z(n11424) );
  XOR U6753 ( .A(n10033), .B(n10492), .Z(n10037) );
  XOR U6754 ( .A(n5100), .B(n5699), .Z(n5104) );
  XOR U6755 ( .A(n5055), .B(n5708), .Z(n5059) );
  XOR U6756 ( .A(n3585), .B(n4284), .Z(n3589) );
  XOR U6757 ( .A(n6508), .B(n7105), .Z(n6512) );
  XOR U6758 ( .A(n7955), .B(n8474), .Z(n7959) );
  XOR U6759 ( .A(n6553), .B(n7096), .Z(n6557) );
  XOR U6760 ( .A(n9378), .B(n9819), .Z(n9382) );
  XOR U6761 ( .A(n8000), .B(n8465), .Z(n8004) );
  XOR U6762 ( .A(n10777), .B(n11140), .Z(n10781) );
  XOR U6763 ( .A(n14757), .B(n14976), .Z(n14761) );
  XOR U6764 ( .A(n12177), .B(n12434), .Z(n12181) );
  XOR U6765 ( .A(n5085), .B(n5702), .Z(n5089) );
  XOR U6766 ( .A(n5130), .B(n5693), .Z(n5134) );
  XOR U6767 ( .A(n10063), .B(n10486), .Z(n10067) );
  XOR U6768 ( .A(n11450), .B(n11795), .Z(n11454) );
  XOR U6769 ( .A(n14109), .B(n14352), .Z(n14113) );
  XOR U6770 ( .A(n12815), .B(n13082), .Z(n12819) );
  XOR U6771 ( .A(n43443), .B(n43655), .Z(n43447) );
  XOR U6772 ( .A(n43224), .B(n43436), .Z(n43228) );
  XOR U6773 ( .A(n42999), .B(n43211), .Z(n43003) );
  XOR U6774 ( .A(n42768), .B(n42980), .Z(n42772) );
  XOR U6775 ( .A(n42531), .B(n42743), .Z(n42535) );
  XOR U6776 ( .A(n42039), .B(n42251), .Z(n42043) );
  XOR U6777 ( .A(n41784), .B(n41996), .Z(n41788) );
  XOR U6778 ( .A(n41523), .B(n41735), .Z(n41527) );
  XOR U6779 ( .A(n41256), .B(n41468), .Z(n41260) );
  XOR U6780 ( .A(n40983), .B(n41195), .Z(n40987) );
  XOR U6781 ( .A(n40704), .B(n40916), .Z(n40708) );
  XOR U6782 ( .A(n40419), .B(n40631), .Z(n40423) );
  XOR U6783 ( .A(n40128), .B(n40340), .Z(n40132) );
  XOR U6784 ( .A(n39831), .B(n40043), .Z(n39835) );
  XOR U6785 ( .A(n39528), .B(n39740), .Z(n39532) );
  XOR U6786 ( .A(n39219), .B(n39431), .Z(n39223) );
  XOR U6787 ( .A(n38904), .B(n39116), .Z(n38908) );
  XOR U6788 ( .A(n38583), .B(n38795), .Z(n38587) );
  XOR U6789 ( .A(n38256), .B(n38468), .Z(n38260) );
  XOR U6790 ( .A(n37923), .B(n38135), .Z(n37927) );
  XOR U6791 ( .A(n37584), .B(n37796), .Z(n37588) );
  XOR U6792 ( .A(n37239), .B(n37451), .Z(n37243) );
  XOR U6793 ( .A(n36888), .B(n37100), .Z(n36892) );
  XOR U6794 ( .A(n36531), .B(n36743), .Z(n36535) );
  XOR U6795 ( .A(n36168), .B(n36380), .Z(n36172) );
  XOR U6796 ( .A(n35799), .B(n36011), .Z(n35803) );
  XOR U6797 ( .A(n35424), .B(n35636), .Z(n35428) );
  XOR U6798 ( .A(n35043), .B(n35255), .Z(n35047) );
  XOR U6799 ( .A(n34656), .B(n34868), .Z(n34660) );
  XOR U6800 ( .A(n34263), .B(n34475), .Z(n34267) );
  XOR U6801 ( .A(n33864), .B(n34076), .Z(n33868) );
  XOR U6802 ( .A(n33459), .B(n33671), .Z(n33463) );
  XOR U6803 ( .A(n33048), .B(n33260), .Z(n33052) );
  XOR U6804 ( .A(n32631), .B(n32843), .Z(n32635) );
  XOR U6805 ( .A(n32208), .B(n32420), .Z(n32212) );
  XOR U6806 ( .A(n31779), .B(n31991), .Z(n31783) );
  XOR U6807 ( .A(n31344), .B(n31556), .Z(n31348) );
  XOR U6808 ( .A(n30903), .B(n31115), .Z(n30907) );
  XOR U6809 ( .A(n30456), .B(n30668), .Z(n30460) );
  XOR U6810 ( .A(n30003), .B(n30215), .Z(n30007) );
  XOR U6811 ( .A(n29544), .B(n29756), .Z(n29548) );
  XOR U6812 ( .A(n29079), .B(n29291), .Z(n29083) );
  XOR U6813 ( .A(n28608), .B(n28820), .Z(n28612) );
  XOR U6814 ( .A(n28131), .B(n28343), .Z(n28135) );
  XOR U6815 ( .A(n27648), .B(n27860), .Z(n27652) );
  XOR U6816 ( .A(n27159), .B(n27371), .Z(n27163) );
  XOR U6817 ( .A(n26662), .B(n26874), .Z(n26666) );
  XOR U6818 ( .A(n26161), .B(n26373), .Z(n26165) );
  XOR U6819 ( .A(n25653), .B(n25865), .Z(n25657) );
  XOR U6820 ( .A(n25139), .B(n25351), .Z(n25143) );
  XOR U6821 ( .A(n24616), .B(n24828), .Z(n24620) );
  XOR U6822 ( .A(n24091), .B(n24303), .Z(n24095) );
  XOR U6823 ( .A(n23560), .B(n23772), .Z(n23564) );
  XOR U6824 ( .A(n23022), .B(n23234), .Z(n23026) );
  XOR U6825 ( .A(n22478), .B(n22690), .Z(n22482) );
  XOR U6826 ( .A(n21929), .B(n22141), .Z(n21933) );
  XOR U6827 ( .A(n21374), .B(n21586), .Z(n21378) );
  XOR U6828 ( .A(n20812), .B(n21024), .Z(n20816) );
  XOR U6829 ( .A(n20245), .B(n20457), .Z(n20249) );
  XOR U6830 ( .A(n19672), .B(n19884), .Z(n19676) );
  XOR U6831 ( .A(n19093), .B(n19305), .Z(n19097) );
  XOR U6832 ( .A(n18404), .B(n18657), .Z(n18408) );
  XOR U6833 ( .A(n17214), .B(n17427), .Z(n17218) );
  XOR U6834 ( .A(n16000), .B(n16213), .Z(n16004) );
  XOR U6835 ( .A(n14134), .B(n14347), .Z(n14138) );
  XOR U6836 ( .A(n10807), .B(n11134), .Z(n10811) );
  XOR U6837 ( .A(n9408), .B(n9813), .Z(n9412) );
  XOR U6838 ( .A(n8030), .B(n8459), .Z(n8034) );
  XOR U6839 ( .A(n7985), .B(n8468), .Z(n7989) );
  XOR U6840 ( .A(n6583), .B(n7090), .Z(n6587) );
  XOR U6841 ( .A(n6538), .B(n7099), .Z(n6542) );
  XOR U6842 ( .A(n2881), .B(n3556), .Z(n2885) );
  XOR U6843 ( .A(n1395), .B(n2094), .Z(n1399) );
  XOR U6844 ( .A(n1375), .B(n2098), .Z(n1379) );
  XOR U6845 ( .A(n12207), .B(n12428), .Z(n12211) );
  XOR U6846 ( .A(n12845), .B(n13076), .Z(n12849) );
  XOR U6847 ( .A(n11480), .B(n11789), .Z(n11484) );
  XOR U6848 ( .A(n10093), .B(n10480), .Z(n10097) );
  XOR U6849 ( .A(n5160), .B(n5687), .Z(n5164) );
  XOR U6850 ( .A(n5115), .B(n5696), .Z(n5119) );
  XOR U6851 ( .A(n3620), .B(n4277), .Z(n3624) );
  XOR U6852 ( .A(n2126), .B(n2831), .Z(n2130) );
  XOR U6853 ( .A(n2911), .B(n3550), .Z(n2915) );
  XOR U6854 ( .A(n1425), .B(n2088), .Z(n1429) );
  XOR U6855 ( .A(n6568), .B(n7093), .Z(n6572) );
  XOR U6856 ( .A(n8015), .B(n8462), .Z(n8019) );
  XOR U6857 ( .A(n6613), .B(n7084), .Z(n6617) );
  XOR U6858 ( .A(n9438), .B(n9807), .Z(n9442) );
  XOR U6859 ( .A(n8060), .B(n8453), .Z(n8064) );
  XOR U6860 ( .A(n10837), .B(n11128), .Z(n10841) );
  XOR U6861 ( .A(n3650), .B(n4271), .Z(n3654) );
  XOR U6862 ( .A(n5145), .B(n5690), .Z(n5149) );
  XOR U6863 ( .A(n5190), .B(n5681), .Z(n5194) );
  XOR U6864 ( .A(n10123), .B(n10474), .Z(n10127) );
  XOR U6865 ( .A(n11510), .B(n11783), .Z(n11514) );
  XOR U6866 ( .A(n44079), .B(n44273), .Z(n44083) );
  XOR U6867 ( .A(n43878), .B(n44072), .Z(n43882) );
  XOR U6868 ( .A(n43671), .B(n43865), .Z(n43675) );
  XOR U6869 ( .A(n43458), .B(n43652), .Z(n43462) );
  XOR U6870 ( .A(n43239), .B(n43433), .Z(n43243) );
  XOR U6871 ( .A(n42783), .B(n42977), .Z(n42787) );
  XOR U6872 ( .A(n42546), .B(n42740), .Z(n42550) );
  XOR U6873 ( .A(n42303), .B(n42497), .Z(n42307) );
  XOR U6874 ( .A(n42054), .B(n42248), .Z(n42058) );
  XOR U6875 ( .A(n41799), .B(n41993), .Z(n41803) );
  XOR U6876 ( .A(n41538), .B(n41732), .Z(n41542) );
  XOR U6877 ( .A(n41271), .B(n41465), .Z(n41275) );
  XOR U6878 ( .A(n40998), .B(n41192), .Z(n41002) );
  XOR U6879 ( .A(n40719), .B(n40913), .Z(n40723) );
  XOR U6880 ( .A(n40434), .B(n40628), .Z(n40438) );
  XOR U6881 ( .A(n40143), .B(n40337), .Z(n40147) );
  XOR U6882 ( .A(n39846), .B(n40040), .Z(n39850) );
  XOR U6883 ( .A(n39543), .B(n39737), .Z(n39547) );
  XOR U6884 ( .A(n39234), .B(n39428), .Z(n39238) );
  XOR U6885 ( .A(n38919), .B(n39113), .Z(n38923) );
  XOR U6886 ( .A(n38598), .B(n38792), .Z(n38602) );
  XOR U6887 ( .A(n38271), .B(n38465), .Z(n38275) );
  XOR U6888 ( .A(n37938), .B(n38132), .Z(n37942) );
  XOR U6889 ( .A(n37599), .B(n37793), .Z(n37603) );
  XOR U6890 ( .A(n37254), .B(n37448), .Z(n37258) );
  XOR U6891 ( .A(n36903), .B(n37097), .Z(n36907) );
  XOR U6892 ( .A(n36546), .B(n36740), .Z(n36550) );
  XOR U6893 ( .A(n36183), .B(n36377), .Z(n36187) );
  XOR U6894 ( .A(n35814), .B(n36008), .Z(n35818) );
  XOR U6895 ( .A(n35439), .B(n35633), .Z(n35443) );
  XOR U6896 ( .A(n35058), .B(n35252), .Z(n35062) );
  XOR U6897 ( .A(n34671), .B(n34865), .Z(n34675) );
  XOR U6898 ( .A(n34278), .B(n34472), .Z(n34282) );
  XOR U6899 ( .A(n33879), .B(n34073), .Z(n33883) );
  XOR U6900 ( .A(n33474), .B(n33668), .Z(n33478) );
  XOR U6901 ( .A(n33063), .B(n33257), .Z(n33067) );
  XOR U6902 ( .A(n32646), .B(n32840), .Z(n32650) );
  XOR U6903 ( .A(n32223), .B(n32417), .Z(n32227) );
  XOR U6904 ( .A(n31794), .B(n31988), .Z(n31798) );
  XOR U6905 ( .A(n31359), .B(n31553), .Z(n31363) );
  XOR U6906 ( .A(n30918), .B(n31112), .Z(n30922) );
  XOR U6907 ( .A(n30471), .B(n30665), .Z(n30475) );
  XOR U6908 ( .A(n30018), .B(n30212), .Z(n30022) );
  XOR U6909 ( .A(n29559), .B(n29753), .Z(n29563) );
  XOR U6910 ( .A(n29094), .B(n29288), .Z(n29098) );
  XOR U6911 ( .A(n28623), .B(n28817), .Z(n28627) );
  XOR U6912 ( .A(n28146), .B(n28340), .Z(n28150) );
  XOR U6913 ( .A(n27663), .B(n27857), .Z(n27667) );
  XOR U6914 ( .A(n27174), .B(n27368), .Z(n27178) );
  XOR U6915 ( .A(n26677), .B(n26871), .Z(n26681) );
  XOR U6916 ( .A(n26176), .B(n26370), .Z(n26180) );
  XOR U6917 ( .A(n25668), .B(n25862), .Z(n25672) );
  XOR U6918 ( .A(n25154), .B(n25348), .Z(n25158) );
  XOR U6919 ( .A(n24631), .B(n24825), .Z(n24635) );
  XOR U6920 ( .A(n24106), .B(n24300), .Z(n24110) );
  XOR U6921 ( .A(n23575), .B(n23769), .Z(n23579) );
  XOR U6922 ( .A(n23037), .B(n23231), .Z(n23041) );
  XOR U6923 ( .A(n22493), .B(n22687), .Z(n22497) );
  XOR U6924 ( .A(n21944), .B(n22138), .Z(n21948) );
  XOR U6925 ( .A(n21389), .B(n21583), .Z(n21393) );
  XOR U6926 ( .A(n20827), .B(n21021), .Z(n20831) );
  XOR U6927 ( .A(n20260), .B(n20454), .Z(n20264) );
  XOR U6928 ( .A(n19687), .B(n19881), .Z(n19691) );
  XOR U6929 ( .A(n19108), .B(n19302), .Z(n19112) );
  XOR U6930 ( .A(n17827), .B(n18022), .Z(n17831) );
  XOR U6931 ( .A(n16625), .B(n16820), .Z(n16629) );
  XOR U6932 ( .A(n15399), .B(n15594), .Z(n15403) );
  XOR U6933 ( .A(n14149), .B(n14344), .Z(n14153) );
  XOR U6934 ( .A(n12875), .B(n13070), .Z(n12879) );
  XOR U6935 ( .A(n10867), .B(n11122), .Z(n10871) );
  XOR U6936 ( .A(n9468), .B(n9801), .Z(n9472) );
  XOR U6937 ( .A(n8090), .B(n8447), .Z(n8094) );
  XOR U6938 ( .A(n8045), .B(n8456), .Z(n8049) );
  XOR U6939 ( .A(n6643), .B(n7078), .Z(n6647) );
  XOR U6940 ( .A(n6598), .B(n7087), .Z(n6602) );
  XOR U6941 ( .A(n2941), .B(n3544), .Z(n2945) );
  XOR U6942 ( .A(n1455), .B(n2082), .Z(n1459) );
  XOR U6943 ( .A(n1410), .B(n2091), .Z(n1414) );
  XOR U6944 ( .A(n11540), .B(n11777), .Z(n11544) );
  XOR U6945 ( .A(n10153), .B(n10468), .Z(n10157) );
  XOR U6946 ( .A(n5220), .B(n5675), .Z(n5224) );
  XOR U6947 ( .A(n5175), .B(n5684), .Z(n5179) );
  XOR U6948 ( .A(n3680), .B(n4265), .Z(n3684) );
  XOR U6949 ( .A(n1440), .B(n2085), .Z(n1444) );
  XOR U6950 ( .A(n2971), .B(n3538), .Z(n2975) );
  XOR U6951 ( .A(n1485), .B(n2076), .Z(n1489) );
  XOR U6952 ( .A(n6628), .B(n7081), .Z(n6632) );
  XOR U6953 ( .A(n8075), .B(n8450), .Z(n8079) );
  XOR U6954 ( .A(n6673), .B(n7072), .Z(n6677) );
  XOR U6955 ( .A(n9498), .B(n9795), .Z(n9502) );
  XOR U6956 ( .A(n8120), .B(n8441), .Z(n8124) );
  XOR U6957 ( .A(n10897), .B(n11116), .Z(n10901) );
  XOR U6958 ( .A(n3710), .B(n4259), .Z(n3714) );
  XOR U6959 ( .A(n5205), .B(n5678), .Z(n5209) );
  XOR U6960 ( .A(n5250), .B(n5669), .Z(n5254) );
  XOR U6961 ( .A(n10183), .B(n10462), .Z(n10187) );
  XOR U6962 ( .A(n11570), .B(n11771), .Z(n11574) );
  XOR U6963 ( .A(n44661), .B(n44837), .Z(n44665) );
  XOR U6964 ( .A(n44478), .B(n44654), .Z(n44482) );
  XOR U6965 ( .A(n44289), .B(n44465), .Z(n44293) );
  XOR U6966 ( .A(n44094), .B(n44270), .Z(n44098) );
  XOR U6967 ( .A(n43893), .B(n44069), .Z(n43897) );
  XOR U6968 ( .A(n43473), .B(n43649), .Z(n43477) );
  XOR U6969 ( .A(n43254), .B(n43430), .Z(n43258) );
  XOR U6970 ( .A(n43029), .B(n43205), .Z(n43033) );
  XOR U6971 ( .A(n42798), .B(n42974), .Z(n42802) );
  XOR U6972 ( .A(n42561), .B(n42737), .Z(n42565) );
  XOR U6973 ( .A(n42318), .B(n42494), .Z(n42322) );
  XOR U6974 ( .A(n42069), .B(n42245), .Z(n42073) );
  XOR U6975 ( .A(n41814), .B(n41990), .Z(n41818) );
  XOR U6976 ( .A(n41553), .B(n41729), .Z(n41557) );
  XOR U6977 ( .A(n41286), .B(n41462), .Z(n41290) );
  XOR U6978 ( .A(n41013), .B(n41189), .Z(n41017) );
  XOR U6979 ( .A(n40734), .B(n40910), .Z(n40738) );
  XOR U6980 ( .A(n40449), .B(n40625), .Z(n40453) );
  XOR U6981 ( .A(n40158), .B(n40334), .Z(n40162) );
  XOR U6982 ( .A(n39861), .B(n40037), .Z(n39865) );
  XOR U6983 ( .A(n39558), .B(n39734), .Z(n39562) );
  XOR U6984 ( .A(n39249), .B(n39425), .Z(n39253) );
  XOR U6985 ( .A(n38934), .B(n39110), .Z(n38938) );
  XOR U6986 ( .A(n38613), .B(n38789), .Z(n38617) );
  XOR U6987 ( .A(n38286), .B(n38462), .Z(n38290) );
  XOR U6988 ( .A(n37953), .B(n38129), .Z(n37957) );
  XOR U6989 ( .A(n37614), .B(n37790), .Z(n37618) );
  XOR U6990 ( .A(n37269), .B(n37445), .Z(n37273) );
  XOR U6991 ( .A(n36918), .B(n37094), .Z(n36922) );
  XOR U6992 ( .A(n36561), .B(n36737), .Z(n36565) );
  XOR U6993 ( .A(n36198), .B(n36374), .Z(n36202) );
  XOR U6994 ( .A(n35829), .B(n36005), .Z(n35833) );
  XOR U6995 ( .A(n35454), .B(n35630), .Z(n35458) );
  XOR U6996 ( .A(n35073), .B(n35249), .Z(n35077) );
  XOR U6997 ( .A(n34686), .B(n34862), .Z(n34690) );
  XOR U6998 ( .A(n34293), .B(n34469), .Z(n34297) );
  XOR U6999 ( .A(n33894), .B(n34070), .Z(n33898) );
  XOR U7000 ( .A(n33489), .B(n33665), .Z(n33493) );
  XOR U7001 ( .A(n33078), .B(n33254), .Z(n33082) );
  XOR U7002 ( .A(n32661), .B(n32837), .Z(n32665) );
  XOR U7003 ( .A(n32238), .B(n32414), .Z(n32242) );
  XOR U7004 ( .A(n31809), .B(n31985), .Z(n31813) );
  XOR U7005 ( .A(n31374), .B(n31550), .Z(n31378) );
  XOR U7006 ( .A(n30933), .B(n31109), .Z(n30937) );
  XOR U7007 ( .A(n30486), .B(n30662), .Z(n30490) );
  XOR U7008 ( .A(n30033), .B(n30209), .Z(n30037) );
  XOR U7009 ( .A(n29574), .B(n29750), .Z(n29578) );
  XOR U7010 ( .A(n29109), .B(n29285), .Z(n29113) );
  XOR U7011 ( .A(n28638), .B(n28814), .Z(n28642) );
  XOR U7012 ( .A(n28161), .B(n28337), .Z(n28165) );
  XOR U7013 ( .A(n27678), .B(n27854), .Z(n27682) );
  XOR U7014 ( .A(n27189), .B(n27365), .Z(n27193) );
  XOR U7015 ( .A(n26692), .B(n26868), .Z(n26696) );
  XOR U7016 ( .A(n26191), .B(n26367), .Z(n26195) );
  XOR U7017 ( .A(n25683), .B(n25859), .Z(n25687) );
  XOR U7018 ( .A(n25169), .B(n25345), .Z(n25173) );
  XOR U7019 ( .A(n24646), .B(n24822), .Z(n24650) );
  XOR U7020 ( .A(n24121), .B(n24297), .Z(n24125) );
  XOR U7021 ( .A(n23590), .B(n23766), .Z(n23594) );
  XOR U7022 ( .A(n23052), .B(n23228), .Z(n23056) );
  XOR U7023 ( .A(n22508), .B(n22684), .Z(n22512) );
  XOR U7024 ( .A(n21959), .B(n22135), .Z(n21963) );
  XOR U7025 ( .A(n21404), .B(n21580), .Z(n21408) );
  XOR U7026 ( .A(n20842), .B(n21018), .Z(n20846) );
  XOR U7027 ( .A(n20275), .B(n20451), .Z(n20279) );
  XOR U7028 ( .A(n19702), .B(n19878), .Z(n19706) );
  XOR U7029 ( .A(n19123), .B(n19299), .Z(n19127) );
  XOR U7030 ( .A(n18434), .B(n18645), .Z(n18438) );
  XOR U7031 ( .A(n17244), .B(n17421), .Z(n17248) );
  XOR U7032 ( .A(n16030), .B(n16207), .Z(n16034) );
  XOR U7033 ( .A(n14792), .B(n14969), .Z(n14796) );
  XOR U7034 ( .A(n13530), .B(n13707), .Z(n13534) );
  XOR U7035 ( .A(n9528), .B(n9789), .Z(n9532) );
  XOR U7036 ( .A(n8150), .B(n8435), .Z(n8154) );
  XOR U7037 ( .A(n8105), .B(n8444), .Z(n8109) );
  XOR U7038 ( .A(n6703), .B(n7066), .Z(n6707) );
  XOR U7039 ( .A(n6658), .B(n7075), .Z(n6662) );
  XOR U7040 ( .A(n3001), .B(n3532), .Z(n3005) );
  XOR U7041 ( .A(n1515), .B(n2070), .Z(n1519) );
  XOR U7042 ( .A(n1470), .B(n2079), .Z(n1474) );
  XOR U7043 ( .A(n12895), .B(n13066), .Z(n12899) );
  XOR U7044 ( .A(n11595), .B(n11766), .Z(n11599) );
  XOR U7045 ( .A(n10213), .B(n10456), .Z(n10217) );
  XOR U7046 ( .A(n5280), .B(n5663), .Z(n5284) );
  XOR U7047 ( .A(n5235), .B(n5672), .Z(n5239) );
  XOR U7048 ( .A(n3740), .B(n4253), .Z(n3744) );
  XOR U7049 ( .A(n1500), .B(n2073), .Z(n1504) );
  XOR U7050 ( .A(n3031), .B(n3526), .Z(n3035) );
  XOR U7051 ( .A(n1545), .B(n2064), .Z(n1549) );
  XOR U7052 ( .A(n6688), .B(n7069), .Z(n6692) );
  XOR U7053 ( .A(n8135), .B(n8438), .Z(n8139) );
  XOR U7054 ( .A(n6733), .B(n7060), .Z(n6737) );
  XOR U7055 ( .A(n9558), .B(n9783), .Z(n9562) );
  XOR U7056 ( .A(n8180), .B(n8429), .Z(n8184) );
  XOR U7057 ( .A(n3770), .B(n4247), .Z(n3774) );
  XOR U7058 ( .A(n5265), .B(n5666), .Z(n5269) );
  XOR U7059 ( .A(n5310), .B(n5657), .Z(n5314) );
  XOR U7060 ( .A(n10243), .B(n10450), .Z(n10247) );
  XOR U7061 ( .A(n45189), .B(n45347), .Z(n45193) );
  XOR U7062 ( .A(n45024), .B(n45182), .Z(n45028) );
  XOR U7063 ( .A(n44853), .B(n45011), .Z(n44857) );
  XOR U7064 ( .A(n44676), .B(n44834), .Z(n44680) );
  XOR U7065 ( .A(n44493), .B(n44651), .Z(n44497) );
  XOR U7066 ( .A(n44109), .B(n44267), .Z(n44113) );
  XOR U7067 ( .A(n43908), .B(n44066), .Z(n43912) );
  XOR U7068 ( .A(n43701), .B(n43859), .Z(n43705) );
  XOR U7069 ( .A(n43488), .B(n43646), .Z(n43492) );
  XOR U7070 ( .A(n43269), .B(n43427), .Z(n43273) );
  XOR U7071 ( .A(n43044), .B(n43202), .Z(n43048) );
  XOR U7072 ( .A(n42813), .B(n42971), .Z(n42817) );
  XOR U7073 ( .A(n42576), .B(n42734), .Z(n42580) );
  XOR U7074 ( .A(n42333), .B(n42491), .Z(n42337) );
  XOR U7075 ( .A(n42084), .B(n42242), .Z(n42088) );
  XOR U7076 ( .A(n41829), .B(n41987), .Z(n41833) );
  XOR U7077 ( .A(n41568), .B(n41726), .Z(n41572) );
  XOR U7078 ( .A(n41301), .B(n41459), .Z(n41305) );
  XOR U7079 ( .A(n41028), .B(n41186), .Z(n41032) );
  XOR U7080 ( .A(n40749), .B(n40907), .Z(n40753) );
  XOR U7081 ( .A(n40464), .B(n40622), .Z(n40468) );
  XOR U7082 ( .A(n40173), .B(n40331), .Z(n40177) );
  XOR U7083 ( .A(n39876), .B(n40034), .Z(n39880) );
  XOR U7084 ( .A(n39573), .B(n39731), .Z(n39577) );
  XOR U7085 ( .A(n39264), .B(n39422), .Z(n39268) );
  XOR U7086 ( .A(n38949), .B(n39107), .Z(n38953) );
  XOR U7087 ( .A(n38628), .B(n38786), .Z(n38632) );
  XOR U7088 ( .A(n38301), .B(n38459), .Z(n38305) );
  XOR U7089 ( .A(n37968), .B(n38126), .Z(n37972) );
  XOR U7090 ( .A(n37629), .B(n37787), .Z(n37633) );
  XOR U7091 ( .A(n37284), .B(n37442), .Z(n37288) );
  XOR U7092 ( .A(n36933), .B(n37091), .Z(n36937) );
  XOR U7093 ( .A(n36576), .B(n36734), .Z(n36580) );
  XOR U7094 ( .A(n36213), .B(n36371), .Z(n36217) );
  XOR U7095 ( .A(n35844), .B(n36002), .Z(n35848) );
  XOR U7096 ( .A(n35469), .B(n35627), .Z(n35473) );
  XOR U7097 ( .A(n35088), .B(n35246), .Z(n35092) );
  XOR U7098 ( .A(n34701), .B(n34859), .Z(n34705) );
  XOR U7099 ( .A(n34308), .B(n34466), .Z(n34312) );
  XOR U7100 ( .A(n33909), .B(n34067), .Z(n33913) );
  XOR U7101 ( .A(n33504), .B(n33662), .Z(n33508) );
  XOR U7102 ( .A(n33093), .B(n33251), .Z(n33097) );
  XOR U7103 ( .A(n32676), .B(n32834), .Z(n32680) );
  XOR U7104 ( .A(n32253), .B(n32411), .Z(n32257) );
  XOR U7105 ( .A(n31824), .B(n31982), .Z(n31828) );
  XOR U7106 ( .A(n31389), .B(n31547), .Z(n31393) );
  XOR U7107 ( .A(n30948), .B(n31106), .Z(n30952) );
  XOR U7108 ( .A(n30501), .B(n30659), .Z(n30505) );
  XOR U7109 ( .A(n30048), .B(n30206), .Z(n30052) );
  XOR U7110 ( .A(n29589), .B(n29747), .Z(n29593) );
  XOR U7111 ( .A(n29124), .B(n29282), .Z(n29128) );
  XOR U7112 ( .A(n28653), .B(n28811), .Z(n28657) );
  XOR U7113 ( .A(n28176), .B(n28334), .Z(n28180) );
  XOR U7114 ( .A(n27693), .B(n27851), .Z(n27697) );
  XOR U7115 ( .A(n27204), .B(n27362), .Z(n27208) );
  XOR U7116 ( .A(n26707), .B(n26865), .Z(n26711) );
  XOR U7117 ( .A(n26206), .B(n26364), .Z(n26210) );
  XOR U7118 ( .A(n25698), .B(n25856), .Z(n25702) );
  XOR U7119 ( .A(n25184), .B(n25342), .Z(n25188) );
  XOR U7120 ( .A(n24661), .B(n24819), .Z(n24665) );
  XOR U7121 ( .A(n24136), .B(n24294), .Z(n24140) );
  XOR U7122 ( .A(n23605), .B(n23763), .Z(n23609) );
  XOR U7123 ( .A(n23067), .B(n23225), .Z(n23071) );
  XOR U7124 ( .A(n22523), .B(n22681), .Z(n22527) );
  XOR U7125 ( .A(n21974), .B(n22132), .Z(n21978) );
  XOR U7126 ( .A(n21419), .B(n21577), .Z(n21423) );
  XOR U7127 ( .A(n20857), .B(n21015), .Z(n20861) );
  XOR U7128 ( .A(n20290), .B(n20448), .Z(n20294) );
  XOR U7129 ( .A(n19717), .B(n19875), .Z(n19721) );
  XOR U7130 ( .A(n19138), .B(n19296), .Z(n19142) );
  XOR U7131 ( .A(n17857), .B(n18016), .Z(n17861) );
  XOR U7132 ( .A(n16655), .B(n16814), .Z(n16659) );
  XOR U7133 ( .A(n15429), .B(n15588), .Z(n15433) );
  XOR U7134 ( .A(n9588), .B(n9777), .Z(n9592) );
  XOR U7135 ( .A(n8210), .B(n8423), .Z(n8214) );
  XOR U7136 ( .A(n8165), .B(n8432), .Z(n8169) );
  XOR U7137 ( .A(n6763), .B(n7054), .Z(n6767) );
  XOR U7138 ( .A(n6718), .B(n7063), .Z(n6722) );
  XOR U7139 ( .A(n3061), .B(n3520), .Z(n3065) );
  XOR U7140 ( .A(n1575), .B(n2058), .Z(n1579) );
  XOR U7141 ( .A(n1530), .B(n2067), .Z(n1534) );
  XOR U7142 ( .A(n14812), .B(n14965), .Z(n14816) );
  XOR U7143 ( .A(n13550), .B(n13703), .Z(n13554) );
  XOR U7144 ( .A(n12262), .B(n12417), .Z(n12266) );
  XOR U7145 ( .A(n10952), .B(n11105), .Z(n10956) );
  XOR U7146 ( .A(n10273), .B(n10444), .Z(n10277) );
  XOR U7147 ( .A(n5340), .B(n5651), .Z(n5344) );
  XOR U7148 ( .A(n5295), .B(n5660), .Z(n5299) );
  XOR U7149 ( .A(n3800), .B(n4241), .Z(n3804) );
  XOR U7150 ( .A(n1560), .B(n2061), .Z(n1564) );
  XOR U7151 ( .A(n3091), .B(n3514), .Z(n3095) );
  XOR U7152 ( .A(n1605), .B(n2052), .Z(n1609) );
  XOR U7153 ( .A(n6748), .B(n7057), .Z(n6752) );
  XOR U7154 ( .A(n8195), .B(n8426), .Z(n8199) );
  XOR U7155 ( .A(n6793), .B(n7048), .Z(n6797) );
  XOR U7156 ( .A(n8240), .B(n8417), .Z(n8244) );
  XOR U7157 ( .A(n10293), .B(n10440), .Z(n10297) );
  XOR U7158 ( .A(n3830), .B(n4235), .Z(n3834) );
  XOR U7159 ( .A(n5325), .B(n5654), .Z(n5329) );
  XOR U7160 ( .A(n5370), .B(n5645), .Z(n5374) );
  XOR U7161 ( .A(n45663), .B(n45803), .Z(n45667) );
  XOR U7162 ( .A(n45516), .B(n45656), .Z(n45520) );
  XOR U7163 ( .A(n45363), .B(n45503), .Z(n45367) );
  XOR U7164 ( .A(n45204), .B(n45344), .Z(n45208) );
  XOR U7165 ( .A(n45039), .B(n45179), .Z(n45043) );
  XOR U7166 ( .A(n44691), .B(n44831), .Z(n44695) );
  XOR U7167 ( .A(n44508), .B(n44648), .Z(n44512) );
  XOR U7168 ( .A(n44319), .B(n44459), .Z(n44323) );
  XOR U7169 ( .A(n44124), .B(n44264), .Z(n44128) );
  XOR U7170 ( .A(n43923), .B(n44063), .Z(n43927) );
  XOR U7171 ( .A(n43716), .B(n43856), .Z(n43720) );
  XOR U7172 ( .A(n43503), .B(n43643), .Z(n43507) );
  XOR U7173 ( .A(n43284), .B(n43424), .Z(n43288) );
  XOR U7174 ( .A(n43059), .B(n43199), .Z(n43063) );
  XOR U7175 ( .A(n42828), .B(n42968), .Z(n42832) );
  XOR U7176 ( .A(n42591), .B(n42731), .Z(n42595) );
  XOR U7177 ( .A(n42348), .B(n42488), .Z(n42352) );
  XOR U7178 ( .A(n42099), .B(n42239), .Z(n42103) );
  XOR U7179 ( .A(n41844), .B(n41984), .Z(n41848) );
  XOR U7180 ( .A(n41583), .B(n41723), .Z(n41587) );
  XOR U7181 ( .A(n41316), .B(n41456), .Z(n41320) );
  XOR U7182 ( .A(n41043), .B(n41183), .Z(n41047) );
  XOR U7183 ( .A(n40764), .B(n40904), .Z(n40768) );
  XOR U7184 ( .A(n40479), .B(n40619), .Z(n40483) );
  XOR U7185 ( .A(n40188), .B(n40328), .Z(n40192) );
  XOR U7186 ( .A(n39891), .B(n40031), .Z(n39895) );
  XOR U7187 ( .A(n39588), .B(n39728), .Z(n39592) );
  XOR U7188 ( .A(n39279), .B(n39419), .Z(n39283) );
  XOR U7189 ( .A(n38964), .B(n39104), .Z(n38968) );
  XOR U7190 ( .A(n38643), .B(n38783), .Z(n38647) );
  XOR U7191 ( .A(n38316), .B(n38456), .Z(n38320) );
  XOR U7192 ( .A(n37983), .B(n38123), .Z(n37987) );
  XOR U7193 ( .A(n37644), .B(n37784), .Z(n37648) );
  XOR U7194 ( .A(n37299), .B(n37439), .Z(n37303) );
  XOR U7195 ( .A(n36948), .B(n37088), .Z(n36952) );
  XOR U7196 ( .A(n36591), .B(n36731), .Z(n36595) );
  XOR U7197 ( .A(n36228), .B(n36368), .Z(n36232) );
  XOR U7198 ( .A(n35859), .B(n35999), .Z(n35863) );
  XOR U7199 ( .A(n35484), .B(n35624), .Z(n35488) );
  XOR U7200 ( .A(n35103), .B(n35243), .Z(n35107) );
  XOR U7201 ( .A(n34716), .B(n34856), .Z(n34720) );
  XOR U7202 ( .A(n34323), .B(n34463), .Z(n34327) );
  XOR U7203 ( .A(n33924), .B(n34064), .Z(n33928) );
  XOR U7204 ( .A(n33519), .B(n33659), .Z(n33523) );
  XOR U7205 ( .A(n33108), .B(n33248), .Z(n33112) );
  XOR U7206 ( .A(n32691), .B(n32831), .Z(n32695) );
  XOR U7207 ( .A(n32268), .B(n32408), .Z(n32272) );
  XOR U7208 ( .A(n31839), .B(n31979), .Z(n31843) );
  XOR U7209 ( .A(n31404), .B(n31544), .Z(n31408) );
  XOR U7210 ( .A(n30963), .B(n31103), .Z(n30967) );
  XOR U7211 ( .A(n30516), .B(n30656), .Z(n30520) );
  XOR U7212 ( .A(n30063), .B(n30203), .Z(n30067) );
  XOR U7213 ( .A(n29604), .B(n29744), .Z(n29608) );
  XOR U7214 ( .A(n29139), .B(n29279), .Z(n29143) );
  XOR U7215 ( .A(n28668), .B(n28808), .Z(n28672) );
  XOR U7216 ( .A(n28191), .B(n28331), .Z(n28195) );
  XOR U7217 ( .A(n27708), .B(n27848), .Z(n27712) );
  XOR U7218 ( .A(n27219), .B(n27359), .Z(n27223) );
  XOR U7219 ( .A(n26722), .B(n26862), .Z(n26726) );
  XOR U7220 ( .A(n26221), .B(n26361), .Z(n26225) );
  XOR U7221 ( .A(n25713), .B(n25853), .Z(n25717) );
  XOR U7222 ( .A(n25199), .B(n25339), .Z(n25203) );
  XOR U7223 ( .A(n24676), .B(n24816), .Z(n24680) );
  XOR U7224 ( .A(n24151), .B(n24291), .Z(n24155) );
  XOR U7225 ( .A(n23620), .B(n23760), .Z(n23624) );
  XOR U7226 ( .A(n23082), .B(n23222), .Z(n23086) );
  XOR U7227 ( .A(n22538), .B(n22678), .Z(n22542) );
  XOR U7228 ( .A(n21989), .B(n22129), .Z(n21993) );
  XOR U7229 ( .A(n21434), .B(n21574), .Z(n21438) );
  XOR U7230 ( .A(n20872), .B(n21012), .Z(n20876) );
  XOR U7231 ( .A(n20305), .B(n20445), .Z(n20309) );
  XOR U7232 ( .A(n19732), .B(n19872), .Z(n19736) );
  XOR U7233 ( .A(n19153), .B(n19293), .Z(n19157) );
  XOR U7234 ( .A(n17872), .B(n18013), .Z(n17876) );
  XOR U7235 ( .A(n16670), .B(n16811), .Z(n16674) );
  XOR U7236 ( .A(n8225), .B(n8420), .Z(n8229) );
  XOR U7237 ( .A(n6823), .B(n7042), .Z(n6827) );
  XOR U7238 ( .A(n6778), .B(n7051), .Z(n6782) );
  XOR U7239 ( .A(n3121), .B(n3508), .Z(n3125) );
  XOR U7240 ( .A(n1635), .B(n2046), .Z(n1639) );
  XOR U7241 ( .A(n1590), .B(n2055), .Z(n1594) );
  XOR U7242 ( .A(n15449), .B(n15584), .Z(n15453) );
  XOR U7243 ( .A(n14199), .B(n14334), .Z(n14203) );
  XOR U7244 ( .A(n12925), .B(n13060), .Z(n12929) );
  XOR U7245 ( .A(n8957), .B(n9092), .Z(n8961) );
  XOR U7246 ( .A(n5400), .B(n5639), .Z(n5404) );
  XOR U7247 ( .A(n5355), .B(n5648), .Z(n5359) );
  XOR U7248 ( .A(n3860), .B(n4229), .Z(n3864) );
  XOR U7249 ( .A(n1620), .B(n2049), .Z(n1624) );
  XOR U7250 ( .A(n3151), .B(n3502), .Z(n3155) );
  XOR U7251 ( .A(n1665), .B(n2040), .Z(n1669) );
  XOR U7252 ( .A(n6808), .B(n7045), .Z(n6812) );
  XOR U7253 ( .A(n8255), .B(n8414), .Z(n8259) );
  XOR U7254 ( .A(n6853), .B(n7036), .Z(n6857) );
  XOR U7255 ( .A(n12282), .B(n12413), .Z(n12286) );
  XOR U7256 ( .A(n10972), .B(n11101), .Z(n10976) );
  XOR U7257 ( .A(n3890), .B(n4223), .Z(n3894) );
  XOR U7258 ( .A(n5385), .B(n5642), .Z(n5389) );
  XOR U7259 ( .A(n5430), .B(n5633), .Z(n5434) );
  XOR U7260 ( .A(n46083), .B(n46205), .Z(n46087) );
  XOR U7261 ( .A(n45954), .B(n46076), .Z(n45958) );
  XOR U7262 ( .A(n45819), .B(n45941), .Z(n45823) );
  XOR U7263 ( .A(n45678), .B(n45800), .Z(n45682) );
  XOR U7264 ( .A(n45531), .B(n45653), .Z(n45535) );
  XOR U7265 ( .A(n45219), .B(n45341), .Z(n45223) );
  XOR U7266 ( .A(n45054), .B(n45176), .Z(n45058) );
  XOR U7267 ( .A(n44883), .B(n45005), .Z(n44887) );
  XOR U7268 ( .A(n44706), .B(n44828), .Z(n44710) );
  XOR U7269 ( .A(n44523), .B(n44645), .Z(n44527) );
  XOR U7270 ( .A(n44334), .B(n44456), .Z(n44338) );
  XOR U7271 ( .A(n44139), .B(n44261), .Z(n44143) );
  XOR U7272 ( .A(n43938), .B(n44060), .Z(n43942) );
  XOR U7273 ( .A(n43731), .B(n43853), .Z(n43735) );
  XOR U7274 ( .A(n43518), .B(n43640), .Z(n43522) );
  XOR U7275 ( .A(n43299), .B(n43421), .Z(n43303) );
  XOR U7276 ( .A(n43074), .B(n43196), .Z(n43078) );
  XOR U7277 ( .A(n42843), .B(n42965), .Z(n42847) );
  XOR U7278 ( .A(n42606), .B(n42728), .Z(n42610) );
  XOR U7279 ( .A(n42363), .B(n42485), .Z(n42367) );
  XOR U7280 ( .A(n42114), .B(n42236), .Z(n42118) );
  XOR U7281 ( .A(n41859), .B(n41981), .Z(n41863) );
  XOR U7282 ( .A(n41598), .B(n41720), .Z(n41602) );
  XOR U7283 ( .A(n41331), .B(n41453), .Z(n41335) );
  XOR U7284 ( .A(n41058), .B(n41180), .Z(n41062) );
  XOR U7285 ( .A(n40779), .B(n40901), .Z(n40783) );
  XOR U7286 ( .A(n40494), .B(n40616), .Z(n40498) );
  XOR U7287 ( .A(n40203), .B(n40325), .Z(n40207) );
  XOR U7288 ( .A(n39906), .B(n40028), .Z(n39910) );
  XOR U7289 ( .A(n39603), .B(n39725), .Z(n39607) );
  XOR U7290 ( .A(n39294), .B(n39416), .Z(n39298) );
  XOR U7291 ( .A(n38979), .B(n39101), .Z(n38983) );
  XOR U7292 ( .A(n38658), .B(n38780), .Z(n38662) );
  XOR U7293 ( .A(n38331), .B(n38453), .Z(n38335) );
  XOR U7294 ( .A(n37998), .B(n38120), .Z(n38002) );
  XOR U7295 ( .A(n37659), .B(n37781), .Z(n37663) );
  XOR U7296 ( .A(n37314), .B(n37436), .Z(n37318) );
  XOR U7297 ( .A(n36963), .B(n37085), .Z(n36967) );
  XOR U7298 ( .A(n36606), .B(n36728), .Z(n36610) );
  XOR U7299 ( .A(n36243), .B(n36365), .Z(n36247) );
  XOR U7300 ( .A(n35874), .B(n35996), .Z(n35878) );
  XOR U7301 ( .A(n35499), .B(n35621), .Z(n35503) );
  XOR U7302 ( .A(n35118), .B(n35240), .Z(n35122) );
  XOR U7303 ( .A(n34731), .B(n34853), .Z(n34735) );
  XOR U7304 ( .A(n34338), .B(n34460), .Z(n34342) );
  XOR U7305 ( .A(n33939), .B(n34061), .Z(n33943) );
  XOR U7306 ( .A(n33534), .B(n33656), .Z(n33538) );
  XOR U7307 ( .A(n33123), .B(n33245), .Z(n33127) );
  XOR U7308 ( .A(n32706), .B(n32828), .Z(n32710) );
  XOR U7309 ( .A(n32283), .B(n32405), .Z(n32287) );
  XOR U7310 ( .A(n31854), .B(n31976), .Z(n31858) );
  XOR U7311 ( .A(n31419), .B(n31541), .Z(n31423) );
  XOR U7312 ( .A(n30978), .B(n31100), .Z(n30982) );
  XOR U7313 ( .A(n30531), .B(n30653), .Z(n30535) );
  XOR U7314 ( .A(n30078), .B(n30200), .Z(n30082) );
  XOR U7315 ( .A(n29619), .B(n29741), .Z(n29623) );
  XOR U7316 ( .A(n29154), .B(n29276), .Z(n29158) );
  XOR U7317 ( .A(n28683), .B(n28805), .Z(n28687) );
  XOR U7318 ( .A(n28206), .B(n28328), .Z(n28210) );
  XOR U7319 ( .A(n27723), .B(n27845), .Z(n27727) );
  XOR U7320 ( .A(n27234), .B(n27356), .Z(n27238) );
  XOR U7321 ( .A(n26737), .B(n26859), .Z(n26741) );
  XOR U7322 ( .A(n26236), .B(n26358), .Z(n26240) );
  XOR U7323 ( .A(n25728), .B(n25850), .Z(n25732) );
  XOR U7324 ( .A(n25214), .B(n25336), .Z(n25218) );
  XOR U7325 ( .A(n24691), .B(n24813), .Z(n24695) );
  XOR U7326 ( .A(n24166), .B(n24288), .Z(n24170) );
  XOR U7327 ( .A(n23635), .B(n23757), .Z(n23639) );
  XOR U7328 ( .A(n23097), .B(n23219), .Z(n23101) );
  XOR U7329 ( .A(n22553), .B(n22675), .Z(n22557) );
  XOR U7330 ( .A(n22004), .B(n22126), .Z(n22008) );
  XOR U7331 ( .A(n21449), .B(n21571), .Z(n21453) );
  XOR U7332 ( .A(n20887), .B(n21009), .Z(n20891) );
  XOR U7333 ( .A(n20320), .B(n20442), .Z(n20324) );
  XOR U7334 ( .A(n19747), .B(n19869), .Z(n19751) );
  XOR U7335 ( .A(n19168), .B(n19290), .Z(n19172) );
  XOR U7336 ( .A(n17887), .B(n18010), .Z(n17891) );
  XOR U7337 ( .A(n6883), .B(n7030), .Z(n6887) );
  XOR U7338 ( .A(n6838), .B(n7039), .Z(n6842) );
  XOR U7339 ( .A(n3181), .B(n3496), .Z(n3185) );
  XOR U7340 ( .A(n1695), .B(n2034), .Z(n1699) );
  XOR U7341 ( .A(n1650), .B(n2043), .Z(n1654) );
  XOR U7342 ( .A(n16690), .B(n16807), .Z(n16694) );
  XOR U7343 ( .A(n15464), .B(n15581), .Z(n15468) );
  XOR U7344 ( .A(n14214), .B(n14331), .Z(n14218) );
  XOR U7345 ( .A(n9648), .B(n9765), .Z(n9652) );
  XOR U7346 ( .A(n5460), .B(n5627), .Z(n5464) );
  XOR U7347 ( .A(n5415), .B(n5636), .Z(n5419) );
  XOR U7348 ( .A(n3920), .B(n4217), .Z(n3924) );
  XOR U7349 ( .A(n1680), .B(n2037), .Z(n1684) );
  XOR U7350 ( .A(n3211), .B(n3490), .Z(n3215) );
  XOR U7351 ( .A(n1725), .B(n2028), .Z(n1729) );
  XOR U7352 ( .A(n6868), .B(n7033), .Z(n6872) );
  XOR U7353 ( .A(n13585), .B(n13696), .Z(n13589) );
  XOR U7354 ( .A(n12297), .B(n12410), .Z(n12301) );
  XOR U7355 ( .A(n10987), .B(n11098), .Z(n10991) );
  XOR U7356 ( .A(n8977), .B(n9088), .Z(n8981) );
  XOR U7357 ( .A(n7607), .B(n7718), .Z(n7611) );
  XOR U7358 ( .A(n3950), .B(n4211), .Z(n3954) );
  XOR U7359 ( .A(n5445), .B(n5630), .Z(n5449) );
  XOR U7360 ( .A(n5490), .B(n5621), .Z(n5494) );
  XOR U7361 ( .A(n46449), .B(n46553), .Z(n46453) );
  XOR U7362 ( .A(n46338), .B(n46442), .Z(n46342) );
  XOR U7363 ( .A(n46221), .B(n46325), .Z(n46225) );
  XOR U7364 ( .A(n46098), .B(n46202), .Z(n46102) );
  XOR U7365 ( .A(n45969), .B(n46073), .Z(n45973) );
  XOR U7366 ( .A(n45693), .B(n45797), .Z(n45697) );
  XOR U7367 ( .A(n45546), .B(n45650), .Z(n45550) );
  XOR U7368 ( .A(n45393), .B(n45497), .Z(n45397) );
  XOR U7369 ( .A(n45234), .B(n45338), .Z(n45238) );
  XOR U7370 ( .A(n45069), .B(n45173), .Z(n45073) );
  XOR U7371 ( .A(n44898), .B(n45002), .Z(n44902) );
  XOR U7372 ( .A(n44721), .B(n44825), .Z(n44725) );
  XOR U7373 ( .A(n44538), .B(n44642), .Z(n44542) );
  XOR U7374 ( .A(n44349), .B(n44453), .Z(n44353) );
  XOR U7375 ( .A(n44154), .B(n44258), .Z(n44158) );
  XOR U7376 ( .A(n43953), .B(n44057), .Z(n43957) );
  XOR U7377 ( .A(n43746), .B(n43850), .Z(n43750) );
  XOR U7378 ( .A(n43533), .B(n43637), .Z(n43537) );
  XOR U7379 ( .A(n43314), .B(n43418), .Z(n43318) );
  XOR U7380 ( .A(n43089), .B(n43193), .Z(n43093) );
  XOR U7381 ( .A(n42858), .B(n42962), .Z(n42862) );
  XOR U7382 ( .A(n42621), .B(n42725), .Z(n42625) );
  XOR U7383 ( .A(n42378), .B(n42482), .Z(n42382) );
  XOR U7384 ( .A(n42129), .B(n42233), .Z(n42133) );
  XOR U7385 ( .A(n41874), .B(n41978), .Z(n41878) );
  XOR U7386 ( .A(n41613), .B(n41717), .Z(n41617) );
  XOR U7387 ( .A(n41346), .B(n41450), .Z(n41350) );
  XOR U7388 ( .A(n41073), .B(n41177), .Z(n41077) );
  XOR U7389 ( .A(n40794), .B(n40898), .Z(n40798) );
  XOR U7390 ( .A(n40509), .B(n40613), .Z(n40513) );
  XOR U7391 ( .A(n40218), .B(n40322), .Z(n40222) );
  XOR U7392 ( .A(n39921), .B(n40025), .Z(n39925) );
  XOR U7393 ( .A(n39618), .B(n39722), .Z(n39622) );
  XOR U7394 ( .A(n39309), .B(n39413), .Z(n39313) );
  XOR U7395 ( .A(n38994), .B(n39098), .Z(n38998) );
  XOR U7396 ( .A(n38673), .B(n38777), .Z(n38677) );
  XOR U7397 ( .A(n38346), .B(n38450), .Z(n38350) );
  XOR U7398 ( .A(n38013), .B(n38117), .Z(n38017) );
  XOR U7399 ( .A(n37674), .B(n37778), .Z(n37678) );
  XOR U7400 ( .A(n37329), .B(n37433), .Z(n37333) );
  XOR U7401 ( .A(n36978), .B(n37082), .Z(n36982) );
  XOR U7402 ( .A(n36621), .B(n36725), .Z(n36625) );
  XOR U7403 ( .A(n36258), .B(n36362), .Z(n36262) );
  XOR U7404 ( .A(n35889), .B(n35993), .Z(n35893) );
  XOR U7405 ( .A(n35514), .B(n35618), .Z(n35518) );
  XOR U7406 ( .A(n35133), .B(n35237), .Z(n35137) );
  XOR U7407 ( .A(n34746), .B(n34850), .Z(n34750) );
  XOR U7408 ( .A(n34353), .B(n34457), .Z(n34357) );
  XOR U7409 ( .A(n33954), .B(n34058), .Z(n33958) );
  XOR U7410 ( .A(n33549), .B(n33653), .Z(n33553) );
  XOR U7411 ( .A(n33138), .B(n33242), .Z(n33142) );
  XOR U7412 ( .A(n32721), .B(n32825), .Z(n32725) );
  XOR U7413 ( .A(n32298), .B(n32402), .Z(n32302) );
  XOR U7414 ( .A(n31869), .B(n31973), .Z(n31873) );
  XOR U7415 ( .A(n31434), .B(n31538), .Z(n31438) );
  XOR U7416 ( .A(n30993), .B(n31097), .Z(n30997) );
  XOR U7417 ( .A(n30546), .B(n30650), .Z(n30550) );
  XOR U7418 ( .A(n30093), .B(n30197), .Z(n30097) );
  XOR U7419 ( .A(n29634), .B(n29738), .Z(n29638) );
  XOR U7420 ( .A(n29169), .B(n29273), .Z(n29173) );
  XOR U7421 ( .A(n28698), .B(n28802), .Z(n28702) );
  XOR U7422 ( .A(n28221), .B(n28325), .Z(n28225) );
  XOR U7423 ( .A(n27738), .B(n27842), .Z(n27742) );
  XOR U7424 ( .A(n27249), .B(n27353), .Z(n27253) );
  XOR U7425 ( .A(n26752), .B(n26856), .Z(n26756) );
  XOR U7426 ( .A(n26251), .B(n26355), .Z(n26255) );
  XOR U7427 ( .A(n25743), .B(n25847), .Z(n25747) );
  XOR U7428 ( .A(n25229), .B(n25333), .Z(n25233) );
  XOR U7429 ( .A(n24706), .B(n24810), .Z(n24710) );
  XOR U7430 ( .A(n24181), .B(n24285), .Z(n24185) );
  XOR U7431 ( .A(n23650), .B(n23754), .Z(n23654) );
  XOR U7432 ( .A(n23112), .B(n23216), .Z(n23116) );
  XOR U7433 ( .A(n22568), .B(n22672), .Z(n22572) );
  XOR U7434 ( .A(n22019), .B(n22123), .Z(n22023) );
  XOR U7435 ( .A(n21464), .B(n21568), .Z(n21468) );
  XOR U7436 ( .A(n20902), .B(n21006), .Z(n20906) );
  XOR U7437 ( .A(n20335), .B(n20439), .Z(n20339) );
  XOR U7438 ( .A(n19762), .B(n19866), .Z(n19766) );
  XOR U7439 ( .A(n19183), .B(n19287), .Z(n19187) );
  XOR U7440 ( .A(n18494), .B(n18621), .Z(n18498) );
  XOR U7441 ( .A(n6898), .B(n7027), .Z(n6902) );
  XOR U7442 ( .A(n3241), .B(n3484), .Z(n3245) );
  XOR U7443 ( .A(n1755), .B(n2022), .Z(n1759) );
  XOR U7444 ( .A(n1710), .B(n2031), .Z(n1714) );
  XOR U7445 ( .A(n17309), .B(n17408), .Z(n17313) );
  XOR U7446 ( .A(n16095), .B(n16194), .Z(n16099) );
  XOR U7447 ( .A(n5475), .B(n5624), .Z(n5479) );
  XOR U7448 ( .A(n3980), .B(n4205), .Z(n3984) );
  XOR U7449 ( .A(n1740), .B(n2025), .Z(n1744) );
  XOR U7450 ( .A(n3271), .B(n3478), .Z(n3275) );
  XOR U7451 ( .A(n1785), .B(n2016), .Z(n1789) );
  XOR U7452 ( .A(n15484), .B(n15577), .Z(n15488) );
  XOR U7453 ( .A(n14234), .B(n14327), .Z(n14238) );
  XOR U7454 ( .A(n12960), .B(n13053), .Z(n12964) );
  XOR U7455 ( .A(n11660), .B(n11753), .Z(n11664) );
  XOR U7456 ( .A(n10338), .B(n10431), .Z(n10342) );
  XOR U7457 ( .A(n8992), .B(n9085), .Z(n8996) );
  XOR U7458 ( .A(n7622), .B(n7715), .Z(n7626) );
  XOR U7459 ( .A(n6228), .B(n6321), .Z(n6232) );
  XOR U7460 ( .A(n4803), .B(n4902), .Z(n4807) );
  XOR U7461 ( .A(n4010), .B(n4199), .Z(n4014) );
  XOR U7462 ( .A(n5505), .B(n5618), .Z(n5509) );
  XOR U7463 ( .A(n46761), .B(n46847), .Z(n46765) );
  XOR U7464 ( .A(n46668), .B(n46754), .Z(n46672) );
  XOR U7465 ( .A(n46569), .B(n46655), .Z(n46573) );
  XOR U7466 ( .A(n46464), .B(n46550), .Z(n46468) );
  XOR U7467 ( .A(n46353), .B(n46439), .Z(n46357) );
  XOR U7468 ( .A(n46113), .B(n46199), .Z(n46117) );
  XOR U7469 ( .A(n45984), .B(n46070), .Z(n45988) );
  XOR U7470 ( .A(n45849), .B(n45935), .Z(n45853) );
  XOR U7471 ( .A(n45708), .B(n45794), .Z(n45712) );
  XOR U7472 ( .A(n45561), .B(n45647), .Z(n45565) );
  XOR U7473 ( .A(n45408), .B(n45494), .Z(n45412) );
  XOR U7474 ( .A(n45249), .B(n45335), .Z(n45253) );
  XOR U7475 ( .A(n45084), .B(n45170), .Z(n45088) );
  XOR U7476 ( .A(n44913), .B(n44999), .Z(n44917) );
  XOR U7477 ( .A(n44736), .B(n44822), .Z(n44740) );
  XOR U7478 ( .A(n44553), .B(n44639), .Z(n44557) );
  XOR U7479 ( .A(n44364), .B(n44450), .Z(n44368) );
  XOR U7480 ( .A(n44169), .B(n44255), .Z(n44173) );
  XOR U7481 ( .A(n43968), .B(n44054), .Z(n43972) );
  XOR U7482 ( .A(n43761), .B(n43847), .Z(n43765) );
  XOR U7483 ( .A(n43548), .B(n43634), .Z(n43552) );
  XOR U7484 ( .A(n43329), .B(n43415), .Z(n43333) );
  XOR U7485 ( .A(n43104), .B(n43190), .Z(n43108) );
  XOR U7486 ( .A(n42873), .B(n42959), .Z(n42877) );
  XOR U7487 ( .A(n42636), .B(n42722), .Z(n42640) );
  XOR U7488 ( .A(n42393), .B(n42479), .Z(n42397) );
  XOR U7489 ( .A(n42144), .B(n42230), .Z(n42148) );
  XOR U7490 ( .A(n41889), .B(n41975), .Z(n41893) );
  XOR U7491 ( .A(n41628), .B(n41714), .Z(n41632) );
  XOR U7492 ( .A(n41361), .B(n41447), .Z(n41365) );
  XOR U7493 ( .A(n41088), .B(n41174), .Z(n41092) );
  XOR U7494 ( .A(n40809), .B(n40895), .Z(n40813) );
  XOR U7495 ( .A(n40524), .B(n40610), .Z(n40528) );
  XOR U7496 ( .A(n40233), .B(n40319), .Z(n40237) );
  XOR U7497 ( .A(n39936), .B(n40022), .Z(n39940) );
  XOR U7498 ( .A(n39633), .B(n39719), .Z(n39637) );
  XOR U7499 ( .A(n39324), .B(n39410), .Z(n39328) );
  XOR U7500 ( .A(n39009), .B(n39095), .Z(n39013) );
  XOR U7501 ( .A(n38688), .B(n38774), .Z(n38692) );
  XOR U7502 ( .A(n38361), .B(n38447), .Z(n38365) );
  XOR U7503 ( .A(n38028), .B(n38114), .Z(n38032) );
  XOR U7504 ( .A(n37689), .B(n37775), .Z(n37693) );
  XOR U7505 ( .A(n37344), .B(n37430), .Z(n37348) );
  XOR U7506 ( .A(n36993), .B(n37079), .Z(n36997) );
  XOR U7507 ( .A(n36636), .B(n36722), .Z(n36640) );
  XOR U7508 ( .A(n36273), .B(n36359), .Z(n36277) );
  XOR U7509 ( .A(n35904), .B(n35990), .Z(n35908) );
  XOR U7510 ( .A(n35529), .B(n35615), .Z(n35533) );
  XOR U7511 ( .A(n35148), .B(n35234), .Z(n35152) );
  XOR U7512 ( .A(n34761), .B(n34847), .Z(n34765) );
  XOR U7513 ( .A(n34368), .B(n34454), .Z(n34372) );
  XOR U7514 ( .A(n33969), .B(n34055), .Z(n33973) );
  XOR U7515 ( .A(n33564), .B(n33650), .Z(n33568) );
  XOR U7516 ( .A(n33153), .B(n33239), .Z(n33157) );
  XOR U7517 ( .A(n32736), .B(n32822), .Z(n32740) );
  XOR U7518 ( .A(n32313), .B(n32399), .Z(n32317) );
  XOR U7519 ( .A(n31884), .B(n31970), .Z(n31888) );
  XOR U7520 ( .A(n31449), .B(n31535), .Z(n31453) );
  XOR U7521 ( .A(n31008), .B(n31094), .Z(n31012) );
  XOR U7522 ( .A(n30561), .B(n30647), .Z(n30565) );
  XOR U7523 ( .A(n30108), .B(n30194), .Z(n30112) );
  XOR U7524 ( .A(n29649), .B(n29735), .Z(n29653) );
  XOR U7525 ( .A(n29184), .B(n29270), .Z(n29188) );
  XOR U7526 ( .A(n28713), .B(n28799), .Z(n28717) );
  XOR U7527 ( .A(n28236), .B(n28322), .Z(n28240) );
  XOR U7528 ( .A(n27753), .B(n27839), .Z(n27757) );
  XOR U7529 ( .A(n27264), .B(n27350), .Z(n27268) );
  XOR U7530 ( .A(n26767), .B(n26853), .Z(n26771) );
  XOR U7531 ( .A(n26266), .B(n26352), .Z(n26270) );
  XOR U7532 ( .A(n25758), .B(n25844), .Z(n25762) );
  XOR U7533 ( .A(n25244), .B(n25330), .Z(n25248) );
  XOR U7534 ( .A(n24721), .B(n24807), .Z(n24725) );
  XOR U7535 ( .A(n24196), .B(n24282), .Z(n24200) );
  XOR U7536 ( .A(n23665), .B(n23751), .Z(n23669) );
  XOR U7537 ( .A(n23127), .B(n23213), .Z(n23131) );
  XOR U7538 ( .A(n22583), .B(n22669), .Z(n22587) );
  XOR U7539 ( .A(n22034), .B(n22120), .Z(n22038) );
  XOR U7540 ( .A(n21479), .B(n21565), .Z(n21483) );
  XOR U7541 ( .A(n20917), .B(n21003), .Z(n20921) );
  XOR U7542 ( .A(n20350), .B(n20436), .Z(n20354) );
  XOR U7543 ( .A(n19777), .B(n19863), .Z(n19781) );
  XOR U7544 ( .A(n19198), .B(n19284), .Z(n19202) );
  XOR U7545 ( .A(n3301), .B(n3472), .Z(n3305) );
  XOR U7546 ( .A(n1815), .B(n2010), .Z(n1819) );
  XOR U7547 ( .A(n1770), .B(n2019), .Z(n1774) );
  XOR U7548 ( .A(n17922), .B(n18003), .Z(n17926) );
  XOR U7549 ( .A(n4040), .B(n4193), .Z(n4044) );
  XOR U7550 ( .A(n1800), .B(n2013), .Z(n1804) );
  XOR U7551 ( .A(n3331), .B(n3466), .Z(n3335) );
  XOR U7552 ( .A(n1845), .B(n2004), .Z(n1849) );
  XOR U7553 ( .A(n17329), .B(n17404), .Z(n17333) );
  XOR U7554 ( .A(n16115), .B(n16190), .Z(n16119) );
  XOR U7555 ( .A(n14877), .B(n14952), .Z(n14881) );
  XOR U7556 ( .A(n13615), .B(n13690), .Z(n13619) );
  XOR U7557 ( .A(n12327), .B(n12404), .Z(n12331) );
  XOR U7558 ( .A(n11017), .B(n11092), .Z(n11021) );
  XOR U7559 ( .A(n9683), .B(n9758), .Z(n9687) );
  XOR U7560 ( .A(n8325), .B(n8400), .Z(n8329) );
  XOR U7561 ( .A(n6943), .B(n7018), .Z(n6947) );
  XOR U7562 ( .A(n5535), .B(n5612), .Z(n5539) );
  XOR U7563 ( .A(n4070), .B(n4187), .Z(n4074) );
  XOR U7564 ( .A(n2641), .B(n2728), .Z(n2645) );
  XOR U7565 ( .A(n47019), .B(n47087), .Z(n47023) );
  XOR U7566 ( .A(n46944), .B(n47012), .Z(n46948) );
  XOR U7567 ( .A(n46863), .B(n46931), .Z(n46867) );
  XOR U7568 ( .A(n46776), .B(n46844), .Z(n46780) );
  XOR U7569 ( .A(n46683), .B(n46751), .Z(n46687) );
  XOR U7570 ( .A(n46479), .B(n46547), .Z(n46483) );
  XOR U7571 ( .A(n46368), .B(n46436), .Z(n46372) );
  XOR U7572 ( .A(n46251), .B(n46319), .Z(n46255) );
  XOR U7573 ( .A(n46128), .B(n46196), .Z(n46132) );
  XOR U7574 ( .A(n45999), .B(n46067), .Z(n46003) );
  XOR U7575 ( .A(n45864), .B(n45932), .Z(n45868) );
  XOR U7576 ( .A(n45723), .B(n45791), .Z(n45727) );
  XOR U7577 ( .A(n45576), .B(n45644), .Z(n45580) );
  XOR U7578 ( .A(n45423), .B(n45491), .Z(n45427) );
  XOR U7579 ( .A(n45264), .B(n45332), .Z(n45268) );
  XOR U7580 ( .A(n45099), .B(n45167), .Z(n45103) );
  XOR U7581 ( .A(n44928), .B(n44996), .Z(n44932) );
  XOR U7582 ( .A(n44751), .B(n44819), .Z(n44755) );
  XOR U7583 ( .A(n44568), .B(n44636), .Z(n44572) );
  XOR U7584 ( .A(n44379), .B(n44447), .Z(n44383) );
  XOR U7585 ( .A(n44184), .B(n44252), .Z(n44188) );
  XOR U7586 ( .A(n43983), .B(n44051), .Z(n43987) );
  XOR U7587 ( .A(n43776), .B(n43844), .Z(n43780) );
  XOR U7588 ( .A(n43563), .B(n43631), .Z(n43567) );
  XOR U7589 ( .A(n43344), .B(n43412), .Z(n43348) );
  XOR U7590 ( .A(n43119), .B(n43187), .Z(n43123) );
  XOR U7591 ( .A(n42888), .B(n42956), .Z(n42892) );
  XOR U7592 ( .A(n42651), .B(n42719), .Z(n42655) );
  XOR U7593 ( .A(n42408), .B(n42476), .Z(n42412) );
  XOR U7594 ( .A(n42159), .B(n42227), .Z(n42163) );
  XOR U7595 ( .A(n41904), .B(n41972), .Z(n41908) );
  XOR U7596 ( .A(n41643), .B(n41711), .Z(n41647) );
  XOR U7597 ( .A(n41376), .B(n41444), .Z(n41380) );
  XOR U7598 ( .A(n41103), .B(n41171), .Z(n41107) );
  XOR U7599 ( .A(n40824), .B(n40892), .Z(n40828) );
  XOR U7600 ( .A(n40539), .B(n40607), .Z(n40543) );
  XOR U7601 ( .A(n40248), .B(n40316), .Z(n40252) );
  XOR U7602 ( .A(n39951), .B(n40019), .Z(n39955) );
  XOR U7603 ( .A(n39648), .B(n39716), .Z(n39652) );
  XOR U7604 ( .A(n39339), .B(n39407), .Z(n39343) );
  XOR U7605 ( .A(n39024), .B(n39092), .Z(n39028) );
  XOR U7606 ( .A(n38703), .B(n38771), .Z(n38707) );
  XOR U7607 ( .A(n38376), .B(n38444), .Z(n38380) );
  XOR U7608 ( .A(n38043), .B(n38111), .Z(n38047) );
  XOR U7609 ( .A(n37704), .B(n37772), .Z(n37708) );
  XOR U7610 ( .A(n37359), .B(n37427), .Z(n37363) );
  XOR U7611 ( .A(n37008), .B(n37076), .Z(n37012) );
  XOR U7612 ( .A(n36651), .B(n36719), .Z(n36655) );
  XOR U7613 ( .A(n36288), .B(n36356), .Z(n36292) );
  XOR U7614 ( .A(n35919), .B(n35987), .Z(n35923) );
  XOR U7615 ( .A(n35544), .B(n35612), .Z(n35548) );
  XOR U7616 ( .A(n35163), .B(n35231), .Z(n35167) );
  XOR U7617 ( .A(n34776), .B(n34844), .Z(n34780) );
  XOR U7618 ( .A(n34383), .B(n34451), .Z(n34387) );
  XOR U7619 ( .A(n33984), .B(n34052), .Z(n33988) );
  XOR U7620 ( .A(n33579), .B(n33647), .Z(n33583) );
  XOR U7621 ( .A(n33168), .B(n33236), .Z(n33172) );
  XOR U7622 ( .A(n32751), .B(n32819), .Z(n32755) );
  XOR U7623 ( .A(n32328), .B(n32396), .Z(n32332) );
  XOR U7624 ( .A(n31899), .B(n31967), .Z(n31903) );
  XOR U7625 ( .A(n31464), .B(n31532), .Z(n31468) );
  XOR U7626 ( .A(n31023), .B(n31091), .Z(n31027) );
  XOR U7627 ( .A(n30576), .B(n30644), .Z(n30580) );
  XOR U7628 ( .A(n30123), .B(n30191), .Z(n30127) );
  XOR U7629 ( .A(n29664), .B(n29732), .Z(n29668) );
  XOR U7630 ( .A(n29199), .B(n29267), .Z(n29203) );
  XOR U7631 ( .A(n28728), .B(n28796), .Z(n28732) );
  XOR U7632 ( .A(n28251), .B(n28319), .Z(n28255) );
  XOR U7633 ( .A(n27768), .B(n27836), .Z(n27772) );
  XOR U7634 ( .A(n27279), .B(n27347), .Z(n27283) );
  XOR U7635 ( .A(n26782), .B(n26850), .Z(n26786) );
  XOR U7636 ( .A(n26281), .B(n26349), .Z(n26285) );
  XOR U7637 ( .A(n25773), .B(n25841), .Z(n25777) );
  XOR U7638 ( .A(n25259), .B(n25327), .Z(n25263) );
  XOR U7639 ( .A(n24736), .B(n24804), .Z(n24740) );
  XOR U7640 ( .A(n24211), .B(n24279), .Z(n24215) );
  XOR U7641 ( .A(n23680), .B(n23748), .Z(n23684) );
  XOR U7642 ( .A(n23142), .B(n23210), .Z(n23146) );
  XOR U7643 ( .A(n22598), .B(n22666), .Z(n22602) );
  XOR U7644 ( .A(n22049), .B(n22117), .Z(n22053) );
  XOR U7645 ( .A(n21494), .B(n21562), .Z(n21498) );
  XOR U7646 ( .A(n20932), .B(n21000), .Z(n20936) );
  XOR U7647 ( .A(n20365), .B(n20433), .Z(n20369) );
  XOR U7648 ( .A(n19792), .B(n19860), .Z(n19796) );
  XOR U7649 ( .A(n19213), .B(n19281), .Z(n19217) );
  XOR U7650 ( .A(n3361), .B(n3460), .Z(n3365) );
  XOR U7651 ( .A(n1875), .B(n1998), .Z(n1879) );
  XOR U7652 ( .A(n1830), .B(n2007), .Z(n1834) );
  XOR U7653 ( .A(n4100), .B(n4181), .Z(n4104) );
  XOR U7654 ( .A(n1860), .B(n2001), .Z(n1864) );
  XOR U7655 ( .A(n17942), .B(n17999), .Z(n17946) );
  XOR U7656 ( .A(n16740), .B(n16797), .Z(n16744) );
  XOR U7657 ( .A(n14892), .B(n14949), .Z(n14896) );
  XOR U7658 ( .A(n13630), .B(n13687), .Z(n13634) );
  XOR U7659 ( .A(n12342), .B(n12401), .Z(n12346) );
  XOR U7660 ( .A(n11032), .B(n11089), .Z(n11036) );
  XOR U7661 ( .A(n9698), .B(n9755), .Z(n9702) );
  XOR U7662 ( .A(n8340), .B(n8397), .Z(n8344) );
  XOR U7663 ( .A(n6958), .B(n7015), .Z(n6962) );
  XOR U7664 ( .A(n5550), .B(n5609), .Z(n5554) );
  XOR U7665 ( .A(n4120), .B(n4177), .Z(n4124) );
  XOR U7666 ( .A(n1930), .B(n1987), .Z(n1934) );
  XOR U7667 ( .A(n1910), .B(n1991), .Z(n1914) );
  XOR U7668 ( .A(n47222), .B(n47272), .Z(n47226) );
  XOR U7669 ( .A(n47166), .B(n47215), .Z(n47170) );
  XOR U7670 ( .A(n47103), .B(n47153), .Z(n47107) );
  XOR U7671 ( .A(n47034), .B(n47084), .Z(n47038) );
  XOR U7672 ( .A(n46959), .B(n47009), .Z(n46963) );
  XOR U7673 ( .A(n46791), .B(n46841), .Z(n46795) );
  XOR U7674 ( .A(n46698), .B(n46748), .Z(n46702) );
  XOR U7675 ( .A(n46599), .B(n46649), .Z(n46603) );
  XOR U7676 ( .A(n46494), .B(n46544), .Z(n46498) );
  XOR U7677 ( .A(n46383), .B(n46433), .Z(n46387) );
  XOR U7678 ( .A(n46266), .B(n46316), .Z(n46270) );
  XOR U7679 ( .A(n46143), .B(n46193), .Z(n46147) );
  XOR U7680 ( .A(n46014), .B(n46064), .Z(n46018) );
  XOR U7681 ( .A(n45879), .B(n45929), .Z(n45883) );
  XOR U7682 ( .A(n45738), .B(n45788), .Z(n45742) );
  XOR U7683 ( .A(n45591), .B(n45641), .Z(n45595) );
  XOR U7684 ( .A(n45438), .B(n45488), .Z(n45442) );
  XOR U7685 ( .A(n45279), .B(n45329), .Z(n45283) );
  XOR U7686 ( .A(n45114), .B(n45164), .Z(n45118) );
  XOR U7687 ( .A(n44943), .B(n44993), .Z(n44947) );
  XOR U7688 ( .A(n44766), .B(n44816), .Z(n44770) );
  XOR U7689 ( .A(n44583), .B(n44633), .Z(n44587) );
  XOR U7690 ( .A(n44394), .B(n44444), .Z(n44398) );
  XOR U7691 ( .A(n44199), .B(n44249), .Z(n44203) );
  XOR U7692 ( .A(n43998), .B(n44048), .Z(n44002) );
  XOR U7693 ( .A(n43791), .B(n43841), .Z(n43795) );
  XOR U7694 ( .A(n43578), .B(n43628), .Z(n43582) );
  XOR U7695 ( .A(n43359), .B(n43409), .Z(n43363) );
  XOR U7696 ( .A(n43134), .B(n43184), .Z(n43138) );
  XOR U7697 ( .A(n42903), .B(n42953), .Z(n42907) );
  XOR U7698 ( .A(n42666), .B(n42716), .Z(n42670) );
  XOR U7699 ( .A(n42423), .B(n42473), .Z(n42427) );
  XOR U7700 ( .A(n42174), .B(n42224), .Z(n42178) );
  XOR U7701 ( .A(n41919), .B(n41969), .Z(n41923) );
  XOR U7702 ( .A(n41658), .B(n41708), .Z(n41662) );
  XOR U7703 ( .A(n41391), .B(n41441), .Z(n41395) );
  XOR U7704 ( .A(n41118), .B(n41168), .Z(n41122) );
  XOR U7705 ( .A(n40839), .B(n40889), .Z(n40843) );
  XOR U7706 ( .A(n40554), .B(n40604), .Z(n40558) );
  XOR U7707 ( .A(n40263), .B(n40313), .Z(n40267) );
  XOR U7708 ( .A(n39966), .B(n40016), .Z(n39970) );
  XOR U7709 ( .A(n39663), .B(n39713), .Z(n39667) );
  XOR U7710 ( .A(n39354), .B(n39404), .Z(n39358) );
  XOR U7711 ( .A(n39039), .B(n39089), .Z(n39043) );
  XOR U7712 ( .A(n38718), .B(n38768), .Z(n38722) );
  XOR U7713 ( .A(n38391), .B(n38441), .Z(n38395) );
  XOR U7714 ( .A(n38058), .B(n38108), .Z(n38062) );
  XOR U7715 ( .A(n37719), .B(n37769), .Z(n37723) );
  XOR U7716 ( .A(n37374), .B(n37424), .Z(n37378) );
  XOR U7717 ( .A(n37023), .B(n37073), .Z(n37027) );
  XOR U7718 ( .A(n36666), .B(n36716), .Z(n36670) );
  XOR U7719 ( .A(n36303), .B(n36353), .Z(n36307) );
  XOR U7720 ( .A(n35934), .B(n35984), .Z(n35938) );
  XOR U7721 ( .A(n35559), .B(n35609), .Z(n35563) );
  XOR U7722 ( .A(n35178), .B(n35228), .Z(n35182) );
  XOR U7723 ( .A(n34791), .B(n34841), .Z(n34795) );
  XOR U7724 ( .A(n34398), .B(n34448), .Z(n34402) );
  XOR U7725 ( .A(n33999), .B(n34049), .Z(n34003) );
  XOR U7726 ( .A(n33594), .B(n33644), .Z(n33598) );
  XOR U7727 ( .A(n33183), .B(n33233), .Z(n33187) );
  XOR U7728 ( .A(n32766), .B(n32816), .Z(n32770) );
  XOR U7729 ( .A(n32343), .B(n32393), .Z(n32347) );
  XOR U7730 ( .A(n31914), .B(n31964), .Z(n31918) );
  XOR U7731 ( .A(n31479), .B(n31529), .Z(n31483) );
  XOR U7732 ( .A(n31038), .B(n31088), .Z(n31042) );
  XOR U7733 ( .A(n30591), .B(n30641), .Z(n30595) );
  XOR U7734 ( .A(n30138), .B(n30188), .Z(n30142) );
  XOR U7735 ( .A(n29679), .B(n29729), .Z(n29683) );
  XOR U7736 ( .A(n29214), .B(n29264), .Z(n29218) );
  XOR U7737 ( .A(n28743), .B(n28793), .Z(n28747) );
  XOR U7738 ( .A(n28266), .B(n28316), .Z(n28270) );
  XOR U7739 ( .A(n27783), .B(n27833), .Z(n27787) );
  XOR U7740 ( .A(n27294), .B(n27344), .Z(n27298) );
  XOR U7741 ( .A(n26797), .B(n26847), .Z(n26801) );
  XOR U7742 ( .A(n26296), .B(n26346), .Z(n26300) );
  XOR U7743 ( .A(n25788), .B(n25838), .Z(n25792) );
  XOR U7744 ( .A(n25274), .B(n25324), .Z(n25278) );
  XOR U7745 ( .A(n24751), .B(n24801), .Z(n24755) );
  XOR U7746 ( .A(n24226), .B(n24276), .Z(n24230) );
  XOR U7747 ( .A(n23695), .B(n23745), .Z(n23699) );
  XOR U7748 ( .A(n23157), .B(n23207), .Z(n23161) );
  XOR U7749 ( .A(n22613), .B(n22663), .Z(n22617) );
  XOR U7750 ( .A(n22064), .B(n22114), .Z(n22068) );
  XOR U7751 ( .A(n21509), .B(n21559), .Z(n21513) );
  XOR U7752 ( .A(n20947), .B(n20997), .Z(n20951) );
  XOR U7753 ( .A(n20380), .B(n20430), .Z(n20384) );
  XOR U7754 ( .A(n19807), .B(n19857), .Z(n19811) );
  XOR U7755 ( .A(n19228), .B(n19278), .Z(n19232) );
  XOR U7756 ( .A(n16135), .B(n16186), .Z(n16139) );
  XOR U7757 ( .A(n1890), .B(n1995), .Z(n1894) );
  XOR U7758 ( .A(n2661), .B(n2724), .Z(n2665) );
  XOR U7759 ( .A(n17957), .B(n17996), .Z(n17961) );
  XOR U7760 ( .A(n15529), .B(n15568), .Z(n15533) );
  XOR U7761 ( .A(n14279), .B(n14318), .Z(n14283) );
  XOR U7762 ( .A(n13005), .B(n13044), .Z(n13009) );
  XOR U7763 ( .A(n11705), .B(n11744), .Z(n11709) );
  XOR U7764 ( .A(n10383), .B(n10422), .Z(n10387) );
  XOR U7765 ( .A(n9037), .B(n9076), .Z(n9041) );
  XOR U7766 ( .A(n7667), .B(n7706), .Z(n7671) );
  XOR U7767 ( .A(n6273), .B(n6312), .Z(n6277) );
  XOR U7768 ( .A(n4853), .B(n4892), .Z(n4857) );
  XOR U7769 ( .A(n3411), .B(n3450), .Z(n3415) );
  XOR U7770 ( .A(n1945), .B(n1984), .Z(n1949) );
  XOR U7771 ( .A(n47372), .B(n47404), .Z(n47376) );
  XOR U7772 ( .A(n47333), .B(n47365), .Z(n47337) );
  XOR U7773 ( .A(n47288), .B(n47320), .Z(n47292) );
  XOR U7774 ( .A(n47237), .B(n47269), .Z(n47241) );
  XOR U7775 ( .A(n47181), .B(n47212), .Z(n47185) );
  XOR U7776 ( .A(n47049), .B(n47081), .Z(n47053) );
  XOR U7777 ( .A(n46974), .B(n47006), .Z(n46978) );
  XOR U7778 ( .A(n46893), .B(n46925), .Z(n46897) );
  XOR U7779 ( .A(n46806), .B(n46838), .Z(n46810) );
  XOR U7780 ( .A(n46713), .B(n46745), .Z(n46717) );
  XOR U7781 ( .A(n46614), .B(n46646), .Z(n46618) );
  XOR U7782 ( .A(n46509), .B(n46541), .Z(n46513) );
  XOR U7783 ( .A(n46398), .B(n46430), .Z(n46402) );
  XOR U7784 ( .A(n46281), .B(n46313), .Z(n46285) );
  XOR U7785 ( .A(n46158), .B(n46190), .Z(n46162) );
  XOR U7786 ( .A(n46029), .B(n46061), .Z(n46033) );
  XOR U7787 ( .A(n45894), .B(n45926), .Z(n45898) );
  XOR U7788 ( .A(n45753), .B(n45785), .Z(n45757) );
  XOR U7789 ( .A(n45606), .B(n45638), .Z(n45610) );
  XOR U7790 ( .A(n45453), .B(n45485), .Z(n45457) );
  XOR U7791 ( .A(n45294), .B(n45326), .Z(n45298) );
  XOR U7792 ( .A(n45129), .B(n45161), .Z(n45133) );
  XOR U7793 ( .A(n44958), .B(n44990), .Z(n44962) );
  XOR U7794 ( .A(n44781), .B(n44813), .Z(n44785) );
  XOR U7795 ( .A(n44598), .B(n44630), .Z(n44602) );
  XOR U7796 ( .A(n44409), .B(n44441), .Z(n44413) );
  XOR U7797 ( .A(n44214), .B(n44246), .Z(n44218) );
  XOR U7798 ( .A(n44013), .B(n44045), .Z(n44017) );
  XOR U7799 ( .A(n43806), .B(n43838), .Z(n43810) );
  XOR U7800 ( .A(n43593), .B(n43625), .Z(n43597) );
  XOR U7801 ( .A(n43374), .B(n43406), .Z(n43378) );
  XOR U7802 ( .A(n43149), .B(n43181), .Z(n43153) );
  XOR U7803 ( .A(n42918), .B(n42950), .Z(n42922) );
  XOR U7804 ( .A(n42681), .B(n42713), .Z(n42685) );
  XOR U7805 ( .A(n42438), .B(n42470), .Z(n42442) );
  XOR U7806 ( .A(n42189), .B(n42221), .Z(n42193) );
  XOR U7807 ( .A(n41934), .B(n41966), .Z(n41938) );
  XOR U7808 ( .A(n41673), .B(n41705), .Z(n41677) );
  XOR U7809 ( .A(n41406), .B(n41438), .Z(n41410) );
  XOR U7810 ( .A(n41133), .B(n41165), .Z(n41137) );
  XOR U7811 ( .A(n40854), .B(n40886), .Z(n40858) );
  XOR U7812 ( .A(n40569), .B(n40601), .Z(n40573) );
  XOR U7813 ( .A(n40278), .B(n40310), .Z(n40282) );
  XOR U7814 ( .A(n39981), .B(n40013), .Z(n39985) );
  XOR U7815 ( .A(n39678), .B(n39710), .Z(n39682) );
  XOR U7816 ( .A(n39369), .B(n39401), .Z(n39373) );
  XOR U7817 ( .A(n39054), .B(n39086), .Z(n39058) );
  XOR U7818 ( .A(n38733), .B(n38765), .Z(n38737) );
  XOR U7819 ( .A(n38406), .B(n38438), .Z(n38410) );
  XOR U7820 ( .A(n38073), .B(n38105), .Z(n38077) );
  XOR U7821 ( .A(n37734), .B(n37766), .Z(n37738) );
  XOR U7822 ( .A(n37389), .B(n37421), .Z(n37393) );
  XOR U7823 ( .A(n37038), .B(n37070), .Z(n37042) );
  XOR U7824 ( .A(n36681), .B(n36713), .Z(n36685) );
  XOR U7825 ( .A(n36318), .B(n36350), .Z(n36322) );
  XOR U7826 ( .A(n35949), .B(n35981), .Z(n35953) );
  XOR U7827 ( .A(n35574), .B(n35606), .Z(n35578) );
  XOR U7828 ( .A(n35193), .B(n35225), .Z(n35197) );
  XOR U7829 ( .A(n34806), .B(n34838), .Z(n34810) );
  XOR U7830 ( .A(n34413), .B(n34445), .Z(n34417) );
  XOR U7831 ( .A(n34014), .B(n34046), .Z(n34018) );
  XOR U7832 ( .A(n33609), .B(n33641), .Z(n33613) );
  XOR U7833 ( .A(n33198), .B(n33230), .Z(n33202) );
  XOR U7834 ( .A(n32781), .B(n32813), .Z(n32785) );
  XOR U7835 ( .A(n32358), .B(n32390), .Z(n32362) );
  XOR U7836 ( .A(n31929), .B(n31961), .Z(n31933) );
  XOR U7837 ( .A(n31494), .B(n31526), .Z(n31498) );
  XOR U7838 ( .A(n31053), .B(n31085), .Z(n31057) );
  XOR U7839 ( .A(n30606), .B(n30638), .Z(n30610) );
  XOR U7840 ( .A(n30153), .B(n30185), .Z(n30157) );
  XOR U7841 ( .A(n29694), .B(n29726), .Z(n29698) );
  XOR U7842 ( .A(n29229), .B(n29261), .Z(n29233) );
  XOR U7843 ( .A(n28758), .B(n28790), .Z(n28762) );
  XOR U7844 ( .A(n28281), .B(n28313), .Z(n28285) );
  XOR U7845 ( .A(n27798), .B(n27830), .Z(n27802) );
  XOR U7846 ( .A(n27309), .B(n27341), .Z(n27313) );
  XOR U7847 ( .A(n26812), .B(n26844), .Z(n26816) );
  XOR U7848 ( .A(n26311), .B(n26343), .Z(n26315) );
  XOR U7849 ( .A(n25803), .B(n25835), .Z(n25807) );
  XOR U7850 ( .A(n25289), .B(n25321), .Z(n25293) );
  XOR U7851 ( .A(n24766), .B(n24798), .Z(n24770) );
  XOR U7852 ( .A(n24241), .B(n24273), .Z(n24245) );
  XOR U7853 ( .A(n23710), .B(n23742), .Z(n23714) );
  XOR U7854 ( .A(n23172), .B(n23204), .Z(n23176) );
  XOR U7855 ( .A(n22628), .B(n22660), .Z(n22632) );
  XOR U7856 ( .A(n22079), .B(n22111), .Z(n22083) );
  XOR U7857 ( .A(n21524), .B(n21556), .Z(n21528) );
  XOR U7858 ( .A(n20962), .B(n20994), .Z(n20966) );
  XOR U7859 ( .A(n20395), .B(n20427), .Z(n20399) );
  XOR U7860 ( .A(n19822), .B(n19854), .Z(n19826) );
  XOR U7861 ( .A(n19243), .B(n19275), .Z(n19247) );
  XOR U7862 ( .A(n17364), .B(n17397), .Z(n17368) );
  XOR U7863 ( .A(n16770), .B(n16791), .Z(n16774) );
  XOR U7864 ( .A(n15544), .B(n15565), .Z(n15548) );
  XOR U7865 ( .A(n14294), .B(n14315), .Z(n14298) );
  XOR U7866 ( .A(n13020), .B(n13041), .Z(n13024) );
  XOR U7867 ( .A(n11720), .B(n11741), .Z(n11724) );
  XOR U7868 ( .A(n10398), .B(n10419), .Z(n10402) );
  XOR U7869 ( .A(n9052), .B(n9073), .Z(n9056) );
  XOR U7870 ( .A(n7682), .B(n7703), .Z(n7686) );
  XOR U7871 ( .A(n6288), .B(n6309), .Z(n6292) );
  XOR U7872 ( .A(n4868), .B(n4889), .Z(n4872) );
  XOR U7873 ( .A(n3426), .B(n3447), .Z(n3430) );
  XOR U7874 ( .A(n1960), .B(n1981), .Z(n1964) );
  XNOR U7875 ( .A(n47472), .B(n47471), .Z(n47458) );
  XOR U7876 ( .A(n47447), .B(n47452), .Z(n47430) );
  XNOR U7877 ( .A(n47424), .B(n47423), .Z(n47398) );
  XNOR U7878 ( .A(n47391), .B(n47390), .Z(n47359) );
  XOR U7879 ( .A(n47348), .B(n47353), .Z(n47313) );
  XOR U7880 ( .A(n47252), .B(n47257), .Z(n47205) );
  XOR U7881 ( .A(n47196), .B(n47201), .Z(n47143) );
  XNOR U7882 ( .A(n47137), .B(n47136), .Z(n47075) );
  XNOR U7883 ( .A(n47068), .B(n47067), .Z(n47000) );
  XOR U7884 ( .A(n46989), .B(n46994), .Z(n46918) );
  XNOR U7885 ( .A(n46912), .B(n46911), .Z(n46832) );
  XNOR U7886 ( .A(n46825), .B(n46824), .Z(n46739) );
  XOR U7887 ( .A(n46728), .B(n46733), .Z(n46639) );
  XNOR U7888 ( .A(n46633), .B(n46632), .Z(n46535) );
  XNOR U7889 ( .A(n46528), .B(n46527), .Z(n46424) );
  XOR U7890 ( .A(n46413), .B(n46418), .Z(n46306) );
  XNOR U7891 ( .A(n46300), .B(n46299), .Z(n46184) );
  XNOR U7892 ( .A(n46177), .B(n46176), .Z(n46055) );
  XOR U7893 ( .A(n46044), .B(n46049), .Z(n45919) );
  XNOR U7894 ( .A(n45913), .B(n45912), .Z(n45779) );
  XNOR U7895 ( .A(n45772), .B(n45771), .Z(n45632) );
  XOR U7896 ( .A(n45621), .B(n45626), .Z(n45478) );
  XNOR U7897 ( .A(n45472), .B(n45471), .Z(n45320) );
  XNOR U7898 ( .A(n45313), .B(n45312), .Z(n45155) );
  XOR U7899 ( .A(n45144), .B(n45149), .Z(n44983) );
  XNOR U7900 ( .A(n44977), .B(n44976), .Z(n44807) );
  XNOR U7901 ( .A(n44800), .B(n44799), .Z(n44624) );
  XOR U7902 ( .A(n44613), .B(n44618), .Z(n44434) );
  XNOR U7903 ( .A(n44428), .B(n44427), .Z(n44240) );
  XNOR U7904 ( .A(n44233), .B(n44232), .Z(n44039) );
  XOR U7905 ( .A(n44028), .B(n44033), .Z(n43831) );
  XNOR U7906 ( .A(n43825), .B(n43824), .Z(n43619) );
  XNOR U7907 ( .A(n43612), .B(n43611), .Z(n43400) );
  XOR U7908 ( .A(n43389), .B(n43394), .Z(n43174) );
  XNOR U7909 ( .A(n43168), .B(n43167), .Z(n42944) );
  XNOR U7910 ( .A(n42937), .B(n42936), .Z(n42707) );
  XOR U7911 ( .A(n42696), .B(n42701), .Z(n42463) );
  XNOR U7912 ( .A(n42457), .B(n42456), .Z(n42215) );
  XNOR U7913 ( .A(n42208), .B(n42207), .Z(n41960) );
  XOR U7914 ( .A(n41949), .B(n41954), .Z(n41698) );
  XNOR U7915 ( .A(n41692), .B(n41691), .Z(n41432) );
  XNOR U7916 ( .A(n41425), .B(n41424), .Z(n41159) );
  XOR U7917 ( .A(n41148), .B(n41153), .Z(n40879) );
  XNOR U7918 ( .A(n40873), .B(n40872), .Z(n40595) );
  XNOR U7919 ( .A(n40588), .B(n40587), .Z(n40304) );
  XOR U7920 ( .A(n40293), .B(n40298), .Z(n40006) );
  XNOR U7921 ( .A(n40000), .B(n39999), .Z(n39704) );
  XNOR U7922 ( .A(n39697), .B(n39696), .Z(n39395) );
  XOR U7923 ( .A(n39384), .B(n39389), .Z(n39079) );
  XNOR U7924 ( .A(n39073), .B(n39072), .Z(n38759) );
  XNOR U7925 ( .A(n38752), .B(n38751), .Z(n38432) );
  XOR U7926 ( .A(n38421), .B(n38426), .Z(n38098) );
  XNOR U7927 ( .A(n38092), .B(n38091), .Z(n37760) );
  XNOR U7928 ( .A(n37753), .B(n37752), .Z(n37415) );
  XOR U7929 ( .A(n37404), .B(n37409), .Z(n37063) );
  XNOR U7930 ( .A(n37057), .B(n37056), .Z(n36707) );
  XNOR U7931 ( .A(n36700), .B(n36699), .Z(n36344) );
  XOR U7932 ( .A(n36333), .B(n36338), .Z(n35974) );
  XNOR U7933 ( .A(n35968), .B(n35967), .Z(n35600) );
  XNOR U7934 ( .A(n35593), .B(n35592), .Z(n35219) );
  XOR U7935 ( .A(n35208), .B(n35213), .Z(n34831) );
  XNOR U7936 ( .A(n34825), .B(n34824), .Z(n34439) );
  XNOR U7937 ( .A(n34432), .B(n34431), .Z(n34040) );
  XOR U7938 ( .A(n34029), .B(n34034), .Z(n33634) );
  XNOR U7939 ( .A(n33628), .B(n33627), .Z(n33224) );
  XNOR U7940 ( .A(n33217), .B(n33216), .Z(n32807) );
  XOR U7941 ( .A(n32796), .B(n32801), .Z(n32383) );
  XNOR U7942 ( .A(n32377), .B(n32376), .Z(n31955) );
  XNOR U7943 ( .A(n31948), .B(n31947), .Z(n31520) );
  XOR U7944 ( .A(n31509), .B(n31514), .Z(n31078) );
  XNOR U7945 ( .A(n31072), .B(n31071), .Z(n30632) );
  XNOR U7946 ( .A(n30625), .B(n30624), .Z(n30179) );
  XOR U7947 ( .A(n30168), .B(n30173), .Z(n29719) );
  XNOR U7948 ( .A(n29713), .B(n29712), .Z(n29255) );
  XNOR U7949 ( .A(n29248), .B(n29247), .Z(n28784) );
  XOR U7950 ( .A(n28773), .B(n28778), .Z(n28306) );
  XNOR U7951 ( .A(n28300), .B(n28299), .Z(n27824) );
  XNOR U7952 ( .A(n27817), .B(n27816), .Z(n27335) );
  XOR U7953 ( .A(n27324), .B(n27329), .Z(n26837) );
  XNOR U7954 ( .A(n26831), .B(n26830), .Z(n26337) );
  XNOR U7955 ( .A(n26330), .B(n26329), .Z(n25829) );
  XOR U7956 ( .A(n25818), .B(n25823), .Z(n25314) );
  XNOR U7957 ( .A(n25308), .B(n25307), .Z(n24792) );
  XNOR U7958 ( .A(n24785), .B(n24784), .Z(n24267) );
  XOR U7959 ( .A(n24256), .B(n24261), .Z(n23735) );
  XNOR U7960 ( .A(n23729), .B(n23728), .Z(n23198) );
  XNOR U7961 ( .A(n23191), .B(n23190), .Z(n22654) );
  XOR U7962 ( .A(n22643), .B(n22648), .Z(n22104) );
  XNOR U7963 ( .A(n22098), .B(n22097), .Z(n21550) );
  XNOR U7964 ( .A(n21543), .B(n21542), .Z(n20988) );
  XOR U7965 ( .A(n20977), .B(n20982), .Z(n20420) );
  XNOR U7966 ( .A(n20414), .B(n20413), .Z(n19848) );
  XNOR U7967 ( .A(n19841), .B(n19840), .Z(n19269) );
  XNOR U7968 ( .A(n19262), .B(n19261), .Z(n18589) );
  XOR U7969 ( .A(n17977), .B(n17992), .Z(n17986) );
  XNOR U7970 ( .A(n26930), .B(n26430), .Z(n26432) );
  XNOR U7971 ( .A(n29340), .B(n28872), .Z(n28874) );
  XNOR U7972 ( .A(n28875), .B(n28401), .Z(n28403) );
  XNOR U7973 ( .A(n28404), .B(n27924), .Z(n27926) );
  XNOR U7974 ( .A(n26453), .B(n25949), .Z(n25951) );
  XNOR U7975 ( .A(n26433), .B(n25929), .Z(n25931) );
  XNOR U7976 ( .A(n27937), .B(n27451), .Z(n27453) );
  XNOR U7977 ( .A(n26945), .B(n26445), .Z(n26447) );
  XNOR U7978 ( .A(n26438), .B(n25934), .Z(n25936) );
  XNOR U7979 ( .A(n25409), .B(n24891), .Z(n24893) );
  XNOR U7980 ( .A(n30714), .B(n30264), .Z(n30266) );
  XNOR U7981 ( .A(n30267), .B(n29811), .Z(n29813) );
  XNOR U7982 ( .A(n29814), .B(n29352), .Z(n29354) );
  XNOR U7983 ( .A(n29355), .B(n28887), .Z(n28889) );
  XNOR U7984 ( .A(n28890), .B(n28416), .Z(n28418) );
  XNOR U7985 ( .A(n27942), .B(n27456), .Z(n27458) );
  XNOR U7986 ( .A(n26463), .B(n25959), .Z(n25961) );
  XNOR U7987 ( .A(n25439), .B(n24921), .Z(n24923) );
  XNOR U7988 ( .A(n24914), .B(n24389), .Z(n24391) );
  XNOR U7989 ( .A(n26448), .B(n25944), .Z(n25946) );
  XNOR U7990 ( .A(n24894), .B(n24369), .Z(n24371) );
  XNOR U7991 ( .A(n29365), .B(n28897), .Z(n28899) );
  XOR U7992 ( .A(n25448), .B(n25907), .Z(n25452) );
  XNOR U7993 ( .A(n25424), .B(n24906), .Z(n24908) );
  XNOR U7994 ( .A(n24899), .B(n24374), .Z(n24376) );
  XNOR U7995 ( .A(n23832), .B(n23298), .Z(n23300) );
  XNOR U7996 ( .A(n24944), .B(n24419), .Z(n24421) );
  XNOR U7997 ( .A(n32034), .B(n31602), .Z(n31604) );
  XNOR U7998 ( .A(n31605), .B(n31167), .Z(n31169) );
  XNOR U7999 ( .A(n31170), .B(n30726), .Z(n30728) );
  XNOR U8000 ( .A(n30729), .B(n30279), .Z(n30281) );
  XNOR U8001 ( .A(n30282), .B(n29826), .Z(n29828) );
  XNOR U8002 ( .A(n29370), .B(n28902), .Z(n28904) );
  XNOR U8003 ( .A(n28905), .B(n28431), .Z(n28433) );
  XNOR U8004 ( .A(n28434), .B(n27954), .Z(n27956) );
  XNOR U8005 ( .A(n27957), .B(n27471), .Z(n27473) );
  XNOR U8006 ( .A(n27474), .B(n26982), .Z(n26984) );
  XNOR U8007 ( .A(n26985), .B(n26485), .Z(n26487) );
  XNOR U8008 ( .A(n26488), .B(n25984), .Z(n25986) );
  XNOR U8009 ( .A(n24924), .B(n24399), .Z(n24401) );
  XNOR U8010 ( .A(n25972), .B(n25461), .Z(n25463) );
  XNOR U8011 ( .A(n25454), .B(n24936), .Z(n24938) );
  XNOR U8012 ( .A(n23862), .B(n23328), .Z(n23330) );
  XNOR U8013 ( .A(n23321), .B(n22780), .Z(n22782) );
  XNOR U8014 ( .A(n24909), .B(n24384), .Z(n24386) );
  XNOR U8015 ( .A(n23301), .B(n22760), .Z(n22762) );
  XNOR U8016 ( .A(n24954), .B(n24429), .Z(n24431) );
  XNOR U8017 ( .A(n30739), .B(n30289), .Z(n30291) );
  XOR U8018 ( .A(n23871), .B(n24347), .Z(n23875) );
  XNOR U8019 ( .A(n23847), .B(n23313), .Z(n23315) );
  XNOR U8020 ( .A(n23306), .B(n22765), .Z(n22767) );
  XNOR U8021 ( .A(n22204), .B(n21652), .Z(n21654) );
  XNOR U8022 ( .A(n24959), .B(n24434), .Z(n24436) );
  XNOR U8023 ( .A(n23892), .B(n23358), .Z(n23360) );
  XNOR U8024 ( .A(n23351), .B(n22810), .Z(n22812) );
  XNOR U8025 ( .A(n33300), .B(n32886), .Z(n32888) );
  XNOR U8026 ( .A(n32889), .B(n32469), .Z(n32471) );
  XNOR U8027 ( .A(n32472), .B(n32046), .Z(n32048) );
  XNOR U8028 ( .A(n32049), .B(n31617), .Z(n31619) );
  XNOR U8029 ( .A(n31620), .B(n31182), .Z(n31184) );
  XNOR U8030 ( .A(n30744), .B(n30294), .Z(n30296) );
  XNOR U8031 ( .A(n30297), .B(n29841), .Z(n29843) );
  XNOR U8032 ( .A(n29844), .B(n29382), .Z(n29384) );
  XNOR U8033 ( .A(n29385), .B(n28917), .Z(n28919) );
  XNOR U8034 ( .A(n28920), .B(n28446), .Z(n28448) );
  XNOR U8035 ( .A(n28449), .B(n27969), .Z(n27971) );
  XNOR U8036 ( .A(n27972), .B(n27486), .Z(n27488) );
  XNOR U8037 ( .A(n27489), .B(n26997), .Z(n26999) );
  XNOR U8038 ( .A(n27000), .B(n26500), .Z(n26502) );
  XNOR U8039 ( .A(n26503), .B(n25999), .Z(n26001) );
  XNOR U8040 ( .A(n25494), .B(n24976), .Z(n24978) );
  XNOR U8041 ( .A(n24452), .B(n23924), .Z(n23926) );
  XNOR U8042 ( .A(n23331), .B(n22790), .Z(n22792) );
  XNOR U8043 ( .A(n23381), .B(n22840), .Z(n22842) );
  XNOR U8044 ( .A(n24412), .B(n23884), .Z(n23886) );
  XNOR U8045 ( .A(n23877), .B(n23343), .Z(n23345) );
  XNOR U8046 ( .A(n22234), .B(n21682), .Z(n21684) );
  XNOR U8047 ( .A(n21675), .B(n21117), .Z(n21119) );
  XNOR U8048 ( .A(n23316), .B(n22775), .Z(n22777) );
  XNOR U8049 ( .A(n21655), .B(n21097), .Z(n21099) );
  XNOR U8050 ( .A(n24969), .B(n24444), .Z(n24446) );
  XNOR U8051 ( .A(n23361), .B(n22820), .Z(n22822) );
  XNOR U8052 ( .A(n32059), .B(n31627), .Z(n31629) );
  XNOR U8053 ( .A(n23927), .B(n23393), .Z(n23395) );
  XOR U8054 ( .A(n22243), .B(n22738), .Z(n22247) );
  XNOR U8055 ( .A(n22219), .B(n21667), .Z(n21669) );
  XNOR U8056 ( .A(n21660), .B(n21102), .Z(n21104) );
  XNOR U8057 ( .A(n20523), .B(n19953), .Z(n19955) );
  XNOR U8058 ( .A(n23907), .B(n23373), .Z(n23375) );
  XNOR U8059 ( .A(n23366), .B(n22825), .Z(n22827) );
  XNOR U8060 ( .A(n22264), .B(n21712), .Z(n21714) );
  XNOR U8061 ( .A(n21705), .B(n21147), .Z(n21149) );
  XNOR U8062 ( .A(n34512), .B(n34116), .Z(n34118) );
  XNOR U8063 ( .A(n34119), .B(n33717), .Z(n33719) );
  XNOR U8064 ( .A(n33720), .B(n33312), .Z(n33314) );
  XNOR U8065 ( .A(n33315), .B(n32901), .Z(n32903) );
  XNOR U8066 ( .A(n32904), .B(n32484), .Z(n32486) );
  XNOR U8067 ( .A(n32064), .B(n31632), .Z(n31634) );
  XNOR U8068 ( .A(n31635), .B(n31197), .Z(n31199) );
  XNOR U8069 ( .A(n31200), .B(n30756), .Z(n30758) );
  XNOR U8070 ( .A(n30759), .B(n30309), .Z(n30311) );
  XNOR U8071 ( .A(n30312), .B(n29856), .Z(n29858) );
  XNOR U8072 ( .A(n29859), .B(n29397), .Z(n29399) );
  XNOR U8073 ( .A(n29400), .B(n28932), .Z(n28934) );
  XNOR U8074 ( .A(n28935), .B(n28461), .Z(n28463) );
  XNOR U8075 ( .A(n28464), .B(n27984), .Z(n27986) );
  XNOR U8076 ( .A(n27987), .B(n27501), .Z(n27503) );
  XNOR U8077 ( .A(n27504), .B(n27012), .Z(n27014) );
  XNOR U8078 ( .A(n27015), .B(n26515), .Z(n26517) );
  XNOR U8079 ( .A(n26518), .B(n26014), .Z(n26016) );
  XNOR U8080 ( .A(n26017), .B(n25506), .Z(n25508) );
  XNOR U8081 ( .A(n25509), .B(n24992), .Z(n24994) );
  XNOR U8082 ( .A(n23947), .B(n23413), .Z(n23415) );
  XNOR U8083 ( .A(n24467), .B(n23939), .Z(n23941) );
  XNOR U8084 ( .A(n22843), .B(n22296), .Z(n22298) );
  XNOR U8085 ( .A(n21685), .B(n21127), .Z(n21129) );
  XNOR U8086 ( .A(n23396), .B(n22855), .Z(n22857) );
  XNOR U8087 ( .A(n21735), .B(n21177), .Z(n21179) );
  XNOR U8088 ( .A(n22803), .B(n22256), .Z(n22258) );
  XNOR U8089 ( .A(n22249), .B(n21697), .Z(n21699) );
  XNOR U8090 ( .A(n20553), .B(n19983), .Z(n19985) );
  XNOR U8091 ( .A(n19976), .B(n19400), .Z(n19402) );
  XNOR U8092 ( .A(n21670), .B(n21112), .Z(n21114) );
  XNOR U8093 ( .A(n23376), .B(n22835), .Z(n22837) );
  XNOR U8094 ( .A(n21715), .B(n21157), .Z(n21159) );
  XNOR U8095 ( .A(n22873), .B(n22326), .Z(n22328) );
  XNOR U8096 ( .A(n33325), .B(n32911), .Z(n32913) );
  XNOR U8097 ( .A(n23942), .B(n23408), .Z(n23410) );
  XNOR U8098 ( .A(n22299), .B(n21747), .Z(n21749) );
  XOR U8099 ( .A(n20562), .B(n21075), .Z(n20566) );
  XNOR U8100 ( .A(n20538), .B(n19968), .Z(n19970) );
  XNOR U8101 ( .A(n19961), .B(n19385), .Z(n19387) );
  XOR U8102 ( .A(n18793), .B(n19365), .Z(n18797) );
  XNOR U8103 ( .A(n22279), .B(n21727), .Z(n21729) );
  XNOR U8104 ( .A(n21720), .B(n21162), .Z(n21164) );
  XNOR U8105 ( .A(n20583), .B(n20013), .Z(n20015) );
  XNOR U8106 ( .A(n20006), .B(n19430), .Z(n19432) );
  XNOR U8107 ( .A(n21765), .B(n21207), .Z(n21209) );
  XNOR U8108 ( .A(n35670), .B(n35292), .Z(n35294) );
  XNOR U8109 ( .A(n35295), .B(n34911), .Z(n34913) );
  XNOR U8110 ( .A(n34914), .B(n34524), .Z(n34526) );
  XNOR U8111 ( .A(n34527), .B(n34131), .Z(n34133) );
  XNOR U8112 ( .A(n34134), .B(n33732), .Z(n33734) );
  XNOR U8113 ( .A(n33330), .B(n32916), .Z(n32918) );
  XNOR U8114 ( .A(n32919), .B(n32499), .Z(n32501) );
  XNOR U8115 ( .A(n32502), .B(n32076), .Z(n32078) );
  XNOR U8116 ( .A(n32079), .B(n31647), .Z(n31649) );
  XNOR U8117 ( .A(n31650), .B(n31212), .Z(n31214) );
  XNOR U8118 ( .A(n31215), .B(n30771), .Z(n30773) );
  XNOR U8119 ( .A(n30774), .B(n30324), .Z(n30326) );
  XNOR U8120 ( .A(n30327), .B(n29871), .Z(n29873) );
  XNOR U8121 ( .A(n29874), .B(n29412), .Z(n29414) );
  XNOR U8122 ( .A(n29415), .B(n28947), .Z(n28949) );
  XNOR U8123 ( .A(n28950), .B(n28476), .Z(n28478) );
  XNOR U8124 ( .A(n28479), .B(n27999), .Z(n28001) );
  XNOR U8125 ( .A(n28002), .B(n27516), .Z(n27518) );
  XNOR U8126 ( .A(n27519), .B(n27027), .Z(n27029) );
  XNOR U8127 ( .A(n27030), .B(n26530), .Z(n26532) );
  XNOR U8128 ( .A(n26533), .B(n26029), .Z(n26031) );
  XNOR U8129 ( .A(n26032), .B(n25521), .Z(n25523) );
  XNOR U8130 ( .A(n25524), .B(n25007), .Z(n25009) );
  XNOR U8131 ( .A(n25010), .B(n24484), .Z(n24486) );
  XNOR U8132 ( .A(n24487), .B(n23959), .Z(n23961) );
  XNOR U8133 ( .A(n23962), .B(n23428), .Z(n23430) );
  XNOR U8134 ( .A(n22858), .B(n22311), .Z(n22313) );
  XNOR U8135 ( .A(n21180), .B(n20615), .Z(n20617) );
  XNOR U8136 ( .A(n19986), .B(n19410), .Z(n19412) );
  XNOR U8137 ( .A(n23431), .B(n22890), .Z(n22892) );
  XNOR U8138 ( .A(n21795), .B(n21237), .Z(n21239) );
  XNOR U8139 ( .A(n21750), .B(n21192), .Z(n21194) );
  XNOR U8140 ( .A(n20036), .B(n19460), .Z(n19462) );
  XNOR U8141 ( .A(n21140), .B(n20575), .Z(n20577) );
  XNOR U8142 ( .A(n20568), .B(n19998), .Z(n20000) );
  XOR U8143 ( .A(n17497), .B(n18088), .Z(n17501) );
  XNOR U8144 ( .A(n21730), .B(n21172), .Z(n21174) );
  XNOR U8145 ( .A(n22334), .B(n21782), .Z(n21784) );
  XNOR U8146 ( .A(n21775), .B(n21217), .Z(n21219) );
  XNOR U8147 ( .A(n21210), .B(n20645), .Z(n20647) );
  XNOR U8148 ( .A(n34537), .B(n34141), .Z(n34143) );
  XNOR U8149 ( .A(n22314), .B(n21762), .Z(n21764) );
  XNOR U8150 ( .A(n20618), .B(n20048), .Z(n20050) );
  XOR U8151 ( .A(n18124), .B(n18769), .Z(n18128) );
  XOR U8152 ( .A(n18828), .B(n19358), .Z(n18832) );
  XOR U8153 ( .A(n18808), .B(n19362), .Z(n18812) );
  XNOR U8154 ( .A(n20598), .B(n20028), .Z(n20030) );
  XNOR U8155 ( .A(n20021), .B(n19445), .Z(n19447) );
  XOR U8156 ( .A(n18853), .B(n19353), .Z(n18857) );
  XNOR U8157 ( .A(n20066), .B(n19490), .Z(n19492) );
  XNOR U8158 ( .A(n36774), .B(n36414), .Z(n36416) );
  XNOR U8159 ( .A(n36417), .B(n36051), .Z(n36053) );
  XNOR U8160 ( .A(n36054), .B(n35682), .Z(n35684) );
  XNOR U8161 ( .A(n35685), .B(n35307), .Z(n35309) );
  XNOR U8162 ( .A(n35310), .B(n34926), .Z(n34928) );
  XNOR U8163 ( .A(n34542), .B(n34146), .Z(n34148) );
  XNOR U8164 ( .A(n34149), .B(n33747), .Z(n33749) );
  XNOR U8165 ( .A(n33750), .B(n33342), .Z(n33344) );
  XNOR U8166 ( .A(n33345), .B(n32931), .Z(n32933) );
  XNOR U8167 ( .A(n32934), .B(n32514), .Z(n32516) );
  XNOR U8168 ( .A(n32517), .B(n32091), .Z(n32093) );
  XNOR U8169 ( .A(n32094), .B(n31662), .Z(n31664) );
  XNOR U8170 ( .A(n31665), .B(n31227), .Z(n31229) );
  XNOR U8171 ( .A(n31230), .B(n30786), .Z(n30788) );
  XNOR U8172 ( .A(n30789), .B(n30339), .Z(n30341) );
  XNOR U8173 ( .A(n30342), .B(n29886), .Z(n29888) );
  XNOR U8174 ( .A(n29889), .B(n29427), .Z(n29429) );
  XNOR U8175 ( .A(n29430), .B(n28962), .Z(n28964) );
  XNOR U8176 ( .A(n28965), .B(n28491), .Z(n28493) );
  XNOR U8177 ( .A(n28494), .B(n28014), .Z(n28016) );
  XNOR U8178 ( .A(n28017), .B(n27531), .Z(n27533) );
  XNOR U8179 ( .A(n27534), .B(n27042), .Z(n27044) );
  XNOR U8180 ( .A(n27045), .B(n26545), .Z(n26547) );
  XNOR U8181 ( .A(n26548), .B(n26044), .Z(n26046) );
  XNOR U8182 ( .A(n26047), .B(n25536), .Z(n25538) );
  XNOR U8183 ( .A(n25539), .B(n25022), .Z(n25024) );
  XNOR U8184 ( .A(n25025), .B(n24499), .Z(n24501) );
  XNOR U8185 ( .A(n24502), .B(n23974), .Z(n23976) );
  XNOR U8186 ( .A(n23977), .B(n23443), .Z(n23445) );
  XNOR U8187 ( .A(n23446), .B(n22905), .Z(n22907) );
  XNOR U8188 ( .A(n22364), .B(n21812), .Z(n21814) );
  XNOR U8189 ( .A(n21805), .B(n21247), .Z(n21249) );
  XNOR U8190 ( .A(n21240), .B(n20675), .Z(n20677) );
  XNOR U8191 ( .A(n21195), .B(n20630), .Z(n20632) );
  XNOR U8192 ( .A(n19463), .B(n18881), .Z(n18883) );
  XNOR U8193 ( .A(n22344), .B(n21792), .Z(n21794) );
  XNOR U8194 ( .A(n21785), .B(n21227), .Z(n21229) );
  XNOR U8195 ( .A(n20096), .B(n19520), .Z(n19522) );
  XNOR U8196 ( .A(n20051), .B(n19475), .Z(n19477) );
  XNOR U8197 ( .A(n19423), .B(n18841), .Z(n18843) );
  XOR U8198 ( .A(n17512), .B(n18085), .Z(n17516) );
  XOR U8199 ( .A(n16290), .B(n16887), .Z(n16294) );
  XNOR U8200 ( .A(n20653), .B(n20083), .Z(n20085) );
  XNOR U8201 ( .A(n20076), .B(n19500), .Z(n19502) );
  XNOR U8202 ( .A(n19493), .B(n18911), .Z(n18913) );
  XNOR U8203 ( .A(n35695), .B(n35317), .Z(n35319) );
  XNOR U8204 ( .A(n21815), .B(n21257), .Z(n21259) );
  XNOR U8205 ( .A(n20633), .B(n20063), .Z(n20065) );
  XOR U8206 ( .A(n18139), .B(n18763), .Z(n18143) );
  XOR U8207 ( .A(n16929), .B(n17484), .Z(n16933) );
  XOR U8208 ( .A(n15049), .B(n15664), .Z(n15053) );
  XOR U8209 ( .A(n18868), .B(n19350), .Z(n18872) );
  XOR U8210 ( .A(n17562), .B(n18075), .Z(n17566) );
  XNOR U8211 ( .A(n20126), .B(n19550), .Z(n19552) );
  XNOR U8212 ( .A(n37824), .B(n37482), .Z(n37484) );
  XNOR U8213 ( .A(n37485), .B(n37137), .Z(n37139) );
  XNOR U8214 ( .A(n37140), .B(n36786), .Z(n36788) );
  XNOR U8215 ( .A(n36789), .B(n36429), .Z(n36431) );
  XNOR U8216 ( .A(n36432), .B(n36066), .Z(n36068) );
  XNOR U8217 ( .A(n35700), .B(n35322), .Z(n35324) );
  XNOR U8218 ( .A(n35325), .B(n34941), .Z(n34943) );
  XNOR U8219 ( .A(n34944), .B(n34554), .Z(n34556) );
  XNOR U8220 ( .A(n34557), .B(n34161), .Z(n34163) );
  XNOR U8221 ( .A(n34164), .B(n33762), .Z(n33764) );
  XNOR U8222 ( .A(n33765), .B(n33357), .Z(n33359) );
  XNOR U8223 ( .A(n33360), .B(n32946), .Z(n32948) );
  XNOR U8224 ( .A(n32949), .B(n32529), .Z(n32531) );
  XNOR U8225 ( .A(n32532), .B(n32106), .Z(n32108) );
  XNOR U8226 ( .A(n32109), .B(n31677), .Z(n31679) );
  XNOR U8227 ( .A(n31680), .B(n31242), .Z(n31244) );
  XNOR U8228 ( .A(n31245), .B(n30801), .Z(n30803) );
  XNOR U8229 ( .A(n30804), .B(n30354), .Z(n30356) );
  XNOR U8230 ( .A(n30357), .B(n29901), .Z(n29903) );
  XNOR U8231 ( .A(n29904), .B(n29442), .Z(n29444) );
  XNOR U8232 ( .A(n29445), .B(n28977), .Z(n28979) );
  XNOR U8233 ( .A(n28980), .B(n28506), .Z(n28508) );
  XNOR U8234 ( .A(n28509), .B(n28029), .Z(n28031) );
  XNOR U8235 ( .A(n28032), .B(n27546), .Z(n27548) );
  XNOR U8236 ( .A(n27549), .B(n27057), .Z(n27059) );
  XNOR U8237 ( .A(n27060), .B(n26560), .Z(n26562) );
  XNOR U8238 ( .A(n26563), .B(n26059), .Z(n26061) );
  XNOR U8239 ( .A(n26062), .B(n25551), .Z(n25553) );
  XNOR U8240 ( .A(n25554), .B(n25037), .Z(n25039) );
  XNOR U8241 ( .A(n25040), .B(n24514), .Z(n24516) );
  XNOR U8242 ( .A(n24517), .B(n23989), .Z(n23991) );
  XNOR U8243 ( .A(n23992), .B(n23458), .Z(n23460) );
  XNOR U8244 ( .A(n23461), .B(n22920), .Z(n22922) );
  XNOR U8245 ( .A(n22923), .B(n22376), .Z(n22378) );
  XNOR U8246 ( .A(n22379), .B(n21827), .Z(n21829) );
  XNOR U8247 ( .A(n21830), .B(n21272), .Z(n21274) );
  XNOR U8248 ( .A(n20683), .B(n20113), .Z(n20115) );
  XNOR U8249 ( .A(n20106), .B(n19530), .Z(n19532) );
  XNOR U8250 ( .A(n19523), .B(n18941), .Z(n18943) );
  XNOR U8251 ( .A(n19478), .B(n18896), .Z(n18898) );
  XOR U8252 ( .A(n18189), .B(n18743), .Z(n18193) );
  XOR U8253 ( .A(n15700), .B(n16273), .Z(n15704) );
  XOR U8254 ( .A(n16345), .B(n16876), .Z(n16349) );
  XNOR U8255 ( .A(n20663), .B(n20093), .Z(n20095) );
  XOR U8256 ( .A(n16305), .B(n16884), .Z(n16309) );
  XOR U8257 ( .A(n18923), .B(n19339), .Z(n18927) );
  XOR U8258 ( .A(n17617), .B(n18064), .Z(n17621) );
  XNOR U8259 ( .A(n20713), .B(n20143), .Z(n20145) );
  XNOR U8260 ( .A(n20136), .B(n19560), .Z(n19562) );
  XNOR U8261 ( .A(n19553), .B(n18971), .Z(n18973) );
  XNOR U8262 ( .A(n36799), .B(n36439), .Z(n36441) );
  XNOR U8263 ( .A(n20693), .B(n20123), .Z(n20125) );
  XOR U8264 ( .A(n16944), .B(n17481), .Z(n16948) );
  XOR U8265 ( .A(n15064), .B(n15661), .Z(n15068) );
  XOR U8266 ( .A(n13794), .B(n14415), .Z(n13798) );
  XOR U8267 ( .A(n17577), .B(n18072), .Z(n17581) );
  XNOR U8268 ( .A(n38820), .B(n38496), .Z(n38498) );
  XNOR U8269 ( .A(n38499), .B(n38169), .Z(n38171) );
  XNOR U8270 ( .A(n38172), .B(n37836), .Z(n37838) );
  XNOR U8271 ( .A(n37839), .B(n37497), .Z(n37499) );
  XNOR U8272 ( .A(n37500), .B(n37152), .Z(n37154) );
  XNOR U8273 ( .A(n36804), .B(n36444), .Z(n36446) );
  XNOR U8274 ( .A(n36447), .B(n36081), .Z(n36083) );
  XNOR U8275 ( .A(n36084), .B(n35712), .Z(n35714) );
  XNOR U8276 ( .A(n35715), .B(n35337), .Z(n35339) );
  XNOR U8277 ( .A(n35340), .B(n34956), .Z(n34958) );
  XNOR U8278 ( .A(n34959), .B(n34569), .Z(n34571) );
  XNOR U8279 ( .A(n34572), .B(n34176), .Z(n34178) );
  XNOR U8280 ( .A(n34179), .B(n33777), .Z(n33779) );
  XNOR U8281 ( .A(n33780), .B(n33372), .Z(n33374) );
  XNOR U8282 ( .A(n33375), .B(n32961), .Z(n32963) );
  XNOR U8283 ( .A(n32964), .B(n32544), .Z(n32546) );
  XNOR U8284 ( .A(n32547), .B(n32121), .Z(n32123) );
  XNOR U8285 ( .A(n32124), .B(n31692), .Z(n31694) );
  XNOR U8286 ( .A(n31695), .B(n31257), .Z(n31259) );
  XNOR U8287 ( .A(n31260), .B(n30816), .Z(n30818) );
  XNOR U8288 ( .A(n30819), .B(n30369), .Z(n30371) );
  XNOR U8289 ( .A(n30372), .B(n29916), .Z(n29918) );
  XNOR U8290 ( .A(n29919), .B(n29457), .Z(n29459) );
  XNOR U8291 ( .A(n29460), .B(n28992), .Z(n28994) );
  XNOR U8292 ( .A(n28995), .B(n28521), .Z(n28523) );
  XNOR U8293 ( .A(n28524), .B(n28044), .Z(n28046) );
  XNOR U8294 ( .A(n28047), .B(n27561), .Z(n27563) );
  XNOR U8295 ( .A(n27564), .B(n27072), .Z(n27074) );
  XNOR U8296 ( .A(n27075), .B(n26575), .Z(n26577) );
  XNOR U8297 ( .A(n26578), .B(n26074), .Z(n26076) );
  XNOR U8298 ( .A(n26077), .B(n25566), .Z(n25568) );
  XNOR U8299 ( .A(n25569), .B(n25052), .Z(n25054) );
  XNOR U8300 ( .A(n25055), .B(n24529), .Z(n24531) );
  XNOR U8301 ( .A(n24532), .B(n24004), .Z(n24006) );
  XNOR U8302 ( .A(n24007), .B(n23473), .Z(n23475) );
  XNOR U8303 ( .A(n23476), .B(n22935), .Z(n22937) );
  XNOR U8304 ( .A(n22938), .B(n22391), .Z(n22393) );
  XNOR U8305 ( .A(n22394), .B(n21842), .Z(n21844) );
  XNOR U8306 ( .A(n21845), .B(n21287), .Z(n21289) );
  XNOR U8307 ( .A(n20728), .B(n20158), .Z(n20160) );
  XNOR U8308 ( .A(n20161), .B(n19585), .Z(n19587) );
  XOR U8309 ( .A(n18953), .B(n19333), .Z(n18957) );
  XOR U8310 ( .A(n17647), .B(n18058), .Z(n17651) );
  XOR U8311 ( .A(n18204), .B(n18737), .Z(n18208) );
  XOR U8312 ( .A(n16994), .B(n17471), .Z(n16998) );
  XOR U8313 ( .A(n15760), .B(n16261), .Z(n15764) );
  XOR U8314 ( .A(n15715), .B(n16270), .Z(n15719) );
  XOR U8315 ( .A(n14457), .B(n15036), .Z(n14461) );
  XOR U8316 ( .A(n12505), .B(n13144), .Z(n12509) );
  XOR U8317 ( .A(n16360), .B(n16873), .Z(n16364) );
  XOR U8318 ( .A(n15114), .B(n15651), .Z(n15118) );
  XNOR U8319 ( .A(n20723), .B(n20153), .Z(n20155) );
  XOR U8320 ( .A(n19003), .B(n19323), .Z(n19007) );
  XOR U8321 ( .A(n13180), .B(n13777), .Z(n13184) );
  XOR U8322 ( .A(n13849), .B(n14404), .Z(n13853) );
  XOR U8323 ( .A(n18234), .B(n18725), .Z(n18238) );
  XOR U8324 ( .A(n17024), .B(n17465), .Z(n17028) );
  XOR U8325 ( .A(n15790), .B(n16255), .Z(n15794) );
  XOR U8326 ( .A(n18983), .B(n19327), .Z(n18987) );
  XOR U8327 ( .A(n17677), .B(n18052), .Z(n17681) );
  XNOR U8328 ( .A(n37849), .B(n37507), .Z(n37509) );
  XOR U8329 ( .A(n13809), .B(n14412), .Z(n13813) );
  XNOR U8330 ( .A(n39762), .B(n39456), .Z(n39458) );
  XNOR U8331 ( .A(n39459), .B(n39147), .Z(n39149) );
  XNOR U8332 ( .A(n39150), .B(n38832), .Z(n38834) );
  XNOR U8333 ( .A(n38835), .B(n38511), .Z(n38513) );
  XNOR U8334 ( .A(n38514), .B(n38184), .Z(n38186) );
  XNOR U8335 ( .A(n37854), .B(n37512), .Z(n37514) );
  XNOR U8336 ( .A(n37515), .B(n37167), .Z(n37169) );
  XNOR U8337 ( .A(n37170), .B(n36816), .Z(n36818) );
  XNOR U8338 ( .A(n36819), .B(n36459), .Z(n36461) );
  XNOR U8339 ( .A(n36462), .B(n36096), .Z(n36098) );
  XNOR U8340 ( .A(n36099), .B(n35727), .Z(n35729) );
  XNOR U8341 ( .A(n35730), .B(n35352), .Z(n35354) );
  XNOR U8342 ( .A(n35355), .B(n34971), .Z(n34973) );
  XNOR U8343 ( .A(n34974), .B(n34584), .Z(n34586) );
  XNOR U8344 ( .A(n34587), .B(n34191), .Z(n34193) );
  XNOR U8345 ( .A(n34194), .B(n33792), .Z(n33794) );
  XNOR U8346 ( .A(n33795), .B(n33387), .Z(n33389) );
  XNOR U8347 ( .A(n33390), .B(n32976), .Z(n32978) );
  XNOR U8348 ( .A(n32979), .B(n32559), .Z(n32561) );
  XNOR U8349 ( .A(n32562), .B(n32136), .Z(n32138) );
  XNOR U8350 ( .A(n32139), .B(n31707), .Z(n31709) );
  XNOR U8351 ( .A(n31710), .B(n31272), .Z(n31274) );
  XNOR U8352 ( .A(n31275), .B(n30831), .Z(n30833) );
  XNOR U8353 ( .A(n30834), .B(n30384), .Z(n30386) );
  XNOR U8354 ( .A(n30387), .B(n29931), .Z(n29933) );
  XNOR U8355 ( .A(n29934), .B(n29472), .Z(n29474) );
  XNOR U8356 ( .A(n29475), .B(n29007), .Z(n29009) );
  XNOR U8357 ( .A(n29010), .B(n28536), .Z(n28538) );
  XNOR U8358 ( .A(n28539), .B(n28059), .Z(n28061) );
  XNOR U8359 ( .A(n28062), .B(n27576), .Z(n27578) );
  XNOR U8360 ( .A(n27579), .B(n27087), .Z(n27089) );
  XNOR U8361 ( .A(n27090), .B(n26590), .Z(n26592) );
  XNOR U8362 ( .A(n26593), .B(n26089), .Z(n26091) );
  XNOR U8363 ( .A(n26092), .B(n25581), .Z(n25583) );
  XNOR U8364 ( .A(n25584), .B(n25067), .Z(n25069) );
  XNOR U8365 ( .A(n25070), .B(n24544), .Z(n24546) );
  XNOR U8366 ( .A(n24547), .B(n24019), .Z(n24021) );
  XNOR U8367 ( .A(n24022), .B(n23488), .Z(n23490) );
  XNOR U8368 ( .A(n23491), .B(n22950), .Z(n22952) );
  XNOR U8369 ( .A(n22953), .B(n22406), .Z(n22408) );
  XNOR U8370 ( .A(n22409), .B(n21857), .Z(n21859) );
  XNOR U8371 ( .A(n21860), .B(n21302), .Z(n21304) );
  XNOR U8372 ( .A(n21305), .B(n20740), .Z(n20742) );
  XNOR U8373 ( .A(n20743), .B(n20173), .Z(n20175) );
  XNOR U8374 ( .A(n19598), .B(n19016), .Z(n19018) );
  XOR U8375 ( .A(n17707), .B(n18046), .Z(n17711) );
  XOR U8376 ( .A(n18264), .B(n18713), .Z(n18268) );
  XOR U8377 ( .A(n17054), .B(n17459), .Z(n17058) );
  XOR U8378 ( .A(n15820), .B(n16249), .Z(n15824) );
  XOR U8379 ( .A(n16395), .B(n16866), .Z(n16399) );
  XOR U8380 ( .A(n15149), .B(n15644), .Z(n15153) );
  XOR U8381 ( .A(n13879), .B(n14398), .Z(n13883) );
  XOR U8382 ( .A(n14472), .B(n15033), .Z(n14476) );
  XOR U8383 ( .A(n12520), .B(n13141), .Z(n12524) );
  XOR U8384 ( .A(n11200), .B(n11845), .Z(n11204) );
  XOR U8385 ( .A(n15129), .B(n15648), .Z(n15133) );
  XOR U8386 ( .A(n13195), .B(n13774), .Z(n13199) );
  XOR U8387 ( .A(n11887), .B(n12492), .Z(n11891) );
  XOR U8388 ( .A(n9863), .B(n10526), .Z(n9867) );
  XOR U8389 ( .A(n13864), .B(n14401), .Z(n13868) );
  XOR U8390 ( .A(n12570), .B(n13131), .Z(n12574) );
  XOR U8391 ( .A(n16425), .B(n16860), .Z(n16429) );
  XOR U8392 ( .A(n15179), .B(n15638), .Z(n15183) );
  XOR U8393 ( .A(n13909), .B(n14392), .Z(n13913) );
  XOR U8394 ( .A(n18294), .B(n18701), .Z(n18298) );
  XOR U8395 ( .A(n17084), .B(n17453), .Z(n17088) );
  XOR U8396 ( .A(n15850), .B(n16243), .Z(n15854) );
  XOR U8397 ( .A(n17737), .B(n18040), .Z(n17741) );
  XNOR U8398 ( .A(n38845), .B(n38521), .Z(n38523) );
  XOR U8399 ( .A(n10562), .B(n11183), .Z(n10566) );
  XNOR U8400 ( .A(n40650), .B(n40362), .Z(n40364) );
  XNOR U8401 ( .A(n40365), .B(n40071), .Z(n40073) );
  XNOR U8402 ( .A(n40074), .B(n39774), .Z(n39776) );
  XNOR U8403 ( .A(n39777), .B(n39471), .Z(n39473) );
  XNOR U8404 ( .A(n39474), .B(n39162), .Z(n39164) );
  XNOR U8405 ( .A(n38850), .B(n38526), .Z(n38528) );
  XNOR U8406 ( .A(n38529), .B(n38199), .Z(n38201) );
  XNOR U8407 ( .A(n38202), .B(n37866), .Z(n37868) );
  XNOR U8408 ( .A(n37869), .B(n37527), .Z(n37529) );
  XNOR U8409 ( .A(n37530), .B(n37182), .Z(n37184) );
  XNOR U8410 ( .A(n37185), .B(n36831), .Z(n36833) );
  XNOR U8411 ( .A(n36834), .B(n36474), .Z(n36476) );
  XNOR U8412 ( .A(n36477), .B(n36111), .Z(n36113) );
  XNOR U8413 ( .A(n36114), .B(n35742), .Z(n35744) );
  XNOR U8414 ( .A(n35745), .B(n35367), .Z(n35369) );
  XNOR U8415 ( .A(n35370), .B(n34986), .Z(n34988) );
  XNOR U8416 ( .A(n34989), .B(n34599), .Z(n34601) );
  XNOR U8417 ( .A(n34602), .B(n34206), .Z(n34208) );
  XNOR U8418 ( .A(n34209), .B(n33807), .Z(n33809) );
  XNOR U8419 ( .A(n33810), .B(n33402), .Z(n33404) );
  XNOR U8420 ( .A(n33405), .B(n32991), .Z(n32993) );
  XNOR U8421 ( .A(n32994), .B(n32574), .Z(n32576) );
  XNOR U8422 ( .A(n32577), .B(n32151), .Z(n32153) );
  XNOR U8423 ( .A(n32154), .B(n31722), .Z(n31724) );
  XNOR U8424 ( .A(n31725), .B(n31287), .Z(n31289) );
  XNOR U8425 ( .A(n31290), .B(n30846), .Z(n30848) );
  XNOR U8426 ( .A(n30849), .B(n30399), .Z(n30401) );
  XNOR U8427 ( .A(n30402), .B(n29946), .Z(n29948) );
  XNOR U8428 ( .A(n29949), .B(n29487), .Z(n29489) );
  XNOR U8429 ( .A(n29490), .B(n29022), .Z(n29024) );
  XNOR U8430 ( .A(n29025), .B(n28551), .Z(n28553) );
  XNOR U8431 ( .A(n28554), .B(n28074), .Z(n28076) );
  XNOR U8432 ( .A(n28077), .B(n27591), .Z(n27593) );
  XNOR U8433 ( .A(n27594), .B(n27102), .Z(n27104) );
  XNOR U8434 ( .A(n27105), .B(n26605), .Z(n26607) );
  XNOR U8435 ( .A(n26608), .B(n26104), .Z(n26106) );
  XNOR U8436 ( .A(n26107), .B(n25596), .Z(n25598) );
  XNOR U8437 ( .A(n25599), .B(n25082), .Z(n25084) );
  XNOR U8438 ( .A(n25085), .B(n24559), .Z(n24561) );
  XNOR U8439 ( .A(n24562), .B(n24034), .Z(n24036) );
  XNOR U8440 ( .A(n24037), .B(n23503), .Z(n23505) );
  XNOR U8441 ( .A(n23506), .B(n22965), .Z(n22967) );
  XNOR U8442 ( .A(n22968), .B(n22421), .Z(n22423) );
  XNOR U8443 ( .A(n22424), .B(n21872), .Z(n21874) );
  XNOR U8444 ( .A(n21875), .B(n21317), .Z(n21319) );
  XNOR U8445 ( .A(n21320), .B(n20755), .Z(n20757) );
  XNOR U8446 ( .A(n20758), .B(n20188), .Z(n20190) );
  XNOR U8447 ( .A(n20191), .B(n19615), .Z(n19617) );
  XNOR U8448 ( .A(n19618), .B(n19036), .Z(n19038) );
  XOR U8449 ( .A(n18324), .B(n18689), .Z(n18328) );
  XOR U8450 ( .A(n17114), .B(n17447), .Z(n17118) );
  XOR U8451 ( .A(n15880), .B(n16237), .Z(n15884) );
  XOR U8452 ( .A(n16455), .B(n16854), .Z(n16459) );
  XOR U8453 ( .A(n15209), .B(n15632), .Z(n15213) );
  XOR U8454 ( .A(n13939), .B(n14386), .Z(n13943) );
  XOR U8455 ( .A(n14532), .B(n15021), .Z(n14536) );
  XOR U8456 ( .A(n13250), .B(n13763), .Z(n13254) );
  XOR U8457 ( .A(n11942), .B(n12481), .Z(n11946) );
  XOR U8458 ( .A(n11215), .B(n11842), .Z(n11219) );
  XOR U8459 ( .A(n11902), .B(n12489), .Z(n11906) );
  XOR U8460 ( .A(n9878), .B(n10523), .Z(n9882) );
  XOR U8461 ( .A(n8512), .B(n9181), .Z(n8516) );
  XOR U8462 ( .A(n12585), .B(n13128), .Z(n12589) );
  XOR U8463 ( .A(n11265), .B(n11832), .Z(n11269) );
  XOR U8464 ( .A(n14562), .B(n15015), .Z(n14566) );
  XOR U8465 ( .A(n13280), .B(n13757), .Z(n13284) );
  XOR U8466 ( .A(n11972), .B(n12475), .Z(n11976) );
  XOR U8467 ( .A(n16485), .B(n16848), .Z(n16489) );
  XOR U8468 ( .A(n15239), .B(n15626), .Z(n15243) );
  XOR U8469 ( .A(n13969), .B(n14380), .Z(n13973) );
  XOR U8470 ( .A(n17144), .B(n17441), .Z(n17148) );
  XOR U8471 ( .A(n15910), .B(n16231), .Z(n15914) );
  XNOR U8472 ( .A(n39787), .B(n39481), .Z(n39483) );
  XOR U8473 ( .A(n10577), .B(n11180), .Z(n10581) );
  XOR U8474 ( .A(n9223), .B(n9850), .Z(n9227) );
  XOR U8475 ( .A(n7127), .B(n7814), .Z(n7131) );
  XOR U8476 ( .A(n9928), .B(n10513), .Z(n9932) );
  XNOR U8477 ( .A(n41484), .B(n41214), .Z(n41216) );
  XNOR U8478 ( .A(n41217), .B(n40941), .Z(n40943) );
  XNOR U8479 ( .A(n40944), .B(n40662), .Z(n40664) );
  XNOR U8480 ( .A(n40665), .B(n40377), .Z(n40379) );
  XNOR U8481 ( .A(n40380), .B(n40086), .Z(n40088) );
  XNOR U8482 ( .A(n39792), .B(n39486), .Z(n39488) );
  XNOR U8483 ( .A(n39489), .B(n39177), .Z(n39179) );
  XNOR U8484 ( .A(n39180), .B(n38862), .Z(n38864) );
  XNOR U8485 ( .A(n38865), .B(n38541), .Z(n38543) );
  XNOR U8486 ( .A(n38544), .B(n38214), .Z(n38216) );
  XNOR U8487 ( .A(n38217), .B(n37881), .Z(n37883) );
  XNOR U8488 ( .A(n37884), .B(n37542), .Z(n37544) );
  XNOR U8489 ( .A(n37545), .B(n37197), .Z(n37199) );
  XNOR U8490 ( .A(n37200), .B(n36846), .Z(n36848) );
  XNOR U8491 ( .A(n36849), .B(n36489), .Z(n36491) );
  XNOR U8492 ( .A(n36492), .B(n36126), .Z(n36128) );
  XNOR U8493 ( .A(n36129), .B(n35757), .Z(n35759) );
  XNOR U8494 ( .A(n35760), .B(n35382), .Z(n35384) );
  XNOR U8495 ( .A(n35385), .B(n35001), .Z(n35003) );
  XNOR U8496 ( .A(n35004), .B(n34614), .Z(n34616) );
  XNOR U8497 ( .A(n34617), .B(n34221), .Z(n34223) );
  XNOR U8498 ( .A(n34224), .B(n33822), .Z(n33824) );
  XNOR U8499 ( .A(n33825), .B(n33417), .Z(n33419) );
  XNOR U8500 ( .A(n33420), .B(n33006), .Z(n33008) );
  XNOR U8501 ( .A(n33009), .B(n32589), .Z(n32591) );
  XNOR U8502 ( .A(n32592), .B(n32166), .Z(n32168) );
  XNOR U8503 ( .A(n32169), .B(n31737), .Z(n31739) );
  XNOR U8504 ( .A(n31740), .B(n31302), .Z(n31304) );
  XNOR U8505 ( .A(n31305), .B(n30861), .Z(n30863) );
  XNOR U8506 ( .A(n30864), .B(n30414), .Z(n30416) );
  XNOR U8507 ( .A(n30417), .B(n29961), .Z(n29963) );
  XNOR U8508 ( .A(n29964), .B(n29502), .Z(n29504) );
  XNOR U8509 ( .A(n29505), .B(n29037), .Z(n29039) );
  XNOR U8510 ( .A(n29040), .B(n28566), .Z(n28568) );
  XNOR U8511 ( .A(n28569), .B(n28089), .Z(n28091) );
  XNOR U8512 ( .A(n28092), .B(n27606), .Z(n27608) );
  XNOR U8513 ( .A(n27609), .B(n27117), .Z(n27119) );
  XNOR U8514 ( .A(n27120), .B(n26620), .Z(n26622) );
  XNOR U8515 ( .A(n26623), .B(n26119), .Z(n26121) );
  XNOR U8516 ( .A(n26122), .B(n25611), .Z(n25613) );
  XNOR U8517 ( .A(n25614), .B(n25097), .Z(n25099) );
  XNOR U8518 ( .A(n25100), .B(n24574), .Z(n24576) );
  XNOR U8519 ( .A(n24577), .B(n24049), .Z(n24051) );
  XNOR U8520 ( .A(n24052), .B(n23518), .Z(n23520) );
  XNOR U8521 ( .A(n23521), .B(n22980), .Z(n22982) );
  XNOR U8522 ( .A(n22983), .B(n22436), .Z(n22438) );
  XNOR U8523 ( .A(n22439), .B(n21887), .Z(n21889) );
  XNOR U8524 ( .A(n21890), .B(n21332), .Z(n21334) );
  XNOR U8525 ( .A(n21335), .B(n20770), .Z(n20772) );
  XNOR U8526 ( .A(n20773), .B(n20203), .Z(n20205) );
  XNOR U8527 ( .A(n20206), .B(n19630), .Z(n19632) );
  XNOR U8528 ( .A(n19633), .B(n19051), .Z(n19053) );
  XOR U8529 ( .A(n18359), .B(n18675), .Z(n18363) );
  XOR U8530 ( .A(n17169), .B(n17436), .Z(n17173) );
  XOR U8531 ( .A(n15940), .B(n16225), .Z(n15944) );
  XOR U8532 ( .A(n16515), .B(n16842), .Z(n16519) );
  XOR U8533 ( .A(n15269), .B(n15620), .Z(n15273) );
  XOR U8534 ( .A(n13999), .B(n14374), .Z(n14003) );
  XOR U8535 ( .A(n14592), .B(n15009), .Z(n14596) );
  XOR U8536 ( .A(n13310), .B(n13751), .Z(n13314) );
  XOR U8537 ( .A(n12002), .B(n12469), .Z(n12006) );
  XOR U8538 ( .A(n12615), .B(n13122), .Z(n12619) );
  XOR U8539 ( .A(n11295), .B(n11826), .Z(n11299) );
  XOR U8540 ( .A(n9953), .B(n10508), .Z(n9957) );
  XOR U8541 ( .A(n7850), .B(n8495), .Z(n7854) );
  XOR U8542 ( .A(n8527), .B(n9178), .Z(n8531) );
  XOR U8543 ( .A(n10612), .B(n11173), .Z(n10616) );
  XOR U8544 ( .A(n7880), .B(n8489), .Z(n7884) );
  XOR U8545 ( .A(n12645), .B(n13116), .Z(n12649) );
  XOR U8546 ( .A(n11325), .B(n11820), .Z(n11329) );
  XOR U8547 ( .A(n9983), .B(n10502), .Z(n9987) );
  XOR U8548 ( .A(n14622), .B(n15003), .Z(n14626) );
  XOR U8549 ( .A(n13340), .B(n13745), .Z(n13344) );
  XOR U8550 ( .A(n12032), .B(n12463), .Z(n12036) );
  XOR U8551 ( .A(n16545), .B(n16836), .Z(n16549) );
  XOR U8552 ( .A(n15299), .B(n15614), .Z(n15303) );
  XOR U8553 ( .A(n14029), .B(n14368), .Z(n14033) );
  XNOR U8554 ( .A(n40675), .B(n40387), .Z(n40389) );
  XOR U8555 ( .A(n9238), .B(n9847), .Z(n9242) );
  XOR U8556 ( .A(n7142), .B(n7811), .Z(n7146) );
  XOR U8557 ( .A(n5728), .B(n6421), .Z(n5732) );
  XOR U8558 ( .A(n9263), .B(n9842), .Z(n9267) );
  XNOR U8559 ( .A(n42264), .B(n42012), .Z(n42014) );
  XNOR U8560 ( .A(n42015), .B(n41757), .Z(n41759) );
  XNOR U8561 ( .A(n41760), .B(n41496), .Z(n41498) );
  XNOR U8562 ( .A(n41499), .B(n41229), .Z(n41231) );
  XNOR U8563 ( .A(n41232), .B(n40956), .Z(n40958) );
  XNOR U8564 ( .A(n40680), .B(n40392), .Z(n40394) );
  XNOR U8565 ( .A(n40395), .B(n40101), .Z(n40103) );
  XNOR U8566 ( .A(n40104), .B(n39804), .Z(n39806) );
  XNOR U8567 ( .A(n39807), .B(n39501), .Z(n39503) );
  XNOR U8568 ( .A(n39504), .B(n39192), .Z(n39194) );
  XNOR U8569 ( .A(n39195), .B(n38877), .Z(n38879) );
  XNOR U8570 ( .A(n38880), .B(n38556), .Z(n38558) );
  XNOR U8571 ( .A(n38559), .B(n38229), .Z(n38231) );
  XNOR U8572 ( .A(n38232), .B(n37896), .Z(n37898) );
  XNOR U8573 ( .A(n37899), .B(n37557), .Z(n37559) );
  XNOR U8574 ( .A(n37560), .B(n37212), .Z(n37214) );
  XNOR U8575 ( .A(n37215), .B(n36861), .Z(n36863) );
  XNOR U8576 ( .A(n36864), .B(n36504), .Z(n36506) );
  XNOR U8577 ( .A(n36507), .B(n36141), .Z(n36143) );
  XNOR U8578 ( .A(n36144), .B(n35772), .Z(n35774) );
  XNOR U8579 ( .A(n35775), .B(n35397), .Z(n35399) );
  XNOR U8580 ( .A(n35400), .B(n35016), .Z(n35018) );
  XNOR U8581 ( .A(n35019), .B(n34629), .Z(n34631) );
  XNOR U8582 ( .A(n34632), .B(n34236), .Z(n34238) );
  XNOR U8583 ( .A(n34239), .B(n33837), .Z(n33839) );
  XNOR U8584 ( .A(n33840), .B(n33432), .Z(n33434) );
  XNOR U8585 ( .A(n33435), .B(n33021), .Z(n33023) );
  XNOR U8586 ( .A(n33024), .B(n32604), .Z(n32606) );
  XNOR U8587 ( .A(n32607), .B(n32181), .Z(n32183) );
  XNOR U8588 ( .A(n32184), .B(n31752), .Z(n31754) );
  XNOR U8589 ( .A(n31755), .B(n31317), .Z(n31319) );
  XNOR U8590 ( .A(n31320), .B(n30876), .Z(n30878) );
  XNOR U8591 ( .A(n30879), .B(n30429), .Z(n30431) );
  XNOR U8592 ( .A(n30432), .B(n29976), .Z(n29978) );
  XNOR U8593 ( .A(n29979), .B(n29517), .Z(n29519) );
  XNOR U8594 ( .A(n29520), .B(n29052), .Z(n29054) );
  XNOR U8595 ( .A(n29055), .B(n28581), .Z(n28583) );
  XNOR U8596 ( .A(n28584), .B(n28104), .Z(n28106) );
  XNOR U8597 ( .A(n28107), .B(n27621), .Z(n27623) );
  XNOR U8598 ( .A(n27624), .B(n27132), .Z(n27134) );
  XNOR U8599 ( .A(n27135), .B(n26635), .Z(n26637) );
  XNOR U8600 ( .A(n26638), .B(n26134), .Z(n26136) );
  XNOR U8601 ( .A(n26137), .B(n25626), .Z(n25628) );
  XNOR U8602 ( .A(n25629), .B(n25112), .Z(n25114) );
  XNOR U8603 ( .A(n25115), .B(n24589), .Z(n24591) );
  XNOR U8604 ( .A(n24592), .B(n24064), .Z(n24066) );
  XNOR U8605 ( .A(n24067), .B(n23533), .Z(n23535) );
  XNOR U8606 ( .A(n23536), .B(n22995), .Z(n22997) );
  XNOR U8607 ( .A(n22998), .B(n22451), .Z(n22453) );
  XNOR U8608 ( .A(n22454), .B(n21902), .Z(n21904) );
  XNOR U8609 ( .A(n21905), .B(n21347), .Z(n21349) );
  XNOR U8610 ( .A(n21350), .B(n20785), .Z(n20787) );
  XNOR U8611 ( .A(n20788), .B(n20218), .Z(n20220) );
  XNOR U8612 ( .A(n20221), .B(n19645), .Z(n19647) );
  XNOR U8613 ( .A(n19648), .B(n19066), .Z(n19068) );
  XOR U8614 ( .A(n17782), .B(n18031), .Z(n17786) );
  XOR U8615 ( .A(n16575), .B(n16830), .Z(n16579) );
  XOR U8616 ( .A(n15329), .B(n15608), .Z(n15333) );
  XOR U8617 ( .A(n14059), .B(n14362), .Z(n14063) );
  XOR U8618 ( .A(n14652), .B(n14997), .Z(n14656) );
  XOR U8619 ( .A(n13370), .B(n13739), .Z(n13374) );
  XOR U8620 ( .A(n12062), .B(n12457), .Z(n12066) );
  XOR U8621 ( .A(n12675), .B(n13110), .Z(n12679) );
  XOR U8622 ( .A(n11355), .B(n11814), .Z(n11359) );
  XOR U8623 ( .A(n10013), .B(n10496), .Z(n10017) );
  XOR U8624 ( .A(n10642), .B(n11167), .Z(n10646) );
  XOR U8625 ( .A(n8602), .B(n9163), .Z(n8606) );
  XOR U8626 ( .A(n7865), .B(n8492), .Z(n7869) );
  XOR U8627 ( .A(n6463), .B(n7114), .Z(n6467) );
  XOR U8628 ( .A(n4293), .B(n5004), .Z(n4297) );
  XOR U8629 ( .A(n15354), .B(n15603), .Z(n15358) );
  XOR U8630 ( .A(n9293), .B(n9836), .Z(n9297) );
  XOR U8631 ( .A(n7197), .B(n7800), .Z(n7201) );
  XOR U8632 ( .A(n5783), .B(n6410), .Z(n5787) );
  XOR U8633 ( .A(n10672), .B(n11161), .Z(n10676) );
  XOR U8634 ( .A(n8632), .B(n9157), .Z(n8636) );
  XOR U8635 ( .A(n12705), .B(n13104), .Z(n12709) );
  XOR U8636 ( .A(n11385), .B(n11808), .Z(n11389) );
  XOR U8637 ( .A(n10043), .B(n10490), .Z(n10047) );
  XOR U8638 ( .A(n14682), .B(n14991), .Z(n14686) );
  XOR U8639 ( .A(n13400), .B(n13733), .Z(n13404) );
  XOR U8640 ( .A(n12092), .B(n12451), .Z(n12096) );
  XOR U8641 ( .A(n14089), .B(n14356), .Z(n14093) );
  XNOR U8642 ( .A(n41509), .B(n41239), .Z(n41241) );
  XOR U8643 ( .A(n5743), .B(n6418), .Z(n5747) );
  XOR U8644 ( .A(n7900), .B(n8485), .Z(n7904) );
  XOR U8645 ( .A(n9323), .B(n9830), .Z(n9327) );
  XNOR U8646 ( .A(n42990), .B(n42756), .Z(n42758) );
  XNOR U8647 ( .A(n42759), .B(n42519), .Z(n42521) );
  XNOR U8648 ( .A(n42522), .B(n42276), .Z(n42278) );
  XNOR U8649 ( .A(n42279), .B(n42027), .Z(n42029) );
  XNOR U8650 ( .A(n42030), .B(n41772), .Z(n41774) );
  XNOR U8651 ( .A(n41514), .B(n41244), .Z(n41246) );
  XNOR U8652 ( .A(n41247), .B(n40971), .Z(n40973) );
  XNOR U8653 ( .A(n40974), .B(n40692), .Z(n40694) );
  XNOR U8654 ( .A(n40695), .B(n40407), .Z(n40409) );
  XNOR U8655 ( .A(n40410), .B(n40116), .Z(n40118) );
  XNOR U8656 ( .A(n40119), .B(n39819), .Z(n39821) );
  XNOR U8657 ( .A(n39822), .B(n39516), .Z(n39518) );
  XNOR U8658 ( .A(n39519), .B(n39207), .Z(n39209) );
  XNOR U8659 ( .A(n39210), .B(n38892), .Z(n38894) );
  XNOR U8660 ( .A(n38895), .B(n38571), .Z(n38573) );
  XNOR U8661 ( .A(n38574), .B(n38244), .Z(n38246) );
  XNOR U8662 ( .A(n38247), .B(n37911), .Z(n37913) );
  XNOR U8663 ( .A(n37914), .B(n37572), .Z(n37574) );
  XNOR U8664 ( .A(n37575), .B(n37227), .Z(n37229) );
  XNOR U8665 ( .A(n37230), .B(n36876), .Z(n36878) );
  XNOR U8666 ( .A(n36879), .B(n36519), .Z(n36521) );
  XNOR U8667 ( .A(n36522), .B(n36156), .Z(n36158) );
  XNOR U8668 ( .A(n36159), .B(n35787), .Z(n35789) );
  XNOR U8669 ( .A(n35790), .B(n35412), .Z(n35414) );
  XNOR U8670 ( .A(n35415), .B(n35031), .Z(n35033) );
  XNOR U8671 ( .A(n35034), .B(n34644), .Z(n34646) );
  XNOR U8672 ( .A(n34647), .B(n34251), .Z(n34253) );
  XNOR U8673 ( .A(n34254), .B(n33852), .Z(n33854) );
  XNOR U8674 ( .A(n33855), .B(n33447), .Z(n33449) );
  XNOR U8675 ( .A(n33450), .B(n33036), .Z(n33038) );
  XNOR U8676 ( .A(n33039), .B(n32619), .Z(n32621) );
  XNOR U8677 ( .A(n32622), .B(n32196), .Z(n32198) );
  XNOR U8678 ( .A(n32199), .B(n31767), .Z(n31769) );
  XNOR U8679 ( .A(n31770), .B(n31332), .Z(n31334) );
  XNOR U8680 ( .A(n31335), .B(n30891), .Z(n30893) );
  XNOR U8681 ( .A(n30894), .B(n30444), .Z(n30446) );
  XNOR U8682 ( .A(n30447), .B(n29991), .Z(n29993) );
  XNOR U8683 ( .A(n29994), .B(n29532), .Z(n29534) );
  XNOR U8684 ( .A(n29535), .B(n29067), .Z(n29069) );
  XNOR U8685 ( .A(n29070), .B(n28596), .Z(n28598) );
  XNOR U8686 ( .A(n28599), .B(n28119), .Z(n28121) );
  XNOR U8687 ( .A(n28122), .B(n27636), .Z(n27638) );
  XNOR U8688 ( .A(n27639), .B(n27147), .Z(n27149) );
  XNOR U8689 ( .A(n27150), .B(n26650), .Z(n26652) );
  XNOR U8690 ( .A(n26653), .B(n26149), .Z(n26151) );
  XNOR U8691 ( .A(n26152), .B(n25641), .Z(n25643) );
  XNOR U8692 ( .A(n25644), .B(n25127), .Z(n25129) );
  XNOR U8693 ( .A(n25130), .B(n24604), .Z(n24606) );
  XNOR U8694 ( .A(n24607), .B(n24079), .Z(n24081) );
  XNOR U8695 ( .A(n24082), .B(n23548), .Z(n23550) );
  XNOR U8696 ( .A(n23551), .B(n23010), .Z(n23012) );
  XNOR U8697 ( .A(n23013), .B(n22466), .Z(n22468) );
  XNOR U8698 ( .A(n22469), .B(n21917), .Z(n21919) );
  XNOR U8699 ( .A(n21920), .B(n21362), .Z(n21364) );
  XNOR U8700 ( .A(n21365), .B(n20800), .Z(n20802) );
  XNOR U8701 ( .A(n20803), .B(n20233), .Z(n20235) );
  XNOR U8702 ( .A(n20236), .B(n19660), .Z(n19662) );
  XNOR U8703 ( .A(n19663), .B(n19081), .Z(n19083) );
  XOR U8704 ( .A(n18389), .B(n18663), .Z(n18393) );
  XOR U8705 ( .A(n17199), .B(n17430), .Z(n17203) );
  XOR U8706 ( .A(n15985), .B(n16216), .Z(n15989) );
  XOR U8707 ( .A(n14119), .B(n14350), .Z(n14123) );
  XOR U8708 ( .A(n14712), .B(n14985), .Z(n14716) );
  XOR U8709 ( .A(n13430), .B(n13727), .Z(n13434) );
  XOR U8710 ( .A(n12122), .B(n12445), .Z(n12126) );
  XOR U8711 ( .A(n12735), .B(n13098), .Z(n12739) );
  XOR U8712 ( .A(n11415), .B(n11802), .Z(n11419) );
  XOR U8713 ( .A(n10073), .B(n10484), .Z(n10077) );
  XOR U8714 ( .A(n10702), .B(n11155), .Z(n10706) );
  XOR U8715 ( .A(n8662), .B(n9151), .Z(n8666) );
  XOR U8716 ( .A(n7227), .B(n7794), .Z(n7231) );
  XOR U8717 ( .A(n5813), .B(n6404), .Z(n5817) );
  XOR U8718 ( .A(n6478), .B(n7111), .Z(n6482) );
  XOR U8719 ( .A(n5050), .B(n5709), .Z(n5054) );
  XOR U8720 ( .A(n4308), .B(n5001), .Z(n4312) );
  XOR U8721 ( .A(n2846), .B(n3563), .Z(n2850) );
  XOR U8722 ( .A(n9353), .B(n9824), .Z(n9357) );
  XOR U8723 ( .A(n7930), .B(n8479), .Z(n7934) );
  XOR U8724 ( .A(n3605), .B(n4280), .Z(n3609) );
  XOR U8725 ( .A(n1365), .B(n2100), .Z(n1369) );
  XOR U8726 ( .A(n5798), .B(n6407), .Z(n5802) );
  XOR U8727 ( .A(n4358), .B(n4991), .Z(n4362) );
  XOR U8728 ( .A(n7257), .B(n7788), .Z(n7261) );
  XOR U8729 ( .A(n5843), .B(n6398), .Z(n5847) );
  XOR U8730 ( .A(n10732), .B(n11149), .Z(n10736) );
  XOR U8731 ( .A(n8692), .B(n9145), .Z(n8696) );
  XOR U8732 ( .A(n12765), .B(n13092), .Z(n12769) );
  XOR U8733 ( .A(n11445), .B(n11796), .Z(n11449) );
  XOR U8734 ( .A(n10103), .B(n10478), .Z(n10107) );
  XOR U8735 ( .A(n14742), .B(n14979), .Z(n14746) );
  XOR U8736 ( .A(n13460), .B(n13721), .Z(n13464) );
  XOR U8737 ( .A(n12152), .B(n12439), .Z(n12156) );
  XNOR U8738 ( .A(n42289), .B(n42037), .Z(n42039) );
  XOR U8739 ( .A(n2901), .B(n3552), .Z(n2905) );
  XOR U8740 ( .A(n7960), .B(n8473), .Z(n7964) );
  XOR U8741 ( .A(n9383), .B(n9818), .Z(n9387) );
  XNOR U8742 ( .A(n43662), .B(n43446), .Z(n43448) );
  XNOR U8743 ( .A(n43449), .B(n43227), .Z(n43229) );
  XNOR U8744 ( .A(n43230), .B(n43002), .Z(n43004) );
  XNOR U8745 ( .A(n43005), .B(n42771), .Z(n42773) );
  XNOR U8746 ( .A(n42774), .B(n42534), .Z(n42536) );
  XNOR U8747 ( .A(n42294), .B(n42042), .Z(n42044) );
  XNOR U8748 ( .A(n42045), .B(n41787), .Z(n41789) );
  XNOR U8749 ( .A(n41790), .B(n41526), .Z(n41528) );
  XNOR U8750 ( .A(n41529), .B(n41259), .Z(n41261) );
  XNOR U8751 ( .A(n41262), .B(n40986), .Z(n40988) );
  XNOR U8752 ( .A(n40989), .B(n40707), .Z(n40709) );
  XNOR U8753 ( .A(n40710), .B(n40422), .Z(n40424) );
  XNOR U8754 ( .A(n40425), .B(n40131), .Z(n40133) );
  XNOR U8755 ( .A(n40134), .B(n39834), .Z(n39836) );
  XNOR U8756 ( .A(n39837), .B(n39531), .Z(n39533) );
  XNOR U8757 ( .A(n39534), .B(n39222), .Z(n39224) );
  XNOR U8758 ( .A(n39225), .B(n38907), .Z(n38909) );
  XNOR U8759 ( .A(n38910), .B(n38586), .Z(n38588) );
  XNOR U8760 ( .A(n38589), .B(n38259), .Z(n38261) );
  XNOR U8761 ( .A(n38262), .B(n37926), .Z(n37928) );
  XNOR U8762 ( .A(n37929), .B(n37587), .Z(n37589) );
  XNOR U8763 ( .A(n37590), .B(n37242), .Z(n37244) );
  XNOR U8764 ( .A(n37245), .B(n36891), .Z(n36893) );
  XNOR U8765 ( .A(n36894), .B(n36534), .Z(n36536) );
  XNOR U8766 ( .A(n36537), .B(n36171), .Z(n36173) );
  XNOR U8767 ( .A(n36174), .B(n35802), .Z(n35804) );
  XNOR U8768 ( .A(n35805), .B(n35427), .Z(n35429) );
  XNOR U8769 ( .A(n35430), .B(n35046), .Z(n35048) );
  XNOR U8770 ( .A(n35049), .B(n34659), .Z(n34661) );
  XNOR U8771 ( .A(n34662), .B(n34266), .Z(n34268) );
  XNOR U8772 ( .A(n34269), .B(n33867), .Z(n33869) );
  XNOR U8773 ( .A(n33870), .B(n33462), .Z(n33464) );
  XNOR U8774 ( .A(n33465), .B(n33051), .Z(n33053) );
  XNOR U8775 ( .A(n33054), .B(n32634), .Z(n32636) );
  XNOR U8776 ( .A(n32637), .B(n32211), .Z(n32213) );
  XNOR U8777 ( .A(n32214), .B(n31782), .Z(n31784) );
  XNOR U8778 ( .A(n31785), .B(n31347), .Z(n31349) );
  XNOR U8779 ( .A(n31350), .B(n30906), .Z(n30908) );
  XNOR U8780 ( .A(n30909), .B(n30459), .Z(n30461) );
  XNOR U8781 ( .A(n30462), .B(n30006), .Z(n30008) );
  XNOR U8782 ( .A(n30009), .B(n29547), .Z(n29549) );
  XNOR U8783 ( .A(n29550), .B(n29082), .Z(n29084) );
  XNOR U8784 ( .A(n29085), .B(n28611), .Z(n28613) );
  XNOR U8785 ( .A(n28614), .B(n28134), .Z(n28136) );
  XNOR U8786 ( .A(n28137), .B(n27651), .Z(n27653) );
  XNOR U8787 ( .A(n27654), .B(n27162), .Z(n27164) );
  XNOR U8788 ( .A(n27165), .B(n26665), .Z(n26667) );
  XNOR U8789 ( .A(n26668), .B(n26164), .Z(n26166) );
  XNOR U8790 ( .A(n26167), .B(n25656), .Z(n25658) );
  XNOR U8791 ( .A(n25659), .B(n25142), .Z(n25144) );
  XNOR U8792 ( .A(n25145), .B(n24619), .Z(n24621) );
  XNOR U8793 ( .A(n24622), .B(n24094), .Z(n24096) );
  XNOR U8794 ( .A(n24097), .B(n23563), .Z(n23565) );
  XNOR U8795 ( .A(n23566), .B(n23025), .Z(n23027) );
  XNOR U8796 ( .A(n23028), .B(n22481), .Z(n22483) );
  XNOR U8797 ( .A(n22484), .B(n21932), .Z(n21934) );
  XNOR U8798 ( .A(n21935), .B(n21377), .Z(n21379) );
  XNOR U8799 ( .A(n21380), .B(n20815), .Z(n20817) );
  XNOR U8800 ( .A(n20818), .B(n20248), .Z(n20250) );
  XNOR U8801 ( .A(n20251), .B(n19675), .Z(n19677) );
  XNOR U8802 ( .A(n19678), .B(n19096), .Z(n19098) );
  XOR U8803 ( .A(n17812), .B(n18025), .Z(n17816) );
  XOR U8804 ( .A(n16610), .B(n16823), .Z(n16614) );
  XOR U8805 ( .A(n15384), .B(n15597), .Z(n15388) );
  XOR U8806 ( .A(n13490), .B(n13715), .Z(n13494) );
  XOR U8807 ( .A(n12182), .B(n12433), .Z(n12186) );
  XOR U8808 ( .A(n12795), .B(n13086), .Z(n12799) );
  XOR U8809 ( .A(n11475), .B(n11790), .Z(n11479) );
  XOR U8810 ( .A(n10133), .B(n10472), .Z(n10137) );
  XOR U8811 ( .A(n10762), .B(n11143), .Z(n10766) );
  XOR U8812 ( .A(n8722), .B(n9139), .Z(n8726) );
  XOR U8813 ( .A(n7287), .B(n7782), .Z(n7291) );
  XOR U8814 ( .A(n5873), .B(n6392), .Z(n5877) );
  XOR U8815 ( .A(n5828), .B(n6401), .Z(n5832) );
  XOR U8816 ( .A(n4388), .B(n4985), .Z(n4392) );
  XOR U8817 ( .A(n4343), .B(n4994), .Z(n4347) );
  XOR U8818 ( .A(n2861), .B(n3560), .Z(n2865) );
  XOR U8819 ( .A(n9413), .B(n9812), .Z(n9417) );
  XOR U8820 ( .A(n7990), .B(n8467), .Z(n7994) );
  XOR U8821 ( .A(n2931), .B(n3546), .Z(n2935) );
  XOR U8822 ( .A(n2886), .B(n3555), .Z(n2890) );
  XOR U8823 ( .A(n1400), .B(n2093), .Z(n1404) );
  XOR U8824 ( .A(n1380), .B(n2097), .Z(n1384) );
  XOR U8825 ( .A(n4373), .B(n4988), .Z(n4377) );
  XOR U8826 ( .A(n5858), .B(n6395), .Z(n5862) );
  XOR U8827 ( .A(n4418), .B(n4979), .Z(n4422) );
  XOR U8828 ( .A(n7317), .B(n7776), .Z(n7321) );
  XOR U8829 ( .A(n5903), .B(n6386), .Z(n5907) );
  XOR U8830 ( .A(n10792), .B(n11137), .Z(n10796) );
  XOR U8831 ( .A(n8752), .B(n9133), .Z(n8756) );
  XOR U8832 ( .A(n12825), .B(n13080), .Z(n12829) );
  XOR U8833 ( .A(n11505), .B(n11784), .Z(n11509) );
  XOR U8834 ( .A(n10163), .B(n10466), .Z(n10167) );
  XOR U8835 ( .A(n12212), .B(n12427), .Z(n12216) );
  XNOR U8836 ( .A(n43015), .B(n42781), .Z(n42783) );
  XOR U8837 ( .A(n2916), .B(n3549), .Z(n2920) );
  XOR U8838 ( .A(n1430), .B(n2087), .Z(n1434) );
  XOR U8839 ( .A(n2961), .B(n3540), .Z(n2965) );
  XOR U8840 ( .A(n8020), .B(n8461), .Z(n8024) );
  XOR U8841 ( .A(n9443), .B(n9806), .Z(n9447) );
  XNOR U8842 ( .A(n44280), .B(n44082), .Z(n44084) );
  XNOR U8843 ( .A(n44085), .B(n43881), .Z(n43883) );
  XNOR U8844 ( .A(n43884), .B(n43674), .Z(n43676) );
  XNOR U8845 ( .A(n43677), .B(n43461), .Z(n43463) );
  XNOR U8846 ( .A(n43464), .B(n43242), .Z(n43244) );
  XNOR U8847 ( .A(n43020), .B(n42786), .Z(n42788) );
  XNOR U8848 ( .A(n42789), .B(n42549), .Z(n42551) );
  XNOR U8849 ( .A(n42552), .B(n42306), .Z(n42308) );
  XNOR U8850 ( .A(n42309), .B(n42057), .Z(n42059) );
  XNOR U8851 ( .A(n42060), .B(n41802), .Z(n41804) );
  XNOR U8852 ( .A(n41805), .B(n41541), .Z(n41543) );
  XNOR U8853 ( .A(n41544), .B(n41274), .Z(n41276) );
  XNOR U8854 ( .A(n41277), .B(n41001), .Z(n41003) );
  XNOR U8855 ( .A(n41004), .B(n40722), .Z(n40724) );
  XNOR U8856 ( .A(n40725), .B(n40437), .Z(n40439) );
  XNOR U8857 ( .A(n40440), .B(n40146), .Z(n40148) );
  XNOR U8858 ( .A(n40149), .B(n39849), .Z(n39851) );
  XNOR U8859 ( .A(n39852), .B(n39546), .Z(n39548) );
  XNOR U8860 ( .A(n39549), .B(n39237), .Z(n39239) );
  XNOR U8861 ( .A(n39240), .B(n38922), .Z(n38924) );
  XNOR U8862 ( .A(n38925), .B(n38601), .Z(n38603) );
  XNOR U8863 ( .A(n38604), .B(n38274), .Z(n38276) );
  XNOR U8864 ( .A(n38277), .B(n37941), .Z(n37943) );
  XNOR U8865 ( .A(n37944), .B(n37602), .Z(n37604) );
  XNOR U8866 ( .A(n37605), .B(n37257), .Z(n37259) );
  XNOR U8867 ( .A(n37260), .B(n36906), .Z(n36908) );
  XNOR U8868 ( .A(n36909), .B(n36549), .Z(n36551) );
  XNOR U8869 ( .A(n36552), .B(n36186), .Z(n36188) );
  XNOR U8870 ( .A(n36189), .B(n35817), .Z(n35819) );
  XNOR U8871 ( .A(n35820), .B(n35442), .Z(n35444) );
  XNOR U8872 ( .A(n35445), .B(n35061), .Z(n35063) );
  XNOR U8873 ( .A(n35064), .B(n34674), .Z(n34676) );
  XNOR U8874 ( .A(n34677), .B(n34281), .Z(n34283) );
  XNOR U8875 ( .A(n34284), .B(n33882), .Z(n33884) );
  XNOR U8876 ( .A(n33885), .B(n33477), .Z(n33479) );
  XNOR U8877 ( .A(n33480), .B(n33066), .Z(n33068) );
  XNOR U8878 ( .A(n33069), .B(n32649), .Z(n32651) );
  XNOR U8879 ( .A(n32652), .B(n32226), .Z(n32228) );
  XNOR U8880 ( .A(n32229), .B(n31797), .Z(n31799) );
  XNOR U8881 ( .A(n31800), .B(n31362), .Z(n31364) );
  XNOR U8882 ( .A(n31365), .B(n30921), .Z(n30923) );
  XNOR U8883 ( .A(n30924), .B(n30474), .Z(n30476) );
  XNOR U8884 ( .A(n30477), .B(n30021), .Z(n30023) );
  XNOR U8885 ( .A(n30024), .B(n29562), .Z(n29564) );
  XNOR U8886 ( .A(n29565), .B(n29097), .Z(n29099) );
  XNOR U8887 ( .A(n29100), .B(n28626), .Z(n28628) );
  XNOR U8888 ( .A(n28629), .B(n28149), .Z(n28151) );
  XNOR U8889 ( .A(n28152), .B(n27666), .Z(n27668) );
  XNOR U8890 ( .A(n27669), .B(n27177), .Z(n27179) );
  XNOR U8891 ( .A(n27180), .B(n26680), .Z(n26682) );
  XNOR U8892 ( .A(n26683), .B(n26179), .Z(n26181) );
  XNOR U8893 ( .A(n26182), .B(n25671), .Z(n25673) );
  XNOR U8894 ( .A(n25674), .B(n25157), .Z(n25159) );
  XNOR U8895 ( .A(n25160), .B(n24634), .Z(n24636) );
  XNOR U8896 ( .A(n24637), .B(n24109), .Z(n24111) );
  XNOR U8897 ( .A(n24112), .B(n23578), .Z(n23580) );
  XNOR U8898 ( .A(n23581), .B(n23040), .Z(n23042) );
  XNOR U8899 ( .A(n23043), .B(n22496), .Z(n22498) );
  XNOR U8900 ( .A(n22499), .B(n21947), .Z(n21949) );
  XNOR U8901 ( .A(n21950), .B(n21392), .Z(n21394) );
  XNOR U8902 ( .A(n21395), .B(n20830), .Z(n20832) );
  XNOR U8903 ( .A(n20833), .B(n20263), .Z(n20265) );
  XNOR U8904 ( .A(n20266), .B(n19690), .Z(n19692) );
  XNOR U8905 ( .A(n19693), .B(n19111), .Z(n19113) );
  XOR U8906 ( .A(n18419), .B(n18651), .Z(n18423) );
  XOR U8907 ( .A(n17229), .B(n17424), .Z(n17233) );
  XOR U8908 ( .A(n16015), .B(n16210), .Z(n16019) );
  XOR U8909 ( .A(n14777), .B(n14972), .Z(n14781) );
  XOR U8910 ( .A(n13515), .B(n13710), .Z(n13519) );
  XOR U8911 ( .A(n12855), .B(n13074), .Z(n12859) );
  XOR U8912 ( .A(n11535), .B(n11778), .Z(n11539) );
  XOR U8913 ( .A(n10193), .B(n10460), .Z(n10197) );
  XOR U8914 ( .A(n10822), .B(n11131), .Z(n10826) );
  XOR U8915 ( .A(n8782), .B(n9127), .Z(n8786) );
  XOR U8916 ( .A(n7347), .B(n7770), .Z(n7351) );
  XOR U8917 ( .A(n5933), .B(n6380), .Z(n5937) );
  XOR U8918 ( .A(n5888), .B(n6389), .Z(n5892) );
  XOR U8919 ( .A(n4448), .B(n4973), .Z(n4452) );
  XOR U8920 ( .A(n4403), .B(n4982), .Z(n4407) );
  XOR U8921 ( .A(n9473), .B(n9800), .Z(n9477) );
  XOR U8922 ( .A(n8050), .B(n8455), .Z(n8054) );
  XOR U8923 ( .A(n2991), .B(n3534), .Z(n2995) );
  XOR U8924 ( .A(n2946), .B(n3543), .Z(n2950) );
  XOR U8925 ( .A(n1460), .B(n2081), .Z(n1464) );
  XOR U8926 ( .A(n1415), .B(n2090), .Z(n1419) );
  XOR U8927 ( .A(n4433), .B(n4976), .Z(n4437) );
  XOR U8928 ( .A(n5918), .B(n6383), .Z(n5922) );
  XOR U8929 ( .A(n4478), .B(n4967), .Z(n4482) );
  XOR U8930 ( .A(n7377), .B(n7764), .Z(n7381) );
  XOR U8931 ( .A(n5963), .B(n6374), .Z(n5967) );
  XOR U8932 ( .A(n10852), .B(n11125), .Z(n10856) );
  XOR U8933 ( .A(n8812), .B(n9121), .Z(n8816) );
  XOR U8934 ( .A(n11565), .B(n11772), .Z(n11569) );
  XOR U8935 ( .A(n10223), .B(n10454), .Z(n10227) );
  XNOR U8936 ( .A(n43687), .B(n43471), .Z(n43473) );
  XOR U8937 ( .A(n1445), .B(n2084), .Z(n1449) );
  XOR U8938 ( .A(n2976), .B(n3537), .Z(n2980) );
  XOR U8939 ( .A(n1490), .B(n2075), .Z(n1494) );
  XOR U8940 ( .A(n3021), .B(n3528), .Z(n3025) );
  XOR U8941 ( .A(n8080), .B(n8449), .Z(n8084) );
  XOR U8942 ( .A(n9503), .B(n9794), .Z(n9507) );
  XNOR U8943 ( .A(n44844), .B(n44664), .Z(n44666) );
  XNOR U8944 ( .A(n44667), .B(n44481), .Z(n44483) );
  XNOR U8945 ( .A(n44484), .B(n44292), .Z(n44294) );
  XNOR U8946 ( .A(n44295), .B(n44097), .Z(n44099) );
  XNOR U8947 ( .A(n44100), .B(n43896), .Z(n43898) );
  XNOR U8948 ( .A(n43692), .B(n43476), .Z(n43478) );
  XNOR U8949 ( .A(n43479), .B(n43257), .Z(n43259) );
  XNOR U8950 ( .A(n43260), .B(n43032), .Z(n43034) );
  XNOR U8951 ( .A(n43035), .B(n42801), .Z(n42803) );
  XNOR U8952 ( .A(n42804), .B(n42564), .Z(n42566) );
  XNOR U8953 ( .A(n42567), .B(n42321), .Z(n42323) );
  XNOR U8954 ( .A(n42324), .B(n42072), .Z(n42074) );
  XNOR U8955 ( .A(n42075), .B(n41817), .Z(n41819) );
  XNOR U8956 ( .A(n41820), .B(n41556), .Z(n41558) );
  XNOR U8957 ( .A(n41559), .B(n41289), .Z(n41291) );
  XNOR U8958 ( .A(n41292), .B(n41016), .Z(n41018) );
  XNOR U8959 ( .A(n41019), .B(n40737), .Z(n40739) );
  XNOR U8960 ( .A(n40740), .B(n40452), .Z(n40454) );
  XNOR U8961 ( .A(n40455), .B(n40161), .Z(n40163) );
  XNOR U8962 ( .A(n40164), .B(n39864), .Z(n39866) );
  XNOR U8963 ( .A(n39867), .B(n39561), .Z(n39563) );
  XNOR U8964 ( .A(n39564), .B(n39252), .Z(n39254) );
  XNOR U8965 ( .A(n39255), .B(n38937), .Z(n38939) );
  XNOR U8966 ( .A(n38940), .B(n38616), .Z(n38618) );
  XNOR U8967 ( .A(n38619), .B(n38289), .Z(n38291) );
  XNOR U8968 ( .A(n38292), .B(n37956), .Z(n37958) );
  XNOR U8969 ( .A(n37959), .B(n37617), .Z(n37619) );
  XNOR U8970 ( .A(n37620), .B(n37272), .Z(n37274) );
  XNOR U8971 ( .A(n37275), .B(n36921), .Z(n36923) );
  XNOR U8972 ( .A(n36924), .B(n36564), .Z(n36566) );
  XNOR U8973 ( .A(n36567), .B(n36201), .Z(n36203) );
  XNOR U8974 ( .A(n36204), .B(n35832), .Z(n35834) );
  XNOR U8975 ( .A(n35835), .B(n35457), .Z(n35459) );
  XNOR U8976 ( .A(n35460), .B(n35076), .Z(n35078) );
  XNOR U8977 ( .A(n35079), .B(n34689), .Z(n34691) );
  XNOR U8978 ( .A(n34692), .B(n34296), .Z(n34298) );
  XNOR U8979 ( .A(n34299), .B(n33897), .Z(n33899) );
  XNOR U8980 ( .A(n33900), .B(n33492), .Z(n33494) );
  XNOR U8981 ( .A(n33495), .B(n33081), .Z(n33083) );
  XNOR U8982 ( .A(n33084), .B(n32664), .Z(n32666) );
  XNOR U8983 ( .A(n32667), .B(n32241), .Z(n32243) );
  XNOR U8984 ( .A(n32244), .B(n31812), .Z(n31814) );
  XNOR U8985 ( .A(n31815), .B(n31377), .Z(n31379) );
  XNOR U8986 ( .A(n31380), .B(n30936), .Z(n30938) );
  XNOR U8987 ( .A(n30939), .B(n30489), .Z(n30491) );
  XNOR U8988 ( .A(n30492), .B(n30036), .Z(n30038) );
  XNOR U8989 ( .A(n30039), .B(n29577), .Z(n29579) );
  XNOR U8990 ( .A(n29580), .B(n29112), .Z(n29114) );
  XNOR U8991 ( .A(n29115), .B(n28641), .Z(n28643) );
  XNOR U8992 ( .A(n28644), .B(n28164), .Z(n28166) );
  XNOR U8993 ( .A(n28167), .B(n27681), .Z(n27683) );
  XNOR U8994 ( .A(n27684), .B(n27192), .Z(n27194) );
  XNOR U8995 ( .A(n27195), .B(n26695), .Z(n26697) );
  XNOR U8996 ( .A(n26698), .B(n26194), .Z(n26196) );
  XNOR U8997 ( .A(n26197), .B(n25686), .Z(n25688) );
  XNOR U8998 ( .A(n25689), .B(n25172), .Z(n25174) );
  XNOR U8999 ( .A(n25175), .B(n24649), .Z(n24651) );
  XNOR U9000 ( .A(n24652), .B(n24124), .Z(n24126) );
  XNOR U9001 ( .A(n24127), .B(n23593), .Z(n23595) );
  XNOR U9002 ( .A(n23596), .B(n23055), .Z(n23057) );
  XNOR U9003 ( .A(n23058), .B(n22511), .Z(n22513) );
  XNOR U9004 ( .A(n22514), .B(n21962), .Z(n21964) );
  XNOR U9005 ( .A(n21965), .B(n21407), .Z(n21409) );
  XNOR U9006 ( .A(n21410), .B(n20845), .Z(n20847) );
  XNOR U9007 ( .A(n20848), .B(n20278), .Z(n20280) );
  XNOR U9008 ( .A(n20281), .B(n19705), .Z(n19707) );
  XNOR U9009 ( .A(n19708), .B(n19126), .Z(n19128) );
  XOR U9010 ( .A(n17842), .B(n18019), .Z(n17846) );
  XOR U9011 ( .A(n16640), .B(n16817), .Z(n16644) );
  XOR U9012 ( .A(n15414), .B(n15591), .Z(n15418) );
  XOR U9013 ( .A(n14164), .B(n14341), .Z(n14168) );
  XOR U9014 ( .A(n12890), .B(n13067), .Z(n12894) );
  XOR U9015 ( .A(n11590), .B(n11767), .Z(n11594) );
  XOR U9016 ( .A(n10253), .B(n10448), .Z(n10257) );
  XOR U9017 ( .A(n10882), .B(n11119), .Z(n10886) );
  XOR U9018 ( .A(n8842), .B(n9115), .Z(n8846) );
  XOR U9019 ( .A(n7407), .B(n7758), .Z(n7411) );
  XOR U9020 ( .A(n5993), .B(n6368), .Z(n5997) );
  XOR U9021 ( .A(n5948), .B(n6377), .Z(n5952) );
  XOR U9022 ( .A(n4508), .B(n4961), .Z(n4512) );
  XOR U9023 ( .A(n4463), .B(n4970), .Z(n4467) );
  XOR U9024 ( .A(n9533), .B(n9788), .Z(n9537) );
  XOR U9025 ( .A(n8110), .B(n8443), .Z(n8114) );
  XOR U9026 ( .A(n3051), .B(n3522), .Z(n3055) );
  XOR U9027 ( .A(n3006), .B(n3531), .Z(n3010) );
  XOR U9028 ( .A(n1520), .B(n2069), .Z(n1524) );
  XOR U9029 ( .A(n1475), .B(n2078), .Z(n1479) );
  XOR U9030 ( .A(n4493), .B(n4964), .Z(n4497) );
  XOR U9031 ( .A(n5978), .B(n6371), .Z(n5982) );
  XOR U9032 ( .A(n4538), .B(n4955), .Z(n4542) );
  XOR U9033 ( .A(n7437), .B(n7752), .Z(n7441) );
  XOR U9034 ( .A(n6023), .B(n6362), .Z(n6027) );
  XOR U9035 ( .A(n10912), .B(n11113), .Z(n10916) );
  XOR U9036 ( .A(n8872), .B(n9109), .Z(n8876) );
  XNOR U9037 ( .A(n44305), .B(n44107), .Z(n44109) );
  XOR U9038 ( .A(n1505), .B(n2072), .Z(n1509) );
  XOR U9039 ( .A(n3036), .B(n3525), .Z(n3040) );
  XOR U9040 ( .A(n1550), .B(n2063), .Z(n1554) );
  XOR U9041 ( .A(n3081), .B(n3516), .Z(n3085) );
  XOR U9042 ( .A(n8140), .B(n8437), .Z(n8144) );
  XOR U9043 ( .A(n9563), .B(n9782), .Z(n9567) );
  XNOR U9044 ( .A(n45354), .B(n45192), .Z(n45194) );
  XNOR U9045 ( .A(n45195), .B(n45027), .Z(n45029) );
  XNOR U9046 ( .A(n45030), .B(n44856), .Z(n44858) );
  XNOR U9047 ( .A(n44859), .B(n44679), .Z(n44681) );
  XNOR U9048 ( .A(n44682), .B(n44496), .Z(n44498) );
  XNOR U9049 ( .A(n44310), .B(n44112), .Z(n44114) );
  XNOR U9050 ( .A(n44115), .B(n43911), .Z(n43913) );
  XNOR U9051 ( .A(n43914), .B(n43704), .Z(n43706) );
  XNOR U9052 ( .A(n43707), .B(n43491), .Z(n43493) );
  XNOR U9053 ( .A(n43494), .B(n43272), .Z(n43274) );
  XNOR U9054 ( .A(n43275), .B(n43047), .Z(n43049) );
  XNOR U9055 ( .A(n43050), .B(n42816), .Z(n42818) );
  XNOR U9056 ( .A(n42819), .B(n42579), .Z(n42581) );
  XNOR U9057 ( .A(n42582), .B(n42336), .Z(n42338) );
  XNOR U9058 ( .A(n42339), .B(n42087), .Z(n42089) );
  XNOR U9059 ( .A(n42090), .B(n41832), .Z(n41834) );
  XNOR U9060 ( .A(n41835), .B(n41571), .Z(n41573) );
  XNOR U9061 ( .A(n41574), .B(n41304), .Z(n41306) );
  XNOR U9062 ( .A(n41307), .B(n41031), .Z(n41033) );
  XNOR U9063 ( .A(n41034), .B(n40752), .Z(n40754) );
  XNOR U9064 ( .A(n40755), .B(n40467), .Z(n40469) );
  XNOR U9065 ( .A(n40470), .B(n40176), .Z(n40178) );
  XNOR U9066 ( .A(n40179), .B(n39879), .Z(n39881) );
  XNOR U9067 ( .A(n39882), .B(n39576), .Z(n39578) );
  XNOR U9068 ( .A(n39579), .B(n39267), .Z(n39269) );
  XNOR U9069 ( .A(n39270), .B(n38952), .Z(n38954) );
  XNOR U9070 ( .A(n38955), .B(n38631), .Z(n38633) );
  XNOR U9071 ( .A(n38634), .B(n38304), .Z(n38306) );
  XNOR U9072 ( .A(n38307), .B(n37971), .Z(n37973) );
  XNOR U9073 ( .A(n37974), .B(n37632), .Z(n37634) );
  XNOR U9074 ( .A(n37635), .B(n37287), .Z(n37289) );
  XNOR U9075 ( .A(n37290), .B(n36936), .Z(n36938) );
  XNOR U9076 ( .A(n36939), .B(n36579), .Z(n36581) );
  XNOR U9077 ( .A(n36582), .B(n36216), .Z(n36218) );
  XNOR U9078 ( .A(n36219), .B(n35847), .Z(n35849) );
  XNOR U9079 ( .A(n35850), .B(n35472), .Z(n35474) );
  XNOR U9080 ( .A(n35475), .B(n35091), .Z(n35093) );
  XNOR U9081 ( .A(n35094), .B(n34704), .Z(n34706) );
  XNOR U9082 ( .A(n34707), .B(n34311), .Z(n34313) );
  XNOR U9083 ( .A(n34314), .B(n33912), .Z(n33914) );
  XNOR U9084 ( .A(n33915), .B(n33507), .Z(n33509) );
  XNOR U9085 ( .A(n33510), .B(n33096), .Z(n33098) );
  XNOR U9086 ( .A(n33099), .B(n32679), .Z(n32681) );
  XNOR U9087 ( .A(n32682), .B(n32256), .Z(n32258) );
  XNOR U9088 ( .A(n32259), .B(n31827), .Z(n31829) );
  XNOR U9089 ( .A(n31830), .B(n31392), .Z(n31394) );
  XNOR U9090 ( .A(n31395), .B(n30951), .Z(n30953) );
  XNOR U9091 ( .A(n30954), .B(n30504), .Z(n30506) );
  XNOR U9092 ( .A(n30507), .B(n30051), .Z(n30053) );
  XNOR U9093 ( .A(n30054), .B(n29592), .Z(n29594) );
  XNOR U9094 ( .A(n29595), .B(n29127), .Z(n29129) );
  XNOR U9095 ( .A(n29130), .B(n28656), .Z(n28658) );
  XNOR U9096 ( .A(n28659), .B(n28179), .Z(n28181) );
  XNOR U9097 ( .A(n28182), .B(n27696), .Z(n27698) );
  XNOR U9098 ( .A(n27699), .B(n27207), .Z(n27209) );
  XNOR U9099 ( .A(n27210), .B(n26710), .Z(n26712) );
  XNOR U9100 ( .A(n26713), .B(n26209), .Z(n26211) );
  XNOR U9101 ( .A(n26212), .B(n25701), .Z(n25703) );
  XNOR U9102 ( .A(n25704), .B(n25187), .Z(n25189) );
  XNOR U9103 ( .A(n25190), .B(n24664), .Z(n24666) );
  XNOR U9104 ( .A(n24667), .B(n24139), .Z(n24141) );
  XNOR U9105 ( .A(n24142), .B(n23608), .Z(n23610) );
  XNOR U9106 ( .A(n23611), .B(n23070), .Z(n23072) );
  XNOR U9107 ( .A(n23073), .B(n22526), .Z(n22528) );
  XNOR U9108 ( .A(n22529), .B(n21977), .Z(n21979) );
  XNOR U9109 ( .A(n21980), .B(n21422), .Z(n21424) );
  XNOR U9110 ( .A(n21425), .B(n20860), .Z(n20862) );
  XNOR U9111 ( .A(n20863), .B(n20293), .Z(n20295) );
  XNOR U9112 ( .A(n20296), .B(n19720), .Z(n19722) );
  XNOR U9113 ( .A(n19723), .B(n19141), .Z(n19143) );
  XOR U9114 ( .A(n18449), .B(n18639), .Z(n18453) );
  XOR U9115 ( .A(n17259), .B(n17418), .Z(n17263) );
  XOR U9116 ( .A(n16045), .B(n16204), .Z(n16049) );
  XOR U9117 ( .A(n14807), .B(n14966), .Z(n14811) );
  XOR U9118 ( .A(n13545), .B(n13704), .Z(n13549) );
  XOR U9119 ( .A(n12257), .B(n12418), .Z(n12261) );
  XOR U9120 ( .A(n10942), .B(n11107), .Z(n10946) );
  XOR U9121 ( .A(n8902), .B(n9103), .Z(n8906) );
  XOR U9122 ( .A(n7467), .B(n7746), .Z(n7471) );
  XOR U9123 ( .A(n6053), .B(n6356), .Z(n6057) );
  XOR U9124 ( .A(n6008), .B(n6365), .Z(n6012) );
  XOR U9125 ( .A(n4568), .B(n4949), .Z(n4572) );
  XOR U9126 ( .A(n4523), .B(n4958), .Z(n4527) );
  XOR U9127 ( .A(n9593), .B(n9776), .Z(n9597) );
  XOR U9128 ( .A(n8170), .B(n8431), .Z(n8174) );
  XOR U9129 ( .A(n3111), .B(n3510), .Z(n3115) );
  XOR U9130 ( .A(n3066), .B(n3519), .Z(n3070) );
  XOR U9131 ( .A(n1580), .B(n2057), .Z(n1584) );
  XOR U9132 ( .A(n1535), .B(n2066), .Z(n1539) );
  XOR U9133 ( .A(n4553), .B(n4952), .Z(n4557) );
  XOR U9134 ( .A(n6038), .B(n6359), .Z(n6042) );
  XOR U9135 ( .A(n4598), .B(n4943), .Z(n4602) );
  XOR U9136 ( .A(n7497), .B(n7740), .Z(n7501) );
  XOR U9137 ( .A(n6083), .B(n6350), .Z(n6087) );
  XOR U9138 ( .A(n8932), .B(n9097), .Z(n8936) );
  XNOR U9139 ( .A(n44869), .B(n44689), .Z(n44691) );
  XOR U9140 ( .A(n10957), .B(n11104), .Z(n10961) );
  XOR U9141 ( .A(n1565), .B(n2060), .Z(n1569) );
  XOR U9142 ( .A(n3096), .B(n3513), .Z(n3100) );
  XOR U9143 ( .A(n1610), .B(n2051), .Z(n1614) );
  XOR U9144 ( .A(n3141), .B(n3504), .Z(n3145) );
  XOR U9145 ( .A(n8200), .B(n8425), .Z(n8204) );
  XOR U9146 ( .A(n9623), .B(n9770), .Z(n9627) );
  XNOR U9147 ( .A(n45810), .B(n45666), .Z(n45668) );
  XNOR U9148 ( .A(n45669), .B(n45519), .Z(n45521) );
  XNOR U9149 ( .A(n45522), .B(n45366), .Z(n45368) );
  XNOR U9150 ( .A(n45369), .B(n45207), .Z(n45209) );
  XNOR U9151 ( .A(n45210), .B(n45042), .Z(n45044) );
  XNOR U9152 ( .A(n44874), .B(n44694), .Z(n44696) );
  XNOR U9153 ( .A(n44697), .B(n44511), .Z(n44513) );
  XNOR U9154 ( .A(n44514), .B(n44322), .Z(n44324) );
  XNOR U9155 ( .A(n44325), .B(n44127), .Z(n44129) );
  XNOR U9156 ( .A(n44130), .B(n43926), .Z(n43928) );
  XNOR U9157 ( .A(n43929), .B(n43719), .Z(n43721) );
  XNOR U9158 ( .A(n43722), .B(n43506), .Z(n43508) );
  XNOR U9159 ( .A(n43509), .B(n43287), .Z(n43289) );
  XNOR U9160 ( .A(n43290), .B(n43062), .Z(n43064) );
  XNOR U9161 ( .A(n43065), .B(n42831), .Z(n42833) );
  XNOR U9162 ( .A(n42834), .B(n42594), .Z(n42596) );
  XNOR U9163 ( .A(n42597), .B(n42351), .Z(n42353) );
  XNOR U9164 ( .A(n42354), .B(n42102), .Z(n42104) );
  XNOR U9165 ( .A(n42105), .B(n41847), .Z(n41849) );
  XNOR U9166 ( .A(n41850), .B(n41586), .Z(n41588) );
  XNOR U9167 ( .A(n41589), .B(n41319), .Z(n41321) );
  XNOR U9168 ( .A(n41322), .B(n41046), .Z(n41048) );
  XNOR U9169 ( .A(n41049), .B(n40767), .Z(n40769) );
  XNOR U9170 ( .A(n40770), .B(n40482), .Z(n40484) );
  XNOR U9171 ( .A(n40485), .B(n40191), .Z(n40193) );
  XNOR U9172 ( .A(n40194), .B(n39894), .Z(n39896) );
  XNOR U9173 ( .A(n39897), .B(n39591), .Z(n39593) );
  XNOR U9174 ( .A(n39594), .B(n39282), .Z(n39284) );
  XNOR U9175 ( .A(n39285), .B(n38967), .Z(n38969) );
  XNOR U9176 ( .A(n38970), .B(n38646), .Z(n38648) );
  XNOR U9177 ( .A(n38649), .B(n38319), .Z(n38321) );
  XNOR U9178 ( .A(n38322), .B(n37986), .Z(n37988) );
  XNOR U9179 ( .A(n37989), .B(n37647), .Z(n37649) );
  XNOR U9180 ( .A(n37650), .B(n37302), .Z(n37304) );
  XNOR U9181 ( .A(n37305), .B(n36951), .Z(n36953) );
  XNOR U9182 ( .A(n36954), .B(n36594), .Z(n36596) );
  XNOR U9183 ( .A(n36597), .B(n36231), .Z(n36233) );
  XNOR U9184 ( .A(n36234), .B(n35862), .Z(n35864) );
  XNOR U9185 ( .A(n35865), .B(n35487), .Z(n35489) );
  XNOR U9186 ( .A(n35490), .B(n35106), .Z(n35108) );
  XNOR U9187 ( .A(n35109), .B(n34719), .Z(n34721) );
  XNOR U9188 ( .A(n34722), .B(n34326), .Z(n34328) );
  XNOR U9189 ( .A(n34329), .B(n33927), .Z(n33929) );
  XNOR U9190 ( .A(n33930), .B(n33522), .Z(n33524) );
  XNOR U9191 ( .A(n33525), .B(n33111), .Z(n33113) );
  XNOR U9192 ( .A(n33114), .B(n32694), .Z(n32696) );
  XNOR U9193 ( .A(n32697), .B(n32271), .Z(n32273) );
  XNOR U9194 ( .A(n32274), .B(n31842), .Z(n31844) );
  XNOR U9195 ( .A(n31845), .B(n31407), .Z(n31409) );
  XNOR U9196 ( .A(n31410), .B(n30966), .Z(n30968) );
  XNOR U9197 ( .A(n30969), .B(n30519), .Z(n30521) );
  XNOR U9198 ( .A(n30522), .B(n30066), .Z(n30068) );
  XNOR U9199 ( .A(n30069), .B(n29607), .Z(n29609) );
  XNOR U9200 ( .A(n29610), .B(n29142), .Z(n29144) );
  XNOR U9201 ( .A(n29145), .B(n28671), .Z(n28673) );
  XNOR U9202 ( .A(n28674), .B(n28194), .Z(n28196) );
  XNOR U9203 ( .A(n28197), .B(n27711), .Z(n27713) );
  XNOR U9204 ( .A(n27714), .B(n27222), .Z(n27224) );
  XNOR U9205 ( .A(n27225), .B(n26725), .Z(n26727) );
  XNOR U9206 ( .A(n26728), .B(n26224), .Z(n26226) );
  XNOR U9207 ( .A(n26227), .B(n25716), .Z(n25718) );
  XNOR U9208 ( .A(n25719), .B(n25202), .Z(n25204) );
  XNOR U9209 ( .A(n25205), .B(n24679), .Z(n24681) );
  XNOR U9210 ( .A(n24682), .B(n24154), .Z(n24156) );
  XNOR U9211 ( .A(n24157), .B(n23623), .Z(n23625) );
  XNOR U9212 ( .A(n23626), .B(n23085), .Z(n23087) );
  XNOR U9213 ( .A(n23088), .B(n22541), .Z(n22543) );
  XNOR U9214 ( .A(n22544), .B(n21992), .Z(n21994) );
  XNOR U9215 ( .A(n21995), .B(n21437), .Z(n21439) );
  XNOR U9216 ( .A(n21440), .B(n20875), .Z(n20877) );
  XNOR U9217 ( .A(n20878), .B(n20308), .Z(n20310) );
  XNOR U9218 ( .A(n20311), .B(n19735), .Z(n19737) );
  XNOR U9219 ( .A(n19738), .B(n19156), .Z(n19158) );
  XOR U9220 ( .A(n18464), .B(n18633), .Z(n18468) );
  XOR U9221 ( .A(n17274), .B(n17415), .Z(n17278) );
  XOR U9222 ( .A(n16060), .B(n16201), .Z(n16064) );
  XOR U9223 ( .A(n14822), .B(n14963), .Z(n14826) );
  XOR U9224 ( .A(n13560), .B(n13701), .Z(n13564) );
  XOR U9225 ( .A(n12272), .B(n12415), .Z(n12276) );
  XOR U9226 ( .A(n7527), .B(n7734), .Z(n7531) );
  XOR U9227 ( .A(n6113), .B(n6344), .Z(n6117) );
  XOR U9228 ( .A(n6068), .B(n6353), .Z(n6072) );
  XOR U9229 ( .A(n4628), .B(n4937), .Z(n4632) );
  XOR U9230 ( .A(n4583), .B(n4946), .Z(n4587) );
  XOR U9231 ( .A(n8230), .B(n8419), .Z(n8234) );
  XOR U9232 ( .A(n3171), .B(n3498), .Z(n3175) );
  XOR U9233 ( .A(n3126), .B(n3507), .Z(n3130) );
  XOR U9234 ( .A(n1640), .B(n2045), .Z(n1644) );
  XOR U9235 ( .A(n1595), .B(n2054), .Z(n1599) );
  XOR U9236 ( .A(n4613), .B(n4940), .Z(n4617) );
  XOR U9237 ( .A(n6098), .B(n6347), .Z(n6102) );
  XOR U9238 ( .A(n4658), .B(n4931), .Z(n4662) );
  XOR U9239 ( .A(n7557), .B(n7728), .Z(n7561) );
  XOR U9240 ( .A(n6143), .B(n6338), .Z(n6147) );
  XNOR U9241 ( .A(n45379), .B(n45217), .Z(n45219) );
  XOR U9242 ( .A(n11630), .B(n11759), .Z(n11634) );
  XOR U9243 ( .A(n10308), .B(n10437), .Z(n10312) );
  XOR U9244 ( .A(n8962), .B(n9091), .Z(n8966) );
  XOR U9245 ( .A(n1625), .B(n2048), .Z(n1629) );
  XOR U9246 ( .A(n3156), .B(n3501), .Z(n3160) );
  XOR U9247 ( .A(n1670), .B(n2039), .Z(n1674) );
  XOR U9248 ( .A(n3201), .B(n3492), .Z(n3205) );
  XOR U9249 ( .A(n8260), .B(n8413), .Z(n8264) );
  XNOR U9250 ( .A(n46212), .B(n46086), .Z(n46088) );
  XNOR U9251 ( .A(n46089), .B(n45957), .Z(n45959) );
  XNOR U9252 ( .A(n45960), .B(n45822), .Z(n45824) );
  XNOR U9253 ( .A(n45825), .B(n45681), .Z(n45683) );
  XNOR U9254 ( .A(n45684), .B(n45534), .Z(n45536) );
  XNOR U9255 ( .A(n45384), .B(n45222), .Z(n45224) );
  XNOR U9256 ( .A(n45225), .B(n45057), .Z(n45059) );
  XNOR U9257 ( .A(n45060), .B(n44886), .Z(n44888) );
  XNOR U9258 ( .A(n44889), .B(n44709), .Z(n44711) );
  XNOR U9259 ( .A(n44712), .B(n44526), .Z(n44528) );
  XNOR U9260 ( .A(n44529), .B(n44337), .Z(n44339) );
  XNOR U9261 ( .A(n44340), .B(n44142), .Z(n44144) );
  XNOR U9262 ( .A(n44145), .B(n43941), .Z(n43943) );
  XNOR U9263 ( .A(n43944), .B(n43734), .Z(n43736) );
  XNOR U9264 ( .A(n43737), .B(n43521), .Z(n43523) );
  XNOR U9265 ( .A(n43524), .B(n43302), .Z(n43304) );
  XNOR U9266 ( .A(n43305), .B(n43077), .Z(n43079) );
  XNOR U9267 ( .A(n43080), .B(n42846), .Z(n42848) );
  XNOR U9268 ( .A(n42849), .B(n42609), .Z(n42611) );
  XNOR U9269 ( .A(n42612), .B(n42366), .Z(n42368) );
  XNOR U9270 ( .A(n42369), .B(n42117), .Z(n42119) );
  XNOR U9271 ( .A(n42120), .B(n41862), .Z(n41864) );
  XNOR U9272 ( .A(n41865), .B(n41601), .Z(n41603) );
  XNOR U9273 ( .A(n41604), .B(n41334), .Z(n41336) );
  XNOR U9274 ( .A(n41337), .B(n41061), .Z(n41063) );
  XNOR U9275 ( .A(n41064), .B(n40782), .Z(n40784) );
  XNOR U9276 ( .A(n40785), .B(n40497), .Z(n40499) );
  XNOR U9277 ( .A(n40500), .B(n40206), .Z(n40208) );
  XNOR U9278 ( .A(n40209), .B(n39909), .Z(n39911) );
  XNOR U9279 ( .A(n39912), .B(n39606), .Z(n39608) );
  XNOR U9280 ( .A(n39609), .B(n39297), .Z(n39299) );
  XNOR U9281 ( .A(n39300), .B(n38982), .Z(n38984) );
  XNOR U9282 ( .A(n38985), .B(n38661), .Z(n38663) );
  XNOR U9283 ( .A(n38664), .B(n38334), .Z(n38336) );
  XNOR U9284 ( .A(n38337), .B(n38001), .Z(n38003) );
  XNOR U9285 ( .A(n38004), .B(n37662), .Z(n37664) );
  XNOR U9286 ( .A(n37665), .B(n37317), .Z(n37319) );
  XNOR U9287 ( .A(n37320), .B(n36966), .Z(n36968) );
  XNOR U9288 ( .A(n36969), .B(n36609), .Z(n36611) );
  XNOR U9289 ( .A(n36612), .B(n36246), .Z(n36248) );
  XNOR U9290 ( .A(n36249), .B(n35877), .Z(n35879) );
  XNOR U9291 ( .A(n35880), .B(n35502), .Z(n35504) );
  XNOR U9292 ( .A(n35505), .B(n35121), .Z(n35123) );
  XNOR U9293 ( .A(n35124), .B(n34734), .Z(n34736) );
  XNOR U9294 ( .A(n34737), .B(n34341), .Z(n34343) );
  XNOR U9295 ( .A(n34344), .B(n33942), .Z(n33944) );
  XNOR U9296 ( .A(n33945), .B(n33537), .Z(n33539) );
  XNOR U9297 ( .A(n33540), .B(n33126), .Z(n33128) );
  XNOR U9298 ( .A(n33129), .B(n32709), .Z(n32711) );
  XNOR U9299 ( .A(n32712), .B(n32286), .Z(n32288) );
  XNOR U9300 ( .A(n32289), .B(n31857), .Z(n31859) );
  XNOR U9301 ( .A(n31860), .B(n31422), .Z(n31424) );
  XNOR U9302 ( .A(n31425), .B(n30981), .Z(n30983) );
  XNOR U9303 ( .A(n30984), .B(n30534), .Z(n30536) );
  XNOR U9304 ( .A(n30537), .B(n30081), .Z(n30083) );
  XNOR U9305 ( .A(n30084), .B(n29622), .Z(n29624) );
  XNOR U9306 ( .A(n29625), .B(n29157), .Z(n29159) );
  XNOR U9307 ( .A(n29160), .B(n28686), .Z(n28688) );
  XNOR U9308 ( .A(n28689), .B(n28209), .Z(n28211) );
  XNOR U9309 ( .A(n28212), .B(n27726), .Z(n27728) );
  XNOR U9310 ( .A(n27729), .B(n27237), .Z(n27239) );
  XNOR U9311 ( .A(n27240), .B(n26740), .Z(n26742) );
  XNOR U9312 ( .A(n26743), .B(n26239), .Z(n26241) );
  XNOR U9313 ( .A(n26242), .B(n25731), .Z(n25733) );
  XNOR U9314 ( .A(n25734), .B(n25217), .Z(n25219) );
  XNOR U9315 ( .A(n25220), .B(n24694), .Z(n24696) );
  XNOR U9316 ( .A(n24697), .B(n24169), .Z(n24171) );
  XNOR U9317 ( .A(n24172), .B(n23638), .Z(n23640) );
  XNOR U9318 ( .A(n23641), .B(n23100), .Z(n23102) );
  XNOR U9319 ( .A(n23103), .B(n22556), .Z(n22558) );
  XNOR U9320 ( .A(n22559), .B(n22007), .Z(n22009) );
  XNOR U9321 ( .A(n22010), .B(n21452), .Z(n21454) );
  XNOR U9322 ( .A(n21455), .B(n20890), .Z(n20892) );
  XNOR U9323 ( .A(n20893), .B(n20323), .Z(n20325) );
  XNOR U9324 ( .A(n20326), .B(n19750), .Z(n19752) );
  XNOR U9325 ( .A(n19753), .B(n19171), .Z(n19173) );
  XOR U9326 ( .A(n18479), .B(n18627), .Z(n18483) );
  XOR U9327 ( .A(n17289), .B(n17412), .Z(n17293) );
  XOR U9328 ( .A(n16075), .B(n16198), .Z(n16079) );
  XOR U9329 ( .A(n14837), .B(n14960), .Z(n14841) );
  XOR U9330 ( .A(n13575), .B(n13698), .Z(n13579) );
  XOR U9331 ( .A(n7587), .B(n7722), .Z(n7591) );
  XOR U9332 ( .A(n6173), .B(n6332), .Z(n6177) );
  XOR U9333 ( .A(n6128), .B(n6341), .Z(n6132) );
  XOR U9334 ( .A(n4688), .B(n4925), .Z(n4692) );
  XOR U9335 ( .A(n4643), .B(n4934), .Z(n4647) );
  XOR U9336 ( .A(n3231), .B(n3486), .Z(n3235) );
  XOR U9337 ( .A(n3186), .B(n3495), .Z(n3190) );
  XOR U9338 ( .A(n1700), .B(n2033), .Z(n1704) );
  XOR U9339 ( .A(n1655), .B(n2042), .Z(n1659) );
  XOR U9340 ( .A(n4673), .B(n4928), .Z(n4677) );
  XOR U9341 ( .A(n6158), .B(n6335), .Z(n6162) );
  XOR U9342 ( .A(n4718), .B(n4919), .Z(n4722) );
  XNOR U9343 ( .A(n45835), .B(n45691), .Z(n45693) );
  XOR U9344 ( .A(n12945), .B(n13056), .Z(n12949) );
  XOR U9345 ( .A(n11645), .B(n11756), .Z(n11649) );
  XOR U9346 ( .A(n10323), .B(n10434), .Z(n10327) );
  XOR U9347 ( .A(n6913), .B(n7024), .Z(n6917) );
  XOR U9348 ( .A(n1685), .B(n2036), .Z(n1689) );
  XOR U9349 ( .A(n3216), .B(n3489), .Z(n3220) );
  XOR U9350 ( .A(n1730), .B(n2027), .Z(n1734) );
  XOR U9351 ( .A(n3261), .B(n3480), .Z(n3265) );
  XNOR U9352 ( .A(n46560), .B(n46452), .Z(n46454) );
  XNOR U9353 ( .A(n46455), .B(n46341), .Z(n46343) );
  XNOR U9354 ( .A(n46344), .B(n46224), .Z(n46226) );
  XNOR U9355 ( .A(n46227), .B(n46101), .Z(n46103) );
  XNOR U9356 ( .A(n46104), .B(n45972), .Z(n45974) );
  XNOR U9357 ( .A(n45840), .B(n45696), .Z(n45698) );
  XNOR U9358 ( .A(n45699), .B(n45549), .Z(n45551) );
  XNOR U9359 ( .A(n45552), .B(n45396), .Z(n45398) );
  XNOR U9360 ( .A(n45399), .B(n45237), .Z(n45239) );
  XNOR U9361 ( .A(n45240), .B(n45072), .Z(n45074) );
  XNOR U9362 ( .A(n45075), .B(n44901), .Z(n44903) );
  XNOR U9363 ( .A(n44904), .B(n44724), .Z(n44726) );
  XNOR U9364 ( .A(n44727), .B(n44541), .Z(n44543) );
  XNOR U9365 ( .A(n44544), .B(n44352), .Z(n44354) );
  XNOR U9366 ( .A(n44355), .B(n44157), .Z(n44159) );
  XNOR U9367 ( .A(n44160), .B(n43956), .Z(n43958) );
  XNOR U9368 ( .A(n43959), .B(n43749), .Z(n43751) );
  XNOR U9369 ( .A(n43752), .B(n43536), .Z(n43538) );
  XNOR U9370 ( .A(n43539), .B(n43317), .Z(n43319) );
  XNOR U9371 ( .A(n43320), .B(n43092), .Z(n43094) );
  XNOR U9372 ( .A(n43095), .B(n42861), .Z(n42863) );
  XNOR U9373 ( .A(n42864), .B(n42624), .Z(n42626) );
  XNOR U9374 ( .A(n42627), .B(n42381), .Z(n42383) );
  XNOR U9375 ( .A(n42384), .B(n42132), .Z(n42134) );
  XNOR U9376 ( .A(n42135), .B(n41877), .Z(n41879) );
  XNOR U9377 ( .A(n41880), .B(n41616), .Z(n41618) );
  XNOR U9378 ( .A(n41619), .B(n41349), .Z(n41351) );
  XNOR U9379 ( .A(n41352), .B(n41076), .Z(n41078) );
  XNOR U9380 ( .A(n41079), .B(n40797), .Z(n40799) );
  XNOR U9381 ( .A(n40800), .B(n40512), .Z(n40514) );
  XNOR U9382 ( .A(n40515), .B(n40221), .Z(n40223) );
  XNOR U9383 ( .A(n40224), .B(n39924), .Z(n39926) );
  XNOR U9384 ( .A(n39927), .B(n39621), .Z(n39623) );
  XNOR U9385 ( .A(n39624), .B(n39312), .Z(n39314) );
  XNOR U9386 ( .A(n39315), .B(n38997), .Z(n38999) );
  XNOR U9387 ( .A(n39000), .B(n38676), .Z(n38678) );
  XNOR U9388 ( .A(n38679), .B(n38349), .Z(n38351) );
  XNOR U9389 ( .A(n38352), .B(n38016), .Z(n38018) );
  XNOR U9390 ( .A(n38019), .B(n37677), .Z(n37679) );
  XNOR U9391 ( .A(n37680), .B(n37332), .Z(n37334) );
  XNOR U9392 ( .A(n37335), .B(n36981), .Z(n36983) );
  XNOR U9393 ( .A(n36984), .B(n36624), .Z(n36626) );
  XNOR U9394 ( .A(n36627), .B(n36261), .Z(n36263) );
  XNOR U9395 ( .A(n36264), .B(n35892), .Z(n35894) );
  XNOR U9396 ( .A(n35895), .B(n35517), .Z(n35519) );
  XNOR U9397 ( .A(n35520), .B(n35136), .Z(n35138) );
  XNOR U9398 ( .A(n35139), .B(n34749), .Z(n34751) );
  XNOR U9399 ( .A(n34752), .B(n34356), .Z(n34358) );
  XNOR U9400 ( .A(n34359), .B(n33957), .Z(n33959) );
  XNOR U9401 ( .A(n33960), .B(n33552), .Z(n33554) );
  XNOR U9402 ( .A(n33555), .B(n33141), .Z(n33143) );
  XNOR U9403 ( .A(n33144), .B(n32724), .Z(n32726) );
  XNOR U9404 ( .A(n32727), .B(n32301), .Z(n32303) );
  XNOR U9405 ( .A(n32304), .B(n31872), .Z(n31874) );
  XNOR U9406 ( .A(n31875), .B(n31437), .Z(n31439) );
  XNOR U9407 ( .A(n31440), .B(n30996), .Z(n30998) );
  XNOR U9408 ( .A(n30999), .B(n30549), .Z(n30551) );
  XNOR U9409 ( .A(n30552), .B(n30096), .Z(n30098) );
  XNOR U9410 ( .A(n30099), .B(n29637), .Z(n29639) );
  XNOR U9411 ( .A(n29640), .B(n29172), .Z(n29174) );
  XNOR U9412 ( .A(n29175), .B(n28701), .Z(n28703) );
  XNOR U9413 ( .A(n28704), .B(n28224), .Z(n28226) );
  XNOR U9414 ( .A(n28227), .B(n27741), .Z(n27743) );
  XNOR U9415 ( .A(n27744), .B(n27252), .Z(n27254) );
  XNOR U9416 ( .A(n27255), .B(n26755), .Z(n26757) );
  XNOR U9417 ( .A(n26758), .B(n26254), .Z(n26256) );
  XNOR U9418 ( .A(n26257), .B(n25746), .Z(n25748) );
  XNOR U9419 ( .A(n25749), .B(n25232), .Z(n25234) );
  XNOR U9420 ( .A(n25235), .B(n24709), .Z(n24711) );
  XNOR U9421 ( .A(n24712), .B(n24184), .Z(n24186) );
  XNOR U9422 ( .A(n24187), .B(n23653), .Z(n23655) );
  XNOR U9423 ( .A(n23656), .B(n23115), .Z(n23117) );
  XNOR U9424 ( .A(n23118), .B(n22571), .Z(n22573) );
  XNOR U9425 ( .A(n22574), .B(n22022), .Z(n22024) );
  XNOR U9426 ( .A(n22025), .B(n21467), .Z(n21469) );
  XNOR U9427 ( .A(n21470), .B(n20905), .Z(n20907) );
  XNOR U9428 ( .A(n20908), .B(n20338), .Z(n20340) );
  XNOR U9429 ( .A(n20341), .B(n19765), .Z(n19767) );
  XNOR U9430 ( .A(n19768), .B(n19186), .Z(n19188) );
  XOR U9431 ( .A(n17902), .B(n18007), .Z(n17906) );
  XOR U9432 ( .A(n16700), .B(n16805), .Z(n16704) );
  XOR U9433 ( .A(n15474), .B(n15579), .Z(n15478) );
  XOR U9434 ( .A(n14224), .B(n14329), .Z(n14228) );
  XOR U9435 ( .A(n9658), .B(n9763), .Z(n9662) );
  XOR U9436 ( .A(n8300), .B(n8405), .Z(n8304) );
  XOR U9437 ( .A(n6188), .B(n6329), .Z(n6192) );
  XOR U9438 ( .A(n4748), .B(n4913), .Z(n4752) );
  XOR U9439 ( .A(n4703), .B(n4922), .Z(n4707) );
  XOR U9440 ( .A(n3291), .B(n3474), .Z(n3295) );
  XOR U9441 ( .A(n3246), .B(n3483), .Z(n3250) );
  XOR U9442 ( .A(n1760), .B(n2021), .Z(n1764) );
  XOR U9443 ( .A(n1715), .B(n2030), .Z(n1719) );
  XOR U9444 ( .A(n4733), .B(n4916), .Z(n4737) );
  XOR U9445 ( .A(n6218), .B(n6323), .Z(n6222) );
  XOR U9446 ( .A(n4778), .B(n4907), .Z(n4782) );
  XNOR U9447 ( .A(n46237), .B(n46111), .Z(n46113) );
  XOR U9448 ( .A(n13600), .B(n13693), .Z(n13604) );
  XOR U9449 ( .A(n12312), .B(n12407), .Z(n12316) );
  XOR U9450 ( .A(n1745), .B(n2024), .Z(n1749) );
  XOR U9451 ( .A(n3276), .B(n3477), .Z(n3280) );
  XOR U9452 ( .A(n1790), .B(n2015), .Z(n1794) );
  XOR U9453 ( .A(n3321), .B(n3468), .Z(n3325) );
  XNOR U9454 ( .A(n46854), .B(n46764), .Z(n46766) );
  XNOR U9455 ( .A(n46767), .B(n46671), .Z(n46673) );
  XNOR U9456 ( .A(n46674), .B(n46572), .Z(n46574) );
  XNOR U9457 ( .A(n46575), .B(n46467), .Z(n46469) );
  XNOR U9458 ( .A(n46470), .B(n46356), .Z(n46358) );
  XNOR U9459 ( .A(n46242), .B(n46116), .Z(n46118) );
  XNOR U9460 ( .A(n46119), .B(n45987), .Z(n45989) );
  XNOR U9461 ( .A(n45990), .B(n45852), .Z(n45854) );
  XNOR U9462 ( .A(n45855), .B(n45711), .Z(n45713) );
  XNOR U9463 ( .A(n45714), .B(n45564), .Z(n45566) );
  XNOR U9464 ( .A(n45567), .B(n45411), .Z(n45413) );
  XNOR U9465 ( .A(n45414), .B(n45252), .Z(n45254) );
  XNOR U9466 ( .A(n45255), .B(n45087), .Z(n45089) );
  XNOR U9467 ( .A(n45090), .B(n44916), .Z(n44918) );
  XNOR U9468 ( .A(n44919), .B(n44739), .Z(n44741) );
  XNOR U9469 ( .A(n44742), .B(n44556), .Z(n44558) );
  XNOR U9470 ( .A(n44559), .B(n44367), .Z(n44369) );
  XNOR U9471 ( .A(n44370), .B(n44172), .Z(n44174) );
  XNOR U9472 ( .A(n44175), .B(n43971), .Z(n43973) );
  XNOR U9473 ( .A(n43974), .B(n43764), .Z(n43766) );
  XNOR U9474 ( .A(n43767), .B(n43551), .Z(n43553) );
  XNOR U9475 ( .A(n43554), .B(n43332), .Z(n43334) );
  XNOR U9476 ( .A(n43335), .B(n43107), .Z(n43109) );
  XNOR U9477 ( .A(n43110), .B(n42876), .Z(n42878) );
  XNOR U9478 ( .A(n42879), .B(n42639), .Z(n42641) );
  XNOR U9479 ( .A(n42642), .B(n42396), .Z(n42398) );
  XNOR U9480 ( .A(n42399), .B(n42147), .Z(n42149) );
  XNOR U9481 ( .A(n42150), .B(n41892), .Z(n41894) );
  XNOR U9482 ( .A(n41895), .B(n41631), .Z(n41633) );
  XNOR U9483 ( .A(n41634), .B(n41364), .Z(n41366) );
  XNOR U9484 ( .A(n41367), .B(n41091), .Z(n41093) );
  XNOR U9485 ( .A(n41094), .B(n40812), .Z(n40814) );
  XNOR U9486 ( .A(n40815), .B(n40527), .Z(n40529) );
  XNOR U9487 ( .A(n40530), .B(n40236), .Z(n40238) );
  XNOR U9488 ( .A(n40239), .B(n39939), .Z(n39941) );
  XNOR U9489 ( .A(n39942), .B(n39636), .Z(n39638) );
  XNOR U9490 ( .A(n39639), .B(n39327), .Z(n39329) );
  XNOR U9491 ( .A(n39330), .B(n39012), .Z(n39014) );
  XNOR U9492 ( .A(n39015), .B(n38691), .Z(n38693) );
  XNOR U9493 ( .A(n38694), .B(n38364), .Z(n38366) );
  XNOR U9494 ( .A(n38367), .B(n38031), .Z(n38033) );
  XNOR U9495 ( .A(n38034), .B(n37692), .Z(n37694) );
  XNOR U9496 ( .A(n37695), .B(n37347), .Z(n37349) );
  XNOR U9497 ( .A(n37350), .B(n36996), .Z(n36998) );
  XNOR U9498 ( .A(n36999), .B(n36639), .Z(n36641) );
  XNOR U9499 ( .A(n36642), .B(n36276), .Z(n36278) );
  XNOR U9500 ( .A(n36279), .B(n35907), .Z(n35909) );
  XNOR U9501 ( .A(n35910), .B(n35532), .Z(n35534) );
  XNOR U9502 ( .A(n35535), .B(n35151), .Z(n35153) );
  XNOR U9503 ( .A(n35154), .B(n34764), .Z(n34766) );
  XNOR U9504 ( .A(n34767), .B(n34371), .Z(n34373) );
  XNOR U9505 ( .A(n34374), .B(n33972), .Z(n33974) );
  XNOR U9506 ( .A(n33975), .B(n33567), .Z(n33569) );
  XNOR U9507 ( .A(n33570), .B(n33156), .Z(n33158) );
  XNOR U9508 ( .A(n33159), .B(n32739), .Z(n32741) );
  XNOR U9509 ( .A(n32742), .B(n32316), .Z(n32318) );
  XNOR U9510 ( .A(n32319), .B(n31887), .Z(n31889) );
  XNOR U9511 ( .A(n31890), .B(n31452), .Z(n31454) );
  XNOR U9512 ( .A(n31455), .B(n31011), .Z(n31013) );
  XNOR U9513 ( .A(n31014), .B(n30564), .Z(n30566) );
  XNOR U9514 ( .A(n30567), .B(n30111), .Z(n30113) );
  XNOR U9515 ( .A(n30114), .B(n29652), .Z(n29654) );
  XNOR U9516 ( .A(n29655), .B(n29187), .Z(n29189) );
  XNOR U9517 ( .A(n29190), .B(n28716), .Z(n28718) );
  XNOR U9518 ( .A(n28719), .B(n28239), .Z(n28241) );
  XNOR U9519 ( .A(n28242), .B(n27756), .Z(n27758) );
  XNOR U9520 ( .A(n27759), .B(n27267), .Z(n27269) );
  XNOR U9521 ( .A(n27270), .B(n26770), .Z(n26772) );
  XNOR U9522 ( .A(n26773), .B(n26269), .Z(n26271) );
  XNOR U9523 ( .A(n26272), .B(n25761), .Z(n25763) );
  XNOR U9524 ( .A(n25764), .B(n25247), .Z(n25249) );
  XNOR U9525 ( .A(n25250), .B(n24724), .Z(n24726) );
  XNOR U9526 ( .A(n24727), .B(n24199), .Z(n24201) );
  XNOR U9527 ( .A(n24202), .B(n23668), .Z(n23670) );
  XNOR U9528 ( .A(n23671), .B(n23130), .Z(n23132) );
  XNOR U9529 ( .A(n23133), .B(n22586), .Z(n22588) );
  XNOR U9530 ( .A(n22589), .B(n22037), .Z(n22039) );
  XNOR U9531 ( .A(n22040), .B(n21482), .Z(n21484) );
  XNOR U9532 ( .A(n21485), .B(n20920), .Z(n20922) );
  XNOR U9533 ( .A(n20923), .B(n20353), .Z(n20355) );
  XNOR U9534 ( .A(n20356), .B(n19780), .Z(n19782) );
  XNOR U9535 ( .A(n19783), .B(n19201), .Z(n19203) );
  XOR U9536 ( .A(n18509), .B(n18615), .Z(n18513) );
  XOR U9537 ( .A(n17319), .B(n17406), .Z(n17323) );
  XOR U9538 ( .A(n16105), .B(n16192), .Z(n16109) );
  XOR U9539 ( .A(n14867), .B(n14954), .Z(n14871) );
  XOR U9540 ( .A(n11665), .B(n11752), .Z(n11669) );
  XOR U9541 ( .A(n10343), .B(n10430), .Z(n10347) );
  XOR U9542 ( .A(n8997), .B(n9084), .Z(n9001) );
  XOR U9543 ( .A(n7627), .B(n7714), .Z(n7631) );
  XOR U9544 ( .A(n6233), .B(n6320), .Z(n6237) );
  XOR U9545 ( .A(n4808), .B(n4901), .Z(n4812) );
  XOR U9546 ( .A(n4763), .B(n4910), .Z(n4767) );
  XOR U9547 ( .A(n3351), .B(n3462), .Z(n3355) );
  XOR U9548 ( .A(n3306), .B(n3471), .Z(n3310) );
  XOR U9549 ( .A(n1820), .B(n2009), .Z(n1824) );
  XOR U9550 ( .A(n1775), .B(n2018), .Z(n1779) );
  XOR U9551 ( .A(n4793), .B(n4904), .Z(n4797) );
  XNOR U9552 ( .A(n46585), .B(n46477), .Z(n46479) );
  XOR U9553 ( .A(n14249), .B(n14324), .Z(n14253) );
  XOR U9554 ( .A(n1805), .B(n2012), .Z(n1809) );
  XOR U9555 ( .A(n3336), .B(n3465), .Z(n3340) );
  XOR U9556 ( .A(n1850), .B(n2003), .Z(n1854) );
  XNOR U9557 ( .A(n47094), .B(n47022), .Z(n47024) );
  XNOR U9558 ( .A(n47025), .B(n46947), .Z(n46949) );
  XNOR U9559 ( .A(n46950), .B(n46866), .Z(n46868) );
  XNOR U9560 ( .A(n46869), .B(n46779), .Z(n46781) );
  XNOR U9561 ( .A(n46782), .B(n46686), .Z(n46688) );
  XNOR U9562 ( .A(n46590), .B(n46482), .Z(n46484) );
  XNOR U9563 ( .A(n46485), .B(n46371), .Z(n46373) );
  XNOR U9564 ( .A(n46374), .B(n46254), .Z(n46256) );
  XNOR U9565 ( .A(n46257), .B(n46131), .Z(n46133) );
  XNOR U9566 ( .A(n46134), .B(n46002), .Z(n46004) );
  XNOR U9567 ( .A(n46005), .B(n45867), .Z(n45869) );
  XNOR U9568 ( .A(n45870), .B(n45726), .Z(n45728) );
  XNOR U9569 ( .A(n45729), .B(n45579), .Z(n45581) );
  XNOR U9570 ( .A(n45582), .B(n45426), .Z(n45428) );
  XNOR U9571 ( .A(n45429), .B(n45267), .Z(n45269) );
  XNOR U9572 ( .A(n45270), .B(n45102), .Z(n45104) );
  XNOR U9573 ( .A(n45105), .B(n44931), .Z(n44933) );
  XNOR U9574 ( .A(n44934), .B(n44754), .Z(n44756) );
  XNOR U9575 ( .A(n44757), .B(n44571), .Z(n44573) );
  XNOR U9576 ( .A(n44574), .B(n44382), .Z(n44384) );
  XNOR U9577 ( .A(n44385), .B(n44187), .Z(n44189) );
  XNOR U9578 ( .A(n44190), .B(n43986), .Z(n43988) );
  XNOR U9579 ( .A(n43989), .B(n43779), .Z(n43781) );
  XNOR U9580 ( .A(n43782), .B(n43566), .Z(n43568) );
  XNOR U9581 ( .A(n43569), .B(n43347), .Z(n43349) );
  XNOR U9582 ( .A(n43350), .B(n43122), .Z(n43124) );
  XNOR U9583 ( .A(n43125), .B(n42891), .Z(n42893) );
  XNOR U9584 ( .A(n42894), .B(n42654), .Z(n42656) );
  XNOR U9585 ( .A(n42657), .B(n42411), .Z(n42413) );
  XNOR U9586 ( .A(n42414), .B(n42162), .Z(n42164) );
  XNOR U9587 ( .A(n42165), .B(n41907), .Z(n41909) );
  XNOR U9588 ( .A(n41910), .B(n41646), .Z(n41648) );
  XNOR U9589 ( .A(n41649), .B(n41379), .Z(n41381) );
  XNOR U9590 ( .A(n41382), .B(n41106), .Z(n41108) );
  XNOR U9591 ( .A(n41109), .B(n40827), .Z(n40829) );
  XNOR U9592 ( .A(n40830), .B(n40542), .Z(n40544) );
  XNOR U9593 ( .A(n40545), .B(n40251), .Z(n40253) );
  XNOR U9594 ( .A(n40254), .B(n39954), .Z(n39956) );
  XNOR U9595 ( .A(n39957), .B(n39651), .Z(n39653) );
  XNOR U9596 ( .A(n39654), .B(n39342), .Z(n39344) );
  XNOR U9597 ( .A(n39345), .B(n39027), .Z(n39029) );
  XNOR U9598 ( .A(n39030), .B(n38706), .Z(n38708) );
  XNOR U9599 ( .A(n38709), .B(n38379), .Z(n38381) );
  XNOR U9600 ( .A(n38382), .B(n38046), .Z(n38048) );
  XNOR U9601 ( .A(n38049), .B(n37707), .Z(n37709) );
  XNOR U9602 ( .A(n37710), .B(n37362), .Z(n37364) );
  XNOR U9603 ( .A(n37365), .B(n37011), .Z(n37013) );
  XNOR U9604 ( .A(n37014), .B(n36654), .Z(n36656) );
  XNOR U9605 ( .A(n36657), .B(n36291), .Z(n36293) );
  XNOR U9606 ( .A(n36294), .B(n35922), .Z(n35924) );
  XNOR U9607 ( .A(n35925), .B(n35547), .Z(n35549) );
  XNOR U9608 ( .A(n35550), .B(n35166), .Z(n35168) );
  XNOR U9609 ( .A(n35169), .B(n34779), .Z(n34781) );
  XNOR U9610 ( .A(n34782), .B(n34386), .Z(n34388) );
  XNOR U9611 ( .A(n34389), .B(n33987), .Z(n33989) );
  XNOR U9612 ( .A(n33990), .B(n33582), .Z(n33584) );
  XNOR U9613 ( .A(n33585), .B(n33171), .Z(n33173) );
  XNOR U9614 ( .A(n33174), .B(n32754), .Z(n32756) );
  XNOR U9615 ( .A(n32757), .B(n32331), .Z(n32333) );
  XNOR U9616 ( .A(n32334), .B(n31902), .Z(n31904) );
  XNOR U9617 ( .A(n31905), .B(n31467), .Z(n31469) );
  XNOR U9618 ( .A(n31470), .B(n31026), .Z(n31028) );
  XNOR U9619 ( .A(n31029), .B(n30579), .Z(n30581) );
  XNOR U9620 ( .A(n30582), .B(n30126), .Z(n30128) );
  XNOR U9621 ( .A(n30129), .B(n29667), .Z(n29669) );
  XNOR U9622 ( .A(n29670), .B(n29202), .Z(n29204) );
  XNOR U9623 ( .A(n29205), .B(n28731), .Z(n28733) );
  XNOR U9624 ( .A(n28734), .B(n28254), .Z(n28256) );
  XNOR U9625 ( .A(n28257), .B(n27771), .Z(n27773) );
  XNOR U9626 ( .A(n27774), .B(n27282), .Z(n27284) );
  XNOR U9627 ( .A(n27285), .B(n26785), .Z(n26787) );
  XNOR U9628 ( .A(n26788), .B(n26284), .Z(n26286) );
  XNOR U9629 ( .A(n26287), .B(n25776), .Z(n25778) );
  XNOR U9630 ( .A(n25779), .B(n25262), .Z(n25264) );
  XNOR U9631 ( .A(n25265), .B(n24739), .Z(n24741) );
  XNOR U9632 ( .A(n24742), .B(n24214), .Z(n24216) );
  XNOR U9633 ( .A(n24217), .B(n23683), .Z(n23685) );
  XNOR U9634 ( .A(n23686), .B(n23145), .Z(n23147) );
  XNOR U9635 ( .A(n23148), .B(n22601), .Z(n22603) );
  XNOR U9636 ( .A(n22604), .B(n22052), .Z(n22054) );
  XNOR U9637 ( .A(n22055), .B(n21497), .Z(n21499) );
  XNOR U9638 ( .A(n21500), .B(n20935), .Z(n20937) );
  XNOR U9639 ( .A(n20938), .B(n20368), .Z(n20370) );
  XNOR U9640 ( .A(n20371), .B(n19795), .Z(n19797) );
  XNOR U9641 ( .A(n19798), .B(n19216), .Z(n19218) );
  XOR U9642 ( .A(n18524), .B(n18609), .Z(n18528) );
  XOR U9643 ( .A(n17334), .B(n17403), .Z(n17338) );
  XOR U9644 ( .A(n16120), .B(n16189), .Z(n16124) );
  XOR U9645 ( .A(n13620), .B(n13689), .Z(n13624) );
  XOR U9646 ( .A(n12332), .B(n12403), .Z(n12336) );
  XOR U9647 ( .A(n11022), .B(n11091), .Z(n11026) );
  XOR U9648 ( .A(n9688), .B(n9757), .Z(n9692) );
  XOR U9649 ( .A(n8330), .B(n8399), .Z(n8334) );
  XOR U9650 ( .A(n6948), .B(n7017), .Z(n6952) );
  XOR U9651 ( .A(n4823), .B(n4898), .Z(n4827) );
  XOR U9652 ( .A(n2646), .B(n2727), .Z(n2650) );
  XOR U9653 ( .A(n3366), .B(n3459), .Z(n3370) );
  XOR U9654 ( .A(n1880), .B(n1997), .Z(n1884) );
  XOR U9655 ( .A(n1835), .B(n2006), .Z(n1839) );
  XNOR U9656 ( .A(n46879), .B(n46789), .Z(n46791) );
  XOR U9657 ( .A(n15514), .B(n15571), .Z(n15518) );
  XOR U9658 ( .A(n1865), .B(n2000), .Z(n1869) );
  XNOR U9659 ( .A(n47279), .B(n47225), .Z(n47227) );
  XNOR U9660 ( .A(n47228), .B(n47169), .Z(n47171) );
  XNOR U9661 ( .A(n47172), .B(n47106), .Z(n47108) );
  XNOR U9662 ( .A(n47109), .B(n47037), .Z(n47039) );
  XNOR U9663 ( .A(n47040), .B(n46962), .Z(n46964) );
  XNOR U9664 ( .A(n46884), .B(n46794), .Z(n46796) );
  XNOR U9665 ( .A(n46797), .B(n46701), .Z(n46703) );
  XNOR U9666 ( .A(n46704), .B(n46602), .Z(n46604) );
  XNOR U9667 ( .A(n46605), .B(n46497), .Z(n46499) );
  XNOR U9668 ( .A(n46500), .B(n46386), .Z(n46388) );
  XNOR U9669 ( .A(n46389), .B(n46269), .Z(n46271) );
  XNOR U9670 ( .A(n46272), .B(n46146), .Z(n46148) );
  XNOR U9671 ( .A(n46149), .B(n46017), .Z(n46019) );
  XNOR U9672 ( .A(n46020), .B(n45882), .Z(n45884) );
  XNOR U9673 ( .A(n45885), .B(n45741), .Z(n45743) );
  XNOR U9674 ( .A(n45744), .B(n45594), .Z(n45596) );
  XNOR U9675 ( .A(n45597), .B(n45441), .Z(n45443) );
  XNOR U9676 ( .A(n45444), .B(n45282), .Z(n45284) );
  XNOR U9677 ( .A(n45285), .B(n45117), .Z(n45119) );
  XNOR U9678 ( .A(n45120), .B(n44946), .Z(n44948) );
  XNOR U9679 ( .A(n44949), .B(n44769), .Z(n44771) );
  XNOR U9680 ( .A(n44772), .B(n44586), .Z(n44588) );
  XNOR U9681 ( .A(n44589), .B(n44397), .Z(n44399) );
  XNOR U9682 ( .A(n44400), .B(n44202), .Z(n44204) );
  XNOR U9683 ( .A(n44205), .B(n44001), .Z(n44003) );
  XNOR U9684 ( .A(n44004), .B(n43794), .Z(n43796) );
  XNOR U9685 ( .A(n43797), .B(n43581), .Z(n43583) );
  XNOR U9686 ( .A(n43584), .B(n43362), .Z(n43364) );
  XNOR U9687 ( .A(n43365), .B(n43137), .Z(n43139) );
  XNOR U9688 ( .A(n43140), .B(n42906), .Z(n42908) );
  XNOR U9689 ( .A(n42909), .B(n42669), .Z(n42671) );
  XNOR U9690 ( .A(n42672), .B(n42426), .Z(n42428) );
  XNOR U9691 ( .A(n42429), .B(n42177), .Z(n42179) );
  XNOR U9692 ( .A(n42180), .B(n41922), .Z(n41924) );
  XNOR U9693 ( .A(n41925), .B(n41661), .Z(n41663) );
  XNOR U9694 ( .A(n41664), .B(n41394), .Z(n41396) );
  XNOR U9695 ( .A(n41397), .B(n41121), .Z(n41123) );
  XNOR U9696 ( .A(n41124), .B(n40842), .Z(n40844) );
  XNOR U9697 ( .A(n40845), .B(n40557), .Z(n40559) );
  XNOR U9698 ( .A(n40560), .B(n40266), .Z(n40268) );
  XNOR U9699 ( .A(n40269), .B(n39969), .Z(n39971) );
  XNOR U9700 ( .A(n39972), .B(n39666), .Z(n39668) );
  XNOR U9701 ( .A(n39669), .B(n39357), .Z(n39359) );
  XNOR U9702 ( .A(n39360), .B(n39042), .Z(n39044) );
  XNOR U9703 ( .A(n39045), .B(n38721), .Z(n38723) );
  XNOR U9704 ( .A(n38724), .B(n38394), .Z(n38396) );
  XNOR U9705 ( .A(n38397), .B(n38061), .Z(n38063) );
  XNOR U9706 ( .A(n38064), .B(n37722), .Z(n37724) );
  XNOR U9707 ( .A(n37725), .B(n37377), .Z(n37379) );
  XNOR U9708 ( .A(n37380), .B(n37026), .Z(n37028) );
  XNOR U9709 ( .A(n37029), .B(n36669), .Z(n36671) );
  XNOR U9710 ( .A(n36672), .B(n36306), .Z(n36308) );
  XNOR U9711 ( .A(n36309), .B(n35937), .Z(n35939) );
  XNOR U9712 ( .A(n35940), .B(n35562), .Z(n35564) );
  XNOR U9713 ( .A(n35565), .B(n35181), .Z(n35183) );
  XNOR U9714 ( .A(n35184), .B(n34794), .Z(n34796) );
  XNOR U9715 ( .A(n34797), .B(n34401), .Z(n34403) );
  XNOR U9716 ( .A(n34404), .B(n34002), .Z(n34004) );
  XNOR U9717 ( .A(n34005), .B(n33597), .Z(n33599) );
  XNOR U9718 ( .A(n33600), .B(n33186), .Z(n33188) );
  XNOR U9719 ( .A(n33189), .B(n32769), .Z(n32771) );
  XNOR U9720 ( .A(n32772), .B(n32346), .Z(n32348) );
  XNOR U9721 ( .A(n32349), .B(n31917), .Z(n31919) );
  XNOR U9722 ( .A(n31920), .B(n31482), .Z(n31484) );
  XNOR U9723 ( .A(n31485), .B(n31041), .Z(n31043) );
  XNOR U9724 ( .A(n31044), .B(n30594), .Z(n30596) );
  XNOR U9725 ( .A(n30597), .B(n30141), .Z(n30143) );
  XNOR U9726 ( .A(n30144), .B(n29682), .Z(n29684) );
  XNOR U9727 ( .A(n29685), .B(n29217), .Z(n29219) );
  XNOR U9728 ( .A(n29220), .B(n28746), .Z(n28748) );
  XNOR U9729 ( .A(n28749), .B(n28269), .Z(n28271) );
  XNOR U9730 ( .A(n28272), .B(n27786), .Z(n27788) );
  XNOR U9731 ( .A(n27789), .B(n27297), .Z(n27299) );
  XNOR U9732 ( .A(n27300), .B(n26800), .Z(n26802) );
  XNOR U9733 ( .A(n26803), .B(n26299), .Z(n26301) );
  XNOR U9734 ( .A(n26302), .B(n25791), .Z(n25793) );
  XNOR U9735 ( .A(n25794), .B(n25277), .Z(n25279) );
  XNOR U9736 ( .A(n25280), .B(n24754), .Z(n24756) );
  XNOR U9737 ( .A(n24757), .B(n24229), .Z(n24231) );
  XNOR U9738 ( .A(n24232), .B(n23698), .Z(n23700) );
  XNOR U9739 ( .A(n23701), .B(n23160), .Z(n23162) );
  XNOR U9740 ( .A(n23163), .B(n22616), .Z(n22618) );
  XNOR U9741 ( .A(n22619), .B(n22067), .Z(n22069) );
  XNOR U9742 ( .A(n22070), .B(n21512), .Z(n21514) );
  XNOR U9743 ( .A(n21515), .B(n20950), .Z(n20952) );
  XNOR U9744 ( .A(n20953), .B(n20383), .Z(n20385) );
  XNOR U9745 ( .A(n20386), .B(n19810), .Z(n19812) );
  XNOR U9746 ( .A(n19813), .B(n19231), .Z(n19233) );
  XOR U9747 ( .A(n18539), .B(n18603), .Z(n18543) );
  XOR U9748 ( .A(n17349), .B(n17400), .Z(n17353) );
  XOR U9749 ( .A(n14897), .B(n14948), .Z(n14901) );
  XOR U9750 ( .A(n13635), .B(n13686), .Z(n13639) );
  XOR U9751 ( .A(n12347), .B(n12400), .Z(n12351) );
  XOR U9752 ( .A(n11037), .B(n11088), .Z(n11041) );
  XOR U9753 ( .A(n9703), .B(n9754), .Z(n9707) );
  XOR U9754 ( .A(n8345), .B(n8396), .Z(n8349) );
  XOR U9755 ( .A(n6963), .B(n7014), .Z(n6967) );
  XOR U9756 ( .A(n5555), .B(n5608), .Z(n5559) );
  XOR U9757 ( .A(n4125), .B(n4176), .Z(n4129) );
  XOR U9758 ( .A(n2671), .B(n2722), .Z(n2675) );
  XOR U9759 ( .A(n1915), .B(n1990), .Z(n1919) );
  XOR U9760 ( .A(n1895), .B(n1994), .Z(n1899) );
  XNOR U9761 ( .A(n47119), .B(n47047), .Z(n47049) );
  XOR U9762 ( .A(n16755), .B(n16794), .Z(n16759) );
  XNOR U9763 ( .A(n47411), .B(n47375), .Z(n47377) );
  XNOR U9764 ( .A(n47378), .B(n47336), .Z(n47338) );
  XNOR U9765 ( .A(n47339), .B(n47291), .Z(n47293) );
  XNOR U9766 ( .A(n47294), .B(n47240), .Z(n47242) );
  XNOR U9767 ( .A(n47243), .B(n47184), .Z(n47186) );
  XNOR U9768 ( .A(n47124), .B(n47052), .Z(n47054) );
  XNOR U9769 ( .A(n47055), .B(n46977), .Z(n46979) );
  XNOR U9770 ( .A(n46980), .B(n46896), .Z(n46898) );
  XNOR U9771 ( .A(n46899), .B(n46809), .Z(n46811) );
  XNOR U9772 ( .A(n46812), .B(n46716), .Z(n46718) );
  XNOR U9773 ( .A(n46719), .B(n46617), .Z(n46619) );
  XNOR U9774 ( .A(n46620), .B(n46512), .Z(n46514) );
  XNOR U9775 ( .A(n46515), .B(n46401), .Z(n46403) );
  XNOR U9776 ( .A(n46404), .B(n46284), .Z(n46286) );
  XNOR U9777 ( .A(n46287), .B(n46161), .Z(n46163) );
  XNOR U9778 ( .A(n46164), .B(n46032), .Z(n46034) );
  XNOR U9779 ( .A(n46035), .B(n45897), .Z(n45899) );
  XNOR U9780 ( .A(n45900), .B(n45756), .Z(n45758) );
  XNOR U9781 ( .A(n45759), .B(n45609), .Z(n45611) );
  XNOR U9782 ( .A(n45612), .B(n45456), .Z(n45458) );
  XNOR U9783 ( .A(n45459), .B(n45297), .Z(n45299) );
  XNOR U9784 ( .A(n45300), .B(n45132), .Z(n45134) );
  XNOR U9785 ( .A(n45135), .B(n44961), .Z(n44963) );
  XNOR U9786 ( .A(n44964), .B(n44784), .Z(n44786) );
  XNOR U9787 ( .A(n44787), .B(n44601), .Z(n44603) );
  XNOR U9788 ( .A(n44604), .B(n44412), .Z(n44414) );
  XNOR U9789 ( .A(n44415), .B(n44217), .Z(n44219) );
  XNOR U9790 ( .A(n44220), .B(n44016), .Z(n44018) );
  XNOR U9791 ( .A(n44019), .B(n43809), .Z(n43811) );
  XNOR U9792 ( .A(n43812), .B(n43596), .Z(n43598) );
  XNOR U9793 ( .A(n43599), .B(n43377), .Z(n43379) );
  XNOR U9794 ( .A(n43380), .B(n43152), .Z(n43154) );
  XNOR U9795 ( .A(n43155), .B(n42921), .Z(n42923) );
  XNOR U9796 ( .A(n42924), .B(n42684), .Z(n42686) );
  XNOR U9797 ( .A(n42687), .B(n42441), .Z(n42443) );
  XNOR U9798 ( .A(n42444), .B(n42192), .Z(n42194) );
  XNOR U9799 ( .A(n42195), .B(n41937), .Z(n41939) );
  XNOR U9800 ( .A(n41940), .B(n41676), .Z(n41678) );
  XNOR U9801 ( .A(n41679), .B(n41409), .Z(n41411) );
  XNOR U9802 ( .A(n41412), .B(n41136), .Z(n41138) );
  XNOR U9803 ( .A(n41139), .B(n40857), .Z(n40859) );
  XNOR U9804 ( .A(n40860), .B(n40572), .Z(n40574) );
  XNOR U9805 ( .A(n40575), .B(n40281), .Z(n40283) );
  XNOR U9806 ( .A(n40284), .B(n39984), .Z(n39986) );
  XNOR U9807 ( .A(n39987), .B(n39681), .Z(n39683) );
  XNOR U9808 ( .A(n39684), .B(n39372), .Z(n39374) );
  XNOR U9809 ( .A(n39375), .B(n39057), .Z(n39059) );
  XNOR U9810 ( .A(n39060), .B(n38736), .Z(n38738) );
  XNOR U9811 ( .A(n38739), .B(n38409), .Z(n38411) );
  XNOR U9812 ( .A(n38412), .B(n38076), .Z(n38078) );
  XNOR U9813 ( .A(n38079), .B(n37737), .Z(n37739) );
  XNOR U9814 ( .A(n37740), .B(n37392), .Z(n37394) );
  XNOR U9815 ( .A(n37395), .B(n37041), .Z(n37043) );
  XNOR U9816 ( .A(n37044), .B(n36684), .Z(n36686) );
  XNOR U9817 ( .A(n36687), .B(n36321), .Z(n36323) );
  XNOR U9818 ( .A(n36324), .B(n35952), .Z(n35954) );
  XNOR U9819 ( .A(n35955), .B(n35577), .Z(n35579) );
  XNOR U9820 ( .A(n35580), .B(n35196), .Z(n35198) );
  XNOR U9821 ( .A(n35199), .B(n34809), .Z(n34811) );
  XNOR U9822 ( .A(n34812), .B(n34416), .Z(n34418) );
  XNOR U9823 ( .A(n34419), .B(n34017), .Z(n34019) );
  XNOR U9824 ( .A(n34020), .B(n33612), .Z(n33614) );
  XNOR U9825 ( .A(n33615), .B(n33201), .Z(n33203) );
  XNOR U9826 ( .A(n33204), .B(n32784), .Z(n32786) );
  XNOR U9827 ( .A(n32787), .B(n32361), .Z(n32363) );
  XNOR U9828 ( .A(n32364), .B(n31932), .Z(n31934) );
  XNOR U9829 ( .A(n31935), .B(n31497), .Z(n31499) );
  XNOR U9830 ( .A(n31500), .B(n31056), .Z(n31058) );
  XNOR U9831 ( .A(n31059), .B(n30609), .Z(n30611) );
  XNOR U9832 ( .A(n30612), .B(n30156), .Z(n30158) );
  XNOR U9833 ( .A(n30159), .B(n29697), .Z(n29699) );
  XNOR U9834 ( .A(n29700), .B(n29232), .Z(n29234) );
  XNOR U9835 ( .A(n29235), .B(n28761), .Z(n28763) );
  XNOR U9836 ( .A(n28764), .B(n28284), .Z(n28286) );
  XNOR U9837 ( .A(n28287), .B(n27801), .Z(n27803) );
  XNOR U9838 ( .A(n27804), .B(n27312), .Z(n27314) );
  XNOR U9839 ( .A(n27315), .B(n26815), .Z(n26817) );
  XNOR U9840 ( .A(n26818), .B(n26314), .Z(n26316) );
  XNOR U9841 ( .A(n26317), .B(n25806), .Z(n25808) );
  XNOR U9842 ( .A(n25809), .B(n25292), .Z(n25294) );
  XNOR U9843 ( .A(n25295), .B(n24769), .Z(n24771) );
  XNOR U9844 ( .A(n24772), .B(n24244), .Z(n24246) );
  XNOR U9845 ( .A(n24247), .B(n23713), .Z(n23715) );
  XNOR U9846 ( .A(n23716), .B(n23175), .Z(n23177) );
  XNOR U9847 ( .A(n23178), .B(n22631), .Z(n22633) );
  XNOR U9848 ( .A(n22634), .B(n22082), .Z(n22084) );
  XNOR U9849 ( .A(n22085), .B(n21527), .Z(n21529) );
  XNOR U9850 ( .A(n21530), .B(n20965), .Z(n20967) );
  XNOR U9851 ( .A(n20968), .B(n20398), .Z(n20400) );
  XNOR U9852 ( .A(n20401), .B(n19825), .Z(n19827) );
  XNOR U9853 ( .A(n19828), .B(n19246), .Z(n19248) );
  XOR U9854 ( .A(n18554), .B(n18597), .Z(n18558) );
  XOR U9855 ( .A(n16150), .B(n16183), .Z(n16154) );
  XOR U9856 ( .A(n14912), .B(n14945), .Z(n14916) );
  XOR U9857 ( .A(n13650), .B(n13683), .Z(n13654) );
  XOR U9858 ( .A(n12362), .B(n12397), .Z(n12366) );
  XOR U9859 ( .A(n11052), .B(n11085), .Z(n11056) );
  XOR U9860 ( .A(n9718), .B(n9751), .Z(n9722) );
  XOR U9861 ( .A(n8360), .B(n8393), .Z(n8364) );
  XOR U9862 ( .A(n6978), .B(n7011), .Z(n6982) );
  XOR U9863 ( .A(n5570), .B(n5605), .Z(n5574) );
  XOR U9864 ( .A(n4140), .B(n4173), .Z(n4144) );
  XOR U9865 ( .A(n2686), .B(n2719), .Z(n2690) );
  XNOR U9866 ( .A(n47304), .B(n47250), .Z(n47252) );
  XOR U9867 ( .A(n17972), .B(n17993), .Z(n17976) );
  XOR U9868 ( .A(n47468), .B(n47473), .Z(n47457) );
  XNOR U9869 ( .A(n47451), .B(n47450), .Z(n47431) );
  XOR U9870 ( .A(n47420), .B(n47425), .Z(n47397) );
  XOR U9871 ( .A(n47387), .B(n47392), .Z(n47358) );
  XNOR U9872 ( .A(n47352), .B(n47351), .Z(n47314) );
  XNOR U9873 ( .A(n47200), .B(n47199), .Z(n47144) );
  XOR U9874 ( .A(n47133), .B(n47138), .Z(n47074) );
  XOR U9875 ( .A(n47064), .B(n47069), .Z(n46999) );
  XNOR U9876 ( .A(n46993), .B(n46992), .Z(n46919) );
  XOR U9877 ( .A(n46908), .B(n46913), .Z(n46831) );
  XOR U9878 ( .A(n46821), .B(n46826), .Z(n46738) );
  XNOR U9879 ( .A(n46732), .B(n46731), .Z(n46640) );
  XOR U9880 ( .A(n46629), .B(n46634), .Z(n46534) );
  XOR U9881 ( .A(n46524), .B(n46529), .Z(n46423) );
  XNOR U9882 ( .A(n46417), .B(n46416), .Z(n46307) );
  XOR U9883 ( .A(n46296), .B(n46301), .Z(n46183) );
  XOR U9884 ( .A(n46173), .B(n46178), .Z(n46054) );
  XNOR U9885 ( .A(n46048), .B(n46047), .Z(n45920) );
  XOR U9886 ( .A(n45909), .B(n45914), .Z(n45778) );
  XOR U9887 ( .A(n45768), .B(n45773), .Z(n45631) );
  XNOR U9888 ( .A(n45625), .B(n45624), .Z(n45479) );
  XOR U9889 ( .A(n45468), .B(n45473), .Z(n45319) );
  XOR U9890 ( .A(n45309), .B(n45314), .Z(n45154) );
  XNOR U9891 ( .A(n45148), .B(n45147), .Z(n44984) );
  XOR U9892 ( .A(n44973), .B(n44978), .Z(n44806) );
  XOR U9893 ( .A(n44796), .B(n44801), .Z(n44623) );
  XNOR U9894 ( .A(n44617), .B(n44616), .Z(n44435) );
  XOR U9895 ( .A(n44424), .B(n44429), .Z(n44239) );
  XOR U9896 ( .A(n44229), .B(n44234), .Z(n44038) );
  XNOR U9897 ( .A(n44032), .B(n44031), .Z(n43832) );
  XOR U9898 ( .A(n43821), .B(n43826), .Z(n43618) );
  XOR U9899 ( .A(n43608), .B(n43613), .Z(n43399) );
  XNOR U9900 ( .A(n43393), .B(n43392), .Z(n43175) );
  XOR U9901 ( .A(n43164), .B(n43169), .Z(n42943) );
  XOR U9902 ( .A(n42933), .B(n42938), .Z(n42706) );
  XNOR U9903 ( .A(n42700), .B(n42699), .Z(n42464) );
  XOR U9904 ( .A(n42453), .B(n42458), .Z(n42214) );
  XOR U9905 ( .A(n42204), .B(n42209), .Z(n41959) );
  XNOR U9906 ( .A(n41953), .B(n41952), .Z(n41699) );
  XOR U9907 ( .A(n41688), .B(n41693), .Z(n41431) );
  XOR U9908 ( .A(n41421), .B(n41426), .Z(n41158) );
  XNOR U9909 ( .A(n41152), .B(n41151), .Z(n40880) );
  XOR U9910 ( .A(n40869), .B(n40874), .Z(n40594) );
  XOR U9911 ( .A(n40584), .B(n40589), .Z(n40303) );
  XNOR U9912 ( .A(n40297), .B(n40296), .Z(n40007) );
  XOR U9913 ( .A(n39996), .B(n40001), .Z(n39703) );
  XOR U9914 ( .A(n39693), .B(n39698), .Z(n39394) );
  XNOR U9915 ( .A(n39388), .B(n39387), .Z(n39080) );
  XOR U9916 ( .A(n39069), .B(n39074), .Z(n38758) );
  XOR U9917 ( .A(n38748), .B(n38753), .Z(n38431) );
  XNOR U9918 ( .A(n38425), .B(n38424), .Z(n38099) );
  XOR U9919 ( .A(n38088), .B(n38093), .Z(n37759) );
  XOR U9920 ( .A(n37749), .B(n37754), .Z(n37414) );
  XNOR U9921 ( .A(n37408), .B(n37407), .Z(n37064) );
  XOR U9922 ( .A(n37053), .B(n37058), .Z(n36706) );
  XOR U9923 ( .A(n36696), .B(n36701), .Z(n36343) );
  XNOR U9924 ( .A(n36337), .B(n36336), .Z(n35975) );
  XOR U9925 ( .A(n35964), .B(n35969), .Z(n35599) );
  XOR U9926 ( .A(n35589), .B(n35594), .Z(n35218) );
  XNOR U9927 ( .A(n35212), .B(n35211), .Z(n34832) );
  XOR U9928 ( .A(n34821), .B(n34826), .Z(n34438) );
  XOR U9929 ( .A(n34428), .B(n34433), .Z(n34039) );
  XNOR U9930 ( .A(n34033), .B(n34032), .Z(n33635) );
  XOR U9931 ( .A(n33624), .B(n33629), .Z(n33223) );
  XOR U9932 ( .A(n33213), .B(n33218), .Z(n32806) );
  XNOR U9933 ( .A(n32800), .B(n32799), .Z(n32384) );
  XOR U9934 ( .A(n32373), .B(n32378), .Z(n31954) );
  XOR U9935 ( .A(n31944), .B(n31949), .Z(n31519) );
  XNOR U9936 ( .A(n31513), .B(n31512), .Z(n31079) );
  XOR U9937 ( .A(n31068), .B(n31073), .Z(n30631) );
  XOR U9938 ( .A(n30621), .B(n30626), .Z(n30178) );
  XNOR U9939 ( .A(n30172), .B(n30171), .Z(n29720) );
  XOR U9940 ( .A(n29709), .B(n29714), .Z(n29254) );
  XOR U9941 ( .A(n29244), .B(n29249), .Z(n28783) );
  XNOR U9942 ( .A(n28777), .B(n28776), .Z(n28307) );
  XOR U9943 ( .A(n28296), .B(n28301), .Z(n27823) );
  XOR U9944 ( .A(n27813), .B(n27818), .Z(n27334) );
  XNOR U9945 ( .A(n27328), .B(n27327), .Z(n26838) );
  XOR U9946 ( .A(n26827), .B(n26832), .Z(n26336) );
  XOR U9947 ( .A(n26326), .B(n26331), .Z(n25828) );
  XNOR U9948 ( .A(n25822), .B(n25821), .Z(n25315) );
  XOR U9949 ( .A(n25304), .B(n25309), .Z(n24791) );
  XOR U9950 ( .A(n24781), .B(n24786), .Z(n24266) );
  XNOR U9951 ( .A(n24260), .B(n24259), .Z(n23736) );
  XOR U9952 ( .A(n23725), .B(n23730), .Z(n23197) );
  XOR U9953 ( .A(n23187), .B(n23192), .Z(n22653) );
  XNOR U9954 ( .A(n22647), .B(n22646), .Z(n22105) );
  XOR U9955 ( .A(n22094), .B(n22099), .Z(n21549) );
  XOR U9956 ( .A(n21539), .B(n21544), .Z(n20987) );
  XNOR U9957 ( .A(n20981), .B(n20980), .Z(n20421) );
  XOR U9958 ( .A(n20410), .B(n20415), .Z(n19847) );
  XOR U9959 ( .A(n19837), .B(n19842), .Z(n19268) );
  XOR U9960 ( .A(n17379), .B(n17394), .Z(n17388) );
  XOR U9961 ( .A(n16165), .B(n16180), .Z(n16174) );
  XOR U9962 ( .A(n14927), .B(n14942), .Z(n14936) );
  XOR U9963 ( .A(n13665), .B(n13680), .Z(n13674) );
  XOR U9964 ( .A(n12377), .B(n12394), .Z(n12386) );
  XOR U9965 ( .A(n11067), .B(n11082), .Z(n11076) );
  XOR U9966 ( .A(n9733), .B(n9748), .Z(n9742) );
  XOR U9967 ( .A(n8375), .B(n8390), .Z(n8384) );
  XOR U9968 ( .A(n6993), .B(n7008), .Z(n7002) );
  XOR U9969 ( .A(n5585), .B(n5602), .Z(n5594) );
  XOR U9970 ( .A(n4155), .B(n4170), .Z(n4164) );
  XOR U9971 ( .A(n2701), .B(n2716), .Z(n2710) );
  XNOR U9972 ( .A(n47264), .B(n47261), .Z(n47209) );
  XNOR U9973 ( .A(n18589), .B(n18586), .Z(n18577) );
  XNOR U9974 ( .A(n27424), .B(n26932), .Z(n26934) );
  XNOR U9975 ( .A(n27429), .B(n26937), .Z(n26939) );
  XNOR U9976 ( .A(n27434), .B(n26942), .Z(n26944) );
  XNOR U9977 ( .A(n29804), .B(n29342), .Z(n29344) );
  XNOR U9978 ( .A(n29345), .B(n28877), .Z(n28879) );
  XNOR U9979 ( .A(n28880), .B(n28406), .Z(n28408) );
  XNOR U9980 ( .A(n27449), .B(n26957), .Z(n26959) );
  XNOR U9981 ( .A(n27439), .B(n26947), .Z(n26949) );
  XNOR U9982 ( .A(n25922), .B(n25411), .Z(n25413) );
  XNOR U9983 ( .A(n25947), .B(n25436), .Z(n25438) );
  XNOR U9984 ( .A(n27444), .B(n26952), .Z(n26954) );
  XNOR U9985 ( .A(n25927), .B(n25416), .Z(n25418) );
  XNOR U9986 ( .A(n25952), .B(n25441), .Z(n25443) );
  XNOR U9987 ( .A(n25932), .B(n25421), .Z(n25423) );
  XNOR U9988 ( .A(n31160), .B(n30716), .Z(n30718) );
  XNOR U9989 ( .A(n30719), .B(n30269), .Z(n30271) );
  XNOR U9990 ( .A(n30272), .B(n29816), .Z(n29818) );
  XNOR U9991 ( .A(n29819), .B(n29357), .Z(n29359) );
  XNOR U9992 ( .A(n29360), .B(n28892), .Z(n28894) );
  XNOR U9993 ( .A(n28895), .B(n28421), .Z(n28423) );
  XNOR U9994 ( .A(n28424), .B(n27944), .Z(n27946) );
  XNOR U9995 ( .A(n27947), .B(n27461), .Z(n27463) );
  XNOR U9996 ( .A(n27464), .B(n26972), .Z(n26974) );
  XNOR U9997 ( .A(n25977), .B(n25466), .Z(n25468) );
  XNOR U9998 ( .A(n25937), .B(n25426), .Z(n25428) );
  XNOR U9999 ( .A(n24362), .B(n23834), .Z(n23836) );
  XNOR U10000 ( .A(n25962), .B(n25451), .Z(n25453) );
  XNOR U10001 ( .A(n25444), .B(n24926), .Z(n24928) );
  XNOR U10002 ( .A(n24387), .B(n23859), .Z(n23861) );
  XNOR U10003 ( .A(n25942), .B(n25431), .Z(n25433) );
  XNOR U10004 ( .A(n24367), .B(n23839), .Z(n23841) );
  XNOR U10005 ( .A(n25967), .B(n25456), .Z(n25458) );
  XNOR U10006 ( .A(n24392), .B(n23864), .Z(n23866) );
  XNOR U10007 ( .A(n24372), .B(n23844), .Z(n23846) );
  XNOR U10008 ( .A(n24417), .B(n23889), .Z(n23891) );
  XNOR U10009 ( .A(n32462), .B(n32036), .Z(n32038) );
  XNOR U10010 ( .A(n32039), .B(n31607), .Z(n31609) );
  XNOR U10011 ( .A(n31610), .B(n31172), .Z(n31174) );
  XNOR U10012 ( .A(n31175), .B(n30731), .Z(n30733) );
  XNOR U10013 ( .A(n30734), .B(n30284), .Z(n30286) );
  XNOR U10014 ( .A(n30287), .B(n29831), .Z(n29833) );
  XNOR U10015 ( .A(n29834), .B(n29372), .Z(n29374) );
  XNOR U10016 ( .A(n29375), .B(n28907), .Z(n28909) );
  XNOR U10017 ( .A(n28910), .B(n28436), .Z(n28438) );
  XNOR U10018 ( .A(n28439), .B(n27959), .Z(n27961) );
  XNOR U10019 ( .A(n27962), .B(n27476), .Z(n27478) );
  XNOR U10020 ( .A(n27479), .B(n26987), .Z(n26989) );
  XNOR U10021 ( .A(n26990), .B(n26490), .Z(n26492) );
  XNOR U10022 ( .A(n26493), .B(n25989), .Z(n25991) );
  XNOR U10023 ( .A(n25992), .B(n25481), .Z(n25483) );
  XNOR U10024 ( .A(n24377), .B(n23849), .Z(n23851) );
  XNOR U10025 ( .A(n22753), .B(n22206), .Z(n22208) );
  XNOR U10026 ( .A(n24422), .B(n23894), .Z(n23896) );
  XNOR U10027 ( .A(n24447), .B(n23919), .Z(n23921) );
  XNOR U10028 ( .A(n25459), .B(n24941), .Z(n24943) );
  XNOR U10029 ( .A(n24402), .B(n23874), .Z(n23876) );
  XNOR U10030 ( .A(n23867), .B(n23333), .Z(n23335) );
  XNOR U10031 ( .A(n22778), .B(n22231), .Z(n22233) );
  XNOR U10032 ( .A(n24382), .B(n23854), .Z(n23856) );
  XNOR U10033 ( .A(n22758), .B(n22211), .Z(n22213) );
  XNOR U10034 ( .A(n24427), .B(n23899), .Z(n23901) );
  XNOR U10035 ( .A(n24407), .B(n23879), .Z(n23881) );
  XNOR U10036 ( .A(n22783), .B(n22236), .Z(n22238) );
  XNOR U10037 ( .A(n22763), .B(n22216), .Z(n22218) );
  XNOR U10038 ( .A(n24432), .B(n23904), .Z(n23906) );
  XNOR U10039 ( .A(n22808), .B(n22261), .Z(n22263) );
  XNOR U10040 ( .A(n33710), .B(n33302), .Z(n33304) );
  XNOR U10041 ( .A(n33305), .B(n32891), .Z(n32893) );
  XNOR U10042 ( .A(n32894), .B(n32474), .Z(n32476) );
  XNOR U10043 ( .A(n32477), .B(n32051), .Z(n32053) );
  XNOR U10044 ( .A(n32054), .B(n31622), .Z(n31624) );
  XNOR U10045 ( .A(n31625), .B(n31187), .Z(n31189) );
  XNOR U10046 ( .A(n31190), .B(n30746), .Z(n30748) );
  XNOR U10047 ( .A(n30749), .B(n30299), .Z(n30301) );
  XNOR U10048 ( .A(n30302), .B(n29846), .Z(n29848) );
  XNOR U10049 ( .A(n29849), .B(n29387), .Z(n29389) );
  XNOR U10050 ( .A(n29390), .B(n28922), .Z(n28924) );
  XNOR U10051 ( .A(n28925), .B(n28451), .Z(n28453) );
  XNOR U10052 ( .A(n28454), .B(n27974), .Z(n27976) );
  XNOR U10053 ( .A(n27977), .B(n27491), .Z(n27493) );
  XNOR U10054 ( .A(n27494), .B(n27002), .Z(n27004) );
  XNOR U10055 ( .A(n27005), .B(n26505), .Z(n26507) );
  XNOR U10056 ( .A(n26508), .B(n26004), .Z(n26006) );
  XNOR U10057 ( .A(n26007), .B(n25496), .Z(n25498) );
  XNOR U10058 ( .A(n25499), .B(n24981), .Z(n24983) );
  XNOR U10059 ( .A(n24457), .B(n23929), .Z(n23931) );
  XNOR U10060 ( .A(n23922), .B(n23388), .Z(n23390) );
  XNOR U10061 ( .A(n22768), .B(n22221), .Z(n22223) );
  XNOR U10062 ( .A(n21090), .B(n20525), .Z(n20527) );
  XNOR U10063 ( .A(n24437), .B(n23909), .Z(n23911) );
  XNOR U10064 ( .A(n22813), .B(n22266), .Z(n22268) );
  XNOR U10065 ( .A(n24462), .B(n23934), .Z(n23936) );
  XNOR U10066 ( .A(n22838), .B(n22291), .Z(n22293) );
  XNOR U10067 ( .A(n23882), .B(n23348), .Z(n23350) );
  XNOR U10068 ( .A(n22793), .B(n22246), .Z(n22248) );
  XNOR U10069 ( .A(n22239), .B(n21687), .Z(n21689) );
  XNOR U10070 ( .A(n21115), .B(n20550), .Z(n20552) );
  XNOR U10071 ( .A(n22773), .B(n22226), .Z(n22228) );
  XNOR U10072 ( .A(n21095), .B(n20530), .Z(n20532) );
  XNOR U10073 ( .A(n24442), .B(n23914), .Z(n23916) );
  XNOR U10074 ( .A(n22818), .B(n22271), .Z(n22273) );
  XNOR U10075 ( .A(n22798), .B(n22251), .Z(n22253) );
  XNOR U10076 ( .A(n21120), .B(n20555), .Z(n20557) );
  XNOR U10077 ( .A(n21100), .B(n20535), .Z(n20537) );
  XNOR U10078 ( .A(n22823), .B(n22276), .Z(n22278) );
  XNOR U10079 ( .A(n21145), .B(n20580), .Z(n20582) );
  XNOR U10080 ( .A(n22868), .B(n22321), .Z(n22323) );
  XNOR U10081 ( .A(n34904), .B(n34514), .Z(n34516) );
  XNOR U10082 ( .A(n34517), .B(n34121), .Z(n34123) );
  XNOR U10083 ( .A(n34124), .B(n33722), .Z(n33724) );
  XNOR U10084 ( .A(n33725), .B(n33317), .Z(n33319) );
  XNOR U10085 ( .A(n33320), .B(n32906), .Z(n32908) );
  XNOR U10086 ( .A(n32909), .B(n32489), .Z(n32491) );
  XNOR U10087 ( .A(n32492), .B(n32066), .Z(n32068) );
  XNOR U10088 ( .A(n32069), .B(n31637), .Z(n31639) );
  XNOR U10089 ( .A(n31640), .B(n31202), .Z(n31204) );
  XNOR U10090 ( .A(n31205), .B(n30761), .Z(n30763) );
  XNOR U10091 ( .A(n30764), .B(n30314), .Z(n30316) );
  XNOR U10092 ( .A(n30317), .B(n29861), .Z(n29863) );
  XNOR U10093 ( .A(n29864), .B(n29402), .Z(n29404) );
  XNOR U10094 ( .A(n29405), .B(n28937), .Z(n28939) );
  XNOR U10095 ( .A(n28940), .B(n28466), .Z(n28468) );
  XNOR U10096 ( .A(n28469), .B(n27989), .Z(n27991) );
  XNOR U10097 ( .A(n27992), .B(n27506), .Z(n27508) );
  XNOR U10098 ( .A(n27509), .B(n27017), .Z(n27019) );
  XNOR U10099 ( .A(n27020), .B(n26520), .Z(n26522) );
  XNOR U10100 ( .A(n26523), .B(n26019), .Z(n26021) );
  XNOR U10101 ( .A(n26022), .B(n25511), .Z(n25513) );
  XNOR U10102 ( .A(n25514), .B(n24997), .Z(n24999) );
  XNOR U10103 ( .A(n24477), .B(n23949), .Z(n23951) );
  XNOR U10104 ( .A(n23952), .B(n23418), .Z(n23420) );
  XNOR U10105 ( .A(n24472), .B(n23944), .Z(n23946) );
  XNOR U10106 ( .A(n23937), .B(n23403), .Z(n23405) );
  XNOR U10107 ( .A(n22848), .B(n22301), .Z(n22303) );
  XNOR U10108 ( .A(n22294), .B(n21742), .Z(n21744) );
  XNOR U10109 ( .A(n21105), .B(n20540), .Z(n20542) );
  XNOR U10110 ( .A(n19373), .B(n18791), .Z(n18793) );
  XNOR U10111 ( .A(n22828), .B(n22281), .Z(n22283) );
  XNOR U10112 ( .A(n21150), .B(n20585), .Z(n20587) );
  XNOR U10113 ( .A(n22853), .B(n22306), .Z(n22308) );
  XNOR U10114 ( .A(n21175), .B(n20610), .Z(n20612) );
  XNOR U10115 ( .A(n22254), .B(n21702), .Z(n21704) );
  XNOR U10116 ( .A(n21130), .B(n20565), .Z(n20567) );
  XNOR U10117 ( .A(n20558), .B(n19988), .Z(n19990) );
  XNOR U10118 ( .A(n19398), .B(n18816), .Z(n18818) );
  XNOR U10119 ( .A(n21110), .B(n20545), .Z(n20547) );
  XNOR U10120 ( .A(n19378), .B(n18796), .Z(n18798) );
  XNOR U10121 ( .A(n22833), .B(n22286), .Z(n22288) );
  XNOR U10122 ( .A(n21155), .B(n20590), .Z(n20592) );
  XNOR U10123 ( .A(n22878), .B(n22331), .Z(n22333) );
  XNOR U10124 ( .A(n22324), .B(n21772), .Z(n21774) );
  XNOR U10125 ( .A(n21135), .B(n20570), .Z(n20572) );
  XNOR U10126 ( .A(n19403), .B(n18821), .Z(n18823) );
  XNOR U10127 ( .A(n19383), .B(n18801), .Z(n18803) );
  XNOR U10128 ( .A(n21160), .B(n20595), .Z(n20597) );
  XNOR U10129 ( .A(n19428), .B(n18846), .Z(n18848) );
  XNOR U10130 ( .A(n22883), .B(n22336), .Z(n22338) );
  XNOR U10131 ( .A(n21205), .B(n20640), .Z(n20642) );
  XNOR U10132 ( .A(n36044), .B(n35672), .Z(n35674) );
  XNOR U10133 ( .A(n35675), .B(n35297), .Z(n35299) );
  XNOR U10134 ( .A(n35300), .B(n34916), .Z(n34918) );
  XNOR U10135 ( .A(n34919), .B(n34529), .Z(n34531) );
  XNOR U10136 ( .A(n34532), .B(n34136), .Z(n34138) );
  XNOR U10137 ( .A(n34139), .B(n33737), .Z(n33739) );
  XNOR U10138 ( .A(n33740), .B(n33332), .Z(n33334) );
  XNOR U10139 ( .A(n33335), .B(n32921), .Z(n32923) );
  XNOR U10140 ( .A(n32924), .B(n32504), .Z(n32506) );
  XNOR U10141 ( .A(n32507), .B(n32081), .Z(n32083) );
  XNOR U10142 ( .A(n32084), .B(n31652), .Z(n31654) );
  XNOR U10143 ( .A(n31655), .B(n31217), .Z(n31219) );
  XNOR U10144 ( .A(n31220), .B(n30776), .Z(n30778) );
  XNOR U10145 ( .A(n30779), .B(n30329), .Z(n30331) );
  XNOR U10146 ( .A(n30332), .B(n29876), .Z(n29878) );
  XNOR U10147 ( .A(n29879), .B(n29417), .Z(n29419) );
  XNOR U10148 ( .A(n29420), .B(n28952), .Z(n28954) );
  XNOR U10149 ( .A(n28955), .B(n28481), .Z(n28483) );
  XNOR U10150 ( .A(n28484), .B(n28004), .Z(n28006) );
  XNOR U10151 ( .A(n28007), .B(n27521), .Z(n27523) );
  XNOR U10152 ( .A(n27524), .B(n27032), .Z(n27034) );
  XNOR U10153 ( .A(n27035), .B(n26535), .Z(n26537) );
  XNOR U10154 ( .A(n26538), .B(n26034), .Z(n26036) );
  XNOR U10155 ( .A(n26037), .B(n25526), .Z(n25528) );
  XNOR U10156 ( .A(n25529), .B(n25012), .Z(n25014) );
  XNOR U10157 ( .A(n25015), .B(n24489), .Z(n24491) );
  XNOR U10158 ( .A(n24492), .B(n23964), .Z(n23966) );
  XNOR U10159 ( .A(n22898), .B(n22351), .Z(n22353) );
  XNOR U10160 ( .A(n22354), .B(n21802), .Z(n21804) );
  XNOR U10161 ( .A(n22863), .B(n22316), .Z(n22318) );
  XNOR U10162 ( .A(n22309), .B(n21757), .Z(n21759) );
  XNOR U10163 ( .A(n21185), .B(n20620), .Z(n20622) );
  XNOR U10164 ( .A(n20613), .B(n20043), .Z(n20045) );
  XNOR U10165 ( .A(n19388), .B(n18806), .Z(n18808) );
  XNOR U10166 ( .A(n21165), .B(n20600), .Z(n20602) );
  XNOR U10167 ( .A(n19433), .B(n18851), .Z(n18853) );
  XNOR U10168 ( .A(n22888), .B(n22341), .Z(n22343) );
  XNOR U10169 ( .A(n21235), .B(n20670), .Z(n20672) );
  XNOR U10170 ( .A(n21190), .B(n20625), .Z(n20627) );
  XNOR U10171 ( .A(n19458), .B(n18876), .Z(n18878) );
  XNOR U10172 ( .A(n20573), .B(n20003), .Z(n20005) );
  XNOR U10173 ( .A(n19413), .B(n18831), .Z(n18833) );
  XNOR U10174 ( .A(n19393), .B(n18811), .Z(n18813) );
  XOR U10175 ( .A(n17502), .B(n18087), .Z(n17506) );
  XNOR U10176 ( .A(n21170), .B(n20605), .Z(n20607) );
  XNOR U10177 ( .A(n19438), .B(n18856), .Z(n18858) );
  XNOR U10178 ( .A(n22893), .B(n22346), .Z(n22348) );
  XNOR U10179 ( .A(n21215), .B(n20650), .Z(n20652) );
  XNOR U10180 ( .A(n20643), .B(n20073), .Z(n20075) );
  XNOR U10181 ( .A(n19418), .B(n18836), .Z(n18838) );
  XOR U10182 ( .A(n18129), .B(n18767), .Z(n18133) );
  XOR U10183 ( .A(n16285), .B(n16888), .Z(n16289) );
  XNOR U10184 ( .A(n19443), .B(n18861), .Z(n18863) );
  XNOR U10185 ( .A(n21220), .B(n20655), .Z(n20657) );
  XNOR U10186 ( .A(n19488), .B(n18906), .Z(n18908) );
  XNOR U10187 ( .A(n37130), .B(n36776), .Z(n36778) );
  XNOR U10188 ( .A(n36779), .B(n36419), .Z(n36421) );
  XNOR U10189 ( .A(n36422), .B(n36056), .Z(n36058) );
  XNOR U10190 ( .A(n36059), .B(n35687), .Z(n35689) );
  XNOR U10191 ( .A(n35690), .B(n35312), .Z(n35314) );
  XNOR U10192 ( .A(n35315), .B(n34931), .Z(n34933) );
  XNOR U10193 ( .A(n34934), .B(n34544), .Z(n34546) );
  XNOR U10194 ( .A(n34547), .B(n34151), .Z(n34153) );
  XNOR U10195 ( .A(n34154), .B(n33752), .Z(n33754) );
  XNOR U10196 ( .A(n33755), .B(n33347), .Z(n33349) );
  XNOR U10197 ( .A(n33350), .B(n32936), .Z(n32938) );
  XNOR U10198 ( .A(n32939), .B(n32519), .Z(n32521) );
  XNOR U10199 ( .A(n32522), .B(n32096), .Z(n32098) );
  XNOR U10200 ( .A(n32099), .B(n31667), .Z(n31669) );
  XNOR U10201 ( .A(n31670), .B(n31232), .Z(n31234) );
  XNOR U10202 ( .A(n31235), .B(n30791), .Z(n30793) );
  XNOR U10203 ( .A(n30794), .B(n30344), .Z(n30346) );
  XNOR U10204 ( .A(n30347), .B(n29891), .Z(n29893) );
  XNOR U10205 ( .A(n29894), .B(n29432), .Z(n29434) );
  XNOR U10206 ( .A(n29435), .B(n28967), .Z(n28969) );
  XNOR U10207 ( .A(n28970), .B(n28496), .Z(n28498) );
  XNOR U10208 ( .A(n28499), .B(n28019), .Z(n28021) );
  XNOR U10209 ( .A(n28022), .B(n27536), .Z(n27538) );
  XNOR U10210 ( .A(n27539), .B(n27047), .Z(n27049) );
  XNOR U10211 ( .A(n27050), .B(n26550), .Z(n26552) );
  XNOR U10212 ( .A(n26553), .B(n26049), .Z(n26051) );
  XNOR U10213 ( .A(n26052), .B(n25541), .Z(n25543) );
  XNOR U10214 ( .A(n25544), .B(n25027), .Z(n25029) );
  XNOR U10215 ( .A(n25030), .B(n24504), .Z(n24506) );
  XNOR U10216 ( .A(n24507), .B(n23979), .Z(n23981) );
  XNOR U10217 ( .A(n23982), .B(n23448), .Z(n23450) );
  XNOR U10218 ( .A(n23451), .B(n22910), .Z(n22912) );
  XNOR U10219 ( .A(n22913), .B(n22366), .Z(n22368) );
  XNOR U10220 ( .A(n21265), .B(n20700), .Z(n20702) );
  XNOR U10221 ( .A(n21245), .B(n20680), .Z(n20682) );
  XNOR U10222 ( .A(n20673), .B(n20103), .Z(n20105) );
  XNOR U10223 ( .A(n21200), .B(n20635), .Z(n20637) );
  XNOR U10224 ( .A(n20628), .B(n20058), .Z(n20060) );
  XNOR U10225 ( .A(n19468), .B(n18886), .Z(n18888) );
  XOR U10226 ( .A(n16924), .B(n17485), .Z(n16928) );
  XNOR U10227 ( .A(n19448), .B(n18866), .Z(n18868) );
  XOR U10228 ( .A(n17557), .B(n18076), .Z(n17561) );
  XNOR U10229 ( .A(n21225), .B(n20660), .Z(n20662) );
  XNOR U10230 ( .A(n21250), .B(n20685), .Z(n20687) );
  XNOR U10231 ( .A(n19518), .B(n18936), .Z(n18938) );
  XOR U10232 ( .A(n18184), .B(n18745), .Z(n18188) );
  XNOR U10233 ( .A(n19473), .B(n18891), .Z(n18893) );
  XOR U10234 ( .A(n17517), .B(n18084), .Z(n17521) );
  XNOR U10235 ( .A(n19453), .B(n18871), .Z(n18873) );
  XNOR U10236 ( .A(n21230), .B(n20665), .Z(n20667) );
  XNOR U10237 ( .A(n19498), .B(n18916), .Z(n18918) );
  XNOR U10238 ( .A(n20703), .B(n20133), .Z(n20135) );
  XNOR U10239 ( .A(n21255), .B(n20690), .Z(n20692) );
  XOR U10240 ( .A(n18144), .B(n18761), .Z(n18148) );
  XOR U10241 ( .A(n16300), .B(n16885), .Z(n16304) );
  XOR U10242 ( .A(n15054), .B(n15663), .Z(n15058) );
  XOR U10243 ( .A(n18214), .B(n18733), .Z(n18218) );
  XNOR U10244 ( .A(n19503), .B(n18921), .Z(n18923) );
  XNOR U10245 ( .A(n19548), .B(n18966), .Z(n18968) );
  XNOR U10246 ( .A(n38162), .B(n37826), .Z(n37828) );
  XNOR U10247 ( .A(n37829), .B(n37487), .Z(n37489) );
  XNOR U10248 ( .A(n37490), .B(n37142), .Z(n37144) );
  XNOR U10249 ( .A(n37145), .B(n36791), .Z(n36793) );
  XNOR U10250 ( .A(n36794), .B(n36434), .Z(n36436) );
  XNOR U10251 ( .A(n36437), .B(n36071), .Z(n36073) );
  XNOR U10252 ( .A(n36074), .B(n35702), .Z(n35704) );
  XNOR U10253 ( .A(n35705), .B(n35327), .Z(n35329) );
  XNOR U10254 ( .A(n35330), .B(n34946), .Z(n34948) );
  XNOR U10255 ( .A(n34949), .B(n34559), .Z(n34561) );
  XNOR U10256 ( .A(n34562), .B(n34166), .Z(n34168) );
  XNOR U10257 ( .A(n34169), .B(n33767), .Z(n33769) );
  XNOR U10258 ( .A(n33770), .B(n33362), .Z(n33364) );
  XNOR U10259 ( .A(n33365), .B(n32951), .Z(n32953) );
  XNOR U10260 ( .A(n32954), .B(n32534), .Z(n32536) );
  XNOR U10261 ( .A(n32537), .B(n32111), .Z(n32113) );
  XNOR U10262 ( .A(n32114), .B(n31682), .Z(n31684) );
  XNOR U10263 ( .A(n31685), .B(n31247), .Z(n31249) );
  XNOR U10264 ( .A(n31250), .B(n30806), .Z(n30808) );
  XNOR U10265 ( .A(n30809), .B(n30359), .Z(n30361) );
  XNOR U10266 ( .A(n30362), .B(n29906), .Z(n29908) );
  XNOR U10267 ( .A(n29909), .B(n29447), .Z(n29449) );
  XNOR U10268 ( .A(n29450), .B(n28982), .Z(n28984) );
  XNOR U10269 ( .A(n28985), .B(n28511), .Z(n28513) );
  XNOR U10270 ( .A(n28514), .B(n28034), .Z(n28036) );
  XNOR U10271 ( .A(n28037), .B(n27551), .Z(n27553) );
  XNOR U10272 ( .A(n27554), .B(n27062), .Z(n27064) );
  XNOR U10273 ( .A(n27065), .B(n26565), .Z(n26567) );
  XNOR U10274 ( .A(n26568), .B(n26064), .Z(n26066) );
  XNOR U10275 ( .A(n26067), .B(n25556), .Z(n25558) );
  XNOR U10276 ( .A(n25559), .B(n25042), .Z(n25044) );
  XNOR U10277 ( .A(n25045), .B(n24519), .Z(n24521) );
  XNOR U10278 ( .A(n24522), .B(n23994), .Z(n23996) );
  XNOR U10279 ( .A(n23997), .B(n23463), .Z(n23465) );
  XNOR U10280 ( .A(n23466), .B(n22925), .Z(n22927) );
  XNOR U10281 ( .A(n22928), .B(n22381), .Z(n22383) );
  XNOR U10282 ( .A(n22384), .B(n21832), .Z(n21834) );
  XNOR U10283 ( .A(n21835), .B(n21277), .Z(n21279) );
  XNOR U10284 ( .A(n21280), .B(n20715), .Z(n20717) );
  XNOR U10285 ( .A(n21260), .B(n20695), .Z(n20697) );
  XNOR U10286 ( .A(n19528), .B(n18946), .Z(n18948) );
  XNOR U10287 ( .A(n19483), .B(n18901), .Z(n18903) );
  XOR U10288 ( .A(n16939), .B(n17482), .Z(n16943) );
  XOR U10289 ( .A(n15705), .B(n16272), .Z(n15709) );
  XOR U10290 ( .A(n13789), .B(n14416), .Z(n13793) );
  XOR U10291 ( .A(n17572), .B(n18073), .Z(n17576) );
  XOR U10292 ( .A(n16350), .B(n16875), .Z(n16354) );
  XNOR U10293 ( .A(n19508), .B(n18926), .Z(n18928) );
  XNOR U10294 ( .A(n19578), .B(n18996), .Z(n18998) );
  XOR U10295 ( .A(n18244), .B(n18721), .Z(n18248) );
  XNOR U10296 ( .A(n19533), .B(n18951), .Z(n18953) );
  XOR U10297 ( .A(n18199), .B(n18739), .Z(n18203) );
  XOR U10298 ( .A(n16989), .B(n17472), .Z(n16993) );
  XOR U10299 ( .A(n14452), .B(n15037), .Z(n14456) );
  XOR U10300 ( .A(n15109), .B(n15652), .Z(n15113) );
  XNOR U10301 ( .A(n19513), .B(n18931), .Z(n18933) );
  XNOR U10302 ( .A(n19558), .B(n18976), .Z(n18978) );
  XNOR U10303 ( .A(n19538), .B(n18956), .Z(n18958) );
  XOR U10304 ( .A(n15069), .B(n15660), .Z(n15073) );
  XOR U10305 ( .A(n17627), .B(n18062), .Z(n17631) );
  XOR U10306 ( .A(n16405), .B(n16864), .Z(n16409) );
  XOR U10307 ( .A(n18274), .B(n18709), .Z(n18278) );
  XNOR U10308 ( .A(n19563), .B(n18981), .Z(n18983) );
  XNOR U10309 ( .A(n39140), .B(n38822), .Z(n38824) );
  XNOR U10310 ( .A(n38825), .B(n38501), .Z(n38503) );
  XNOR U10311 ( .A(n38504), .B(n38174), .Z(n38176) );
  XNOR U10312 ( .A(n38177), .B(n37841), .Z(n37843) );
  XNOR U10313 ( .A(n37844), .B(n37502), .Z(n37504) );
  XNOR U10314 ( .A(n37505), .B(n37157), .Z(n37159) );
  XNOR U10315 ( .A(n37160), .B(n36806), .Z(n36808) );
  XNOR U10316 ( .A(n36809), .B(n36449), .Z(n36451) );
  XNOR U10317 ( .A(n36452), .B(n36086), .Z(n36088) );
  XNOR U10318 ( .A(n36089), .B(n35717), .Z(n35719) );
  XNOR U10319 ( .A(n35720), .B(n35342), .Z(n35344) );
  XNOR U10320 ( .A(n35345), .B(n34961), .Z(n34963) );
  XNOR U10321 ( .A(n34964), .B(n34574), .Z(n34576) );
  XNOR U10322 ( .A(n34577), .B(n34181), .Z(n34183) );
  XNOR U10323 ( .A(n34184), .B(n33782), .Z(n33784) );
  XNOR U10324 ( .A(n33785), .B(n33377), .Z(n33379) );
  XNOR U10325 ( .A(n33380), .B(n32966), .Z(n32968) );
  XNOR U10326 ( .A(n32969), .B(n32549), .Z(n32551) );
  XNOR U10327 ( .A(n32552), .B(n32126), .Z(n32128) );
  XNOR U10328 ( .A(n32129), .B(n31697), .Z(n31699) );
  XNOR U10329 ( .A(n31700), .B(n31262), .Z(n31264) );
  XNOR U10330 ( .A(n31265), .B(n30821), .Z(n30823) );
  XNOR U10331 ( .A(n30824), .B(n30374), .Z(n30376) );
  XNOR U10332 ( .A(n30377), .B(n29921), .Z(n29923) );
  XNOR U10333 ( .A(n29924), .B(n29462), .Z(n29464) );
  XNOR U10334 ( .A(n29465), .B(n28997), .Z(n28999) );
  XNOR U10335 ( .A(n29000), .B(n28526), .Z(n28528) );
  XNOR U10336 ( .A(n28529), .B(n28049), .Z(n28051) );
  XNOR U10337 ( .A(n28052), .B(n27566), .Z(n27568) );
  XNOR U10338 ( .A(n27569), .B(n27077), .Z(n27079) );
  XNOR U10339 ( .A(n27080), .B(n26580), .Z(n26582) );
  XNOR U10340 ( .A(n26583), .B(n26079), .Z(n26081) );
  XNOR U10341 ( .A(n26082), .B(n25571), .Z(n25573) );
  XNOR U10342 ( .A(n25574), .B(n25057), .Z(n25059) );
  XNOR U10343 ( .A(n25060), .B(n24534), .Z(n24536) );
  XNOR U10344 ( .A(n24537), .B(n24009), .Z(n24011) );
  XNOR U10345 ( .A(n24012), .B(n23478), .Z(n23480) );
  XNOR U10346 ( .A(n23481), .B(n22940), .Z(n22942) );
  XNOR U10347 ( .A(n22943), .B(n22396), .Z(n22398) );
  XNOR U10348 ( .A(n22399), .B(n21847), .Z(n21849) );
  XNOR U10349 ( .A(n21850), .B(n21292), .Z(n21294) );
  XNOR U10350 ( .A(n21295), .B(n20730), .Z(n20732) );
  XNOR U10351 ( .A(n20733), .B(n20163), .Z(n20165) );
  XNOR U10352 ( .A(n19588), .B(n19006), .Z(n19008) );
  XNOR U10353 ( .A(n19543), .B(n18961), .Z(n18963) );
  XOR U10354 ( .A(n15720), .B(n16269), .Z(n15724) );
  XOR U10355 ( .A(n13804), .B(n14413), .Z(n13808) );
  XOR U10356 ( .A(n12510), .B(n13143), .Z(n12514) );
  XOR U10357 ( .A(n16365), .B(n16872), .Z(n16369) );
  XNOR U10358 ( .A(n19568), .B(n18986), .Z(n18988) );
  XOR U10359 ( .A(n18304), .B(n18697), .Z(n18308) );
  XNOR U10360 ( .A(n19593), .B(n19011), .Z(n19013) );
  XOR U10361 ( .A(n17657), .B(n18056), .Z(n17661) );
  XOR U10362 ( .A(n16435), .B(n16858), .Z(n16439) );
  XOR U10363 ( .A(n17004), .B(n17469), .Z(n17008) );
  XOR U10364 ( .A(n15770), .B(n16259), .Z(n15774) );
  XOR U10365 ( .A(n14512), .B(n15025), .Z(n14516) );
  XOR U10366 ( .A(n14467), .B(n15034), .Z(n14471) );
  XOR U10367 ( .A(n13185), .B(n13776), .Z(n13189) );
  XOR U10368 ( .A(n11195), .B(n11846), .Z(n11199) );
  XOR U10369 ( .A(n15124), .B(n15649), .Z(n15128) );
  XOR U10370 ( .A(n13854), .B(n14403), .Z(n13858) );
  XNOR U10371 ( .A(n19573), .B(n18991), .Z(n18993) );
  XOR U10372 ( .A(n11882), .B(n12493), .Z(n11886) );
  XOR U10373 ( .A(n12565), .B(n13132), .Z(n12569) );
  XOR U10374 ( .A(n17034), .B(n17463), .Z(n17038) );
  XOR U10375 ( .A(n15800), .B(n16253), .Z(n15804) );
  XOR U10376 ( .A(n14542), .B(n15019), .Z(n14546) );
  XOR U10377 ( .A(n17687), .B(n18050), .Z(n17691) );
  XOR U10378 ( .A(n16465), .B(n16852), .Z(n16469) );
  XNOR U10379 ( .A(n40064), .B(n39764), .Z(n39766) );
  XNOR U10380 ( .A(n39767), .B(n39461), .Z(n39463) );
  XNOR U10381 ( .A(n39464), .B(n39152), .Z(n39154) );
  XNOR U10382 ( .A(n39155), .B(n38837), .Z(n38839) );
  XNOR U10383 ( .A(n38840), .B(n38516), .Z(n38518) );
  XNOR U10384 ( .A(n38519), .B(n38189), .Z(n38191) );
  XNOR U10385 ( .A(n38192), .B(n37856), .Z(n37858) );
  XNOR U10386 ( .A(n37859), .B(n37517), .Z(n37519) );
  XNOR U10387 ( .A(n37520), .B(n37172), .Z(n37174) );
  XNOR U10388 ( .A(n37175), .B(n36821), .Z(n36823) );
  XNOR U10389 ( .A(n36824), .B(n36464), .Z(n36466) );
  XNOR U10390 ( .A(n36467), .B(n36101), .Z(n36103) );
  XNOR U10391 ( .A(n36104), .B(n35732), .Z(n35734) );
  XNOR U10392 ( .A(n35735), .B(n35357), .Z(n35359) );
  XNOR U10393 ( .A(n35360), .B(n34976), .Z(n34978) );
  XNOR U10394 ( .A(n34979), .B(n34589), .Z(n34591) );
  XNOR U10395 ( .A(n34592), .B(n34196), .Z(n34198) );
  XNOR U10396 ( .A(n34199), .B(n33797), .Z(n33799) );
  XNOR U10397 ( .A(n33800), .B(n33392), .Z(n33394) );
  XNOR U10398 ( .A(n33395), .B(n32981), .Z(n32983) );
  XNOR U10399 ( .A(n32984), .B(n32564), .Z(n32566) );
  XNOR U10400 ( .A(n32567), .B(n32141), .Z(n32143) );
  XNOR U10401 ( .A(n32144), .B(n31712), .Z(n31714) );
  XNOR U10402 ( .A(n31715), .B(n31277), .Z(n31279) );
  XNOR U10403 ( .A(n31280), .B(n30836), .Z(n30838) );
  XNOR U10404 ( .A(n30839), .B(n30389), .Z(n30391) );
  XNOR U10405 ( .A(n30392), .B(n29936), .Z(n29938) );
  XNOR U10406 ( .A(n29939), .B(n29477), .Z(n29479) );
  XNOR U10407 ( .A(n29480), .B(n29012), .Z(n29014) );
  XNOR U10408 ( .A(n29015), .B(n28541), .Z(n28543) );
  XNOR U10409 ( .A(n28544), .B(n28064), .Z(n28066) );
  XNOR U10410 ( .A(n28067), .B(n27581), .Z(n27583) );
  XNOR U10411 ( .A(n27584), .B(n27092), .Z(n27094) );
  XNOR U10412 ( .A(n27095), .B(n26595), .Z(n26597) );
  XNOR U10413 ( .A(n26598), .B(n26094), .Z(n26096) );
  XNOR U10414 ( .A(n26097), .B(n25586), .Z(n25588) );
  XNOR U10415 ( .A(n25589), .B(n25072), .Z(n25074) );
  XNOR U10416 ( .A(n25075), .B(n24549), .Z(n24551) );
  XNOR U10417 ( .A(n24552), .B(n24024), .Z(n24026) );
  XNOR U10418 ( .A(n24027), .B(n23493), .Z(n23495) );
  XNOR U10419 ( .A(n23496), .B(n22955), .Z(n22957) );
  XNOR U10420 ( .A(n22958), .B(n22411), .Z(n22413) );
  XNOR U10421 ( .A(n22414), .B(n21862), .Z(n21864) );
  XNOR U10422 ( .A(n21865), .B(n21307), .Z(n21309) );
  XNOR U10423 ( .A(n21310), .B(n20745), .Z(n20747) );
  XNOR U10424 ( .A(n20748), .B(n20178), .Z(n20180) );
  XNOR U10425 ( .A(n19608), .B(n19026), .Z(n19028) );
  XNOR U10426 ( .A(n19603), .B(n19021), .Z(n19023) );
  XOR U10427 ( .A(n12525), .B(n13140), .Z(n12529) );
  XOR U10428 ( .A(n17717), .B(n18044), .Z(n17721) );
  XOR U10429 ( .A(n16495), .B(n16846), .Z(n16499) );
  XOR U10430 ( .A(n17064), .B(n17457), .Z(n17068) );
  XOR U10431 ( .A(n15830), .B(n16247), .Z(n15834) );
  XOR U10432 ( .A(n14572), .B(n15013), .Z(n14576) );
  XOR U10433 ( .A(n15159), .B(n15642), .Z(n15163) );
  XOR U10434 ( .A(n13889), .B(n14396), .Z(n13893) );
  XOR U10435 ( .A(n12595), .B(n13126), .Z(n12599) );
  XOR U10436 ( .A(n13200), .B(n13773), .Z(n13204) );
  XOR U10437 ( .A(n11210), .B(n11843), .Z(n11214) );
  XOR U10438 ( .A(n9868), .B(n10525), .Z(n9872) );
  XOR U10439 ( .A(n13869), .B(n14400), .Z(n13873) );
  XOR U10440 ( .A(n17742), .B(n18039), .Z(n17746) );
  XOR U10441 ( .A(n11897), .B(n12490), .Z(n11901) );
  XOR U10442 ( .A(n10567), .B(n11182), .Z(n10571) );
  XOR U10443 ( .A(n8507), .B(n9182), .Z(n8511) );
  XOR U10444 ( .A(n12580), .B(n13129), .Z(n12584) );
  XOR U10445 ( .A(n11260), .B(n11833), .Z(n11264) );
  XOR U10446 ( .A(n15189), .B(n15636), .Z(n15193) );
  XOR U10447 ( .A(n13919), .B(n14390), .Z(n13923) );
  XOR U10448 ( .A(n12625), .B(n13120), .Z(n12629) );
  XOR U10449 ( .A(n17094), .B(n17451), .Z(n17098) );
  XOR U10450 ( .A(n15860), .B(n16241), .Z(n15864) );
  XOR U10451 ( .A(n14602), .B(n15007), .Z(n14606) );
  XOR U10452 ( .A(n16525), .B(n16840), .Z(n16529) );
  XNOR U10453 ( .A(n40934), .B(n40652), .Z(n40654) );
  XNOR U10454 ( .A(n40655), .B(n40367), .Z(n40369) );
  XNOR U10455 ( .A(n40370), .B(n40076), .Z(n40078) );
  XNOR U10456 ( .A(n40079), .B(n39779), .Z(n39781) );
  XNOR U10457 ( .A(n39782), .B(n39476), .Z(n39478) );
  XNOR U10458 ( .A(n39479), .B(n39167), .Z(n39169) );
  XNOR U10459 ( .A(n39170), .B(n38852), .Z(n38854) );
  XNOR U10460 ( .A(n38855), .B(n38531), .Z(n38533) );
  XNOR U10461 ( .A(n38534), .B(n38204), .Z(n38206) );
  XNOR U10462 ( .A(n38207), .B(n37871), .Z(n37873) );
  XNOR U10463 ( .A(n37874), .B(n37532), .Z(n37534) );
  XNOR U10464 ( .A(n37535), .B(n37187), .Z(n37189) );
  XNOR U10465 ( .A(n37190), .B(n36836), .Z(n36838) );
  XNOR U10466 ( .A(n36839), .B(n36479), .Z(n36481) );
  XNOR U10467 ( .A(n36482), .B(n36116), .Z(n36118) );
  XNOR U10468 ( .A(n36119), .B(n35747), .Z(n35749) );
  XNOR U10469 ( .A(n35750), .B(n35372), .Z(n35374) );
  XNOR U10470 ( .A(n35375), .B(n34991), .Z(n34993) );
  XNOR U10471 ( .A(n34994), .B(n34604), .Z(n34606) );
  XNOR U10472 ( .A(n34607), .B(n34211), .Z(n34213) );
  XNOR U10473 ( .A(n34214), .B(n33812), .Z(n33814) );
  XNOR U10474 ( .A(n33815), .B(n33407), .Z(n33409) );
  XNOR U10475 ( .A(n33410), .B(n32996), .Z(n32998) );
  XNOR U10476 ( .A(n32999), .B(n32579), .Z(n32581) );
  XNOR U10477 ( .A(n32582), .B(n32156), .Z(n32158) );
  XNOR U10478 ( .A(n32159), .B(n31727), .Z(n31729) );
  XNOR U10479 ( .A(n31730), .B(n31292), .Z(n31294) );
  XNOR U10480 ( .A(n31295), .B(n30851), .Z(n30853) );
  XNOR U10481 ( .A(n30854), .B(n30404), .Z(n30406) );
  XNOR U10482 ( .A(n30407), .B(n29951), .Z(n29953) );
  XNOR U10483 ( .A(n29954), .B(n29492), .Z(n29494) );
  XNOR U10484 ( .A(n29495), .B(n29027), .Z(n29029) );
  XNOR U10485 ( .A(n29030), .B(n28556), .Z(n28558) );
  XNOR U10486 ( .A(n28559), .B(n28079), .Z(n28081) );
  XNOR U10487 ( .A(n28082), .B(n27596), .Z(n27598) );
  XNOR U10488 ( .A(n27599), .B(n27107), .Z(n27109) );
  XNOR U10489 ( .A(n27110), .B(n26610), .Z(n26612) );
  XNOR U10490 ( .A(n26613), .B(n26109), .Z(n26111) );
  XNOR U10491 ( .A(n26112), .B(n25601), .Z(n25603) );
  XNOR U10492 ( .A(n25604), .B(n25087), .Z(n25089) );
  XNOR U10493 ( .A(n25090), .B(n24564), .Z(n24566) );
  XNOR U10494 ( .A(n24567), .B(n24039), .Z(n24041) );
  XNOR U10495 ( .A(n24042), .B(n23508), .Z(n23510) );
  XNOR U10496 ( .A(n23511), .B(n22970), .Z(n22972) );
  XNOR U10497 ( .A(n22973), .B(n22426), .Z(n22428) );
  XNOR U10498 ( .A(n22429), .B(n21877), .Z(n21879) );
  XNOR U10499 ( .A(n21880), .B(n21322), .Z(n21324) );
  XNOR U10500 ( .A(n21325), .B(n20760), .Z(n20762) );
  XNOR U10501 ( .A(n20763), .B(n20193), .Z(n20195) );
  XNOR U10502 ( .A(n20196), .B(n19620), .Z(n19622) );
  XNOR U10503 ( .A(n19623), .B(n19041), .Z(n19043) );
  XOR U10504 ( .A(n18349), .B(n18679), .Z(n18353) );
  XOR U10505 ( .A(n9218), .B(n9851), .Z(n9222) );
  XOR U10506 ( .A(n16555), .B(n16834), .Z(n16559) );
  XOR U10507 ( .A(n17124), .B(n17445), .Z(n17128) );
  XOR U10508 ( .A(n15890), .B(n16235), .Z(n15894) );
  XOR U10509 ( .A(n14632), .B(n15001), .Z(n14636) );
  XOR U10510 ( .A(n15219), .B(n15630), .Z(n15223) );
  XOR U10511 ( .A(n13949), .B(n14384), .Z(n13953) );
  XOR U10512 ( .A(n12655), .B(n13114), .Z(n12659) );
  XOR U10513 ( .A(n13260), .B(n13761), .Z(n13264) );
  XOR U10514 ( .A(n11952), .B(n12479), .Z(n11956) );
  XOR U10515 ( .A(n10622), .B(n11171), .Z(n10626) );
  XOR U10516 ( .A(n9883), .B(n10522), .Z(n9887) );
  XOR U10517 ( .A(n10582), .B(n11179), .Z(n10586) );
  XOR U10518 ( .A(n8522), .B(n9179), .Z(n8526) );
  XOR U10519 ( .A(n7132), .B(n7813), .Z(n7136) );
  XOR U10520 ( .A(n11275), .B(n11830), .Z(n11279) );
  XOR U10521 ( .A(n9933), .B(n10512), .Z(n9937) );
  XOR U10522 ( .A(n8567), .B(n9170), .Z(n8571) );
  XOR U10523 ( .A(n13290), .B(n13755), .Z(n13294) );
  XOR U10524 ( .A(n11982), .B(n12473), .Z(n11986) );
  XOR U10525 ( .A(n10652), .B(n11165), .Z(n10656) );
  XOR U10526 ( .A(n15249), .B(n15624), .Z(n15253) );
  XOR U10527 ( .A(n13979), .B(n14378), .Z(n13983) );
  XOR U10528 ( .A(n12685), .B(n13108), .Z(n12689) );
  XOR U10529 ( .A(n17154), .B(n17439), .Z(n17158) );
  XOR U10530 ( .A(n15920), .B(n16229), .Z(n15924) );
  XOR U10531 ( .A(n14662), .B(n14995), .Z(n14666) );
  XNOR U10532 ( .A(n41750), .B(n41486), .Z(n41488) );
  XNOR U10533 ( .A(n41489), .B(n41219), .Z(n41221) );
  XNOR U10534 ( .A(n41222), .B(n40946), .Z(n40948) );
  XNOR U10535 ( .A(n40949), .B(n40667), .Z(n40669) );
  XNOR U10536 ( .A(n40670), .B(n40382), .Z(n40384) );
  XNOR U10537 ( .A(n40385), .B(n40091), .Z(n40093) );
  XNOR U10538 ( .A(n40094), .B(n39794), .Z(n39796) );
  XNOR U10539 ( .A(n39797), .B(n39491), .Z(n39493) );
  XNOR U10540 ( .A(n39494), .B(n39182), .Z(n39184) );
  XNOR U10541 ( .A(n39185), .B(n38867), .Z(n38869) );
  XNOR U10542 ( .A(n38870), .B(n38546), .Z(n38548) );
  XNOR U10543 ( .A(n38549), .B(n38219), .Z(n38221) );
  XNOR U10544 ( .A(n38222), .B(n37886), .Z(n37888) );
  XNOR U10545 ( .A(n37889), .B(n37547), .Z(n37549) );
  XNOR U10546 ( .A(n37550), .B(n37202), .Z(n37204) );
  XNOR U10547 ( .A(n37205), .B(n36851), .Z(n36853) );
  XNOR U10548 ( .A(n36854), .B(n36494), .Z(n36496) );
  XNOR U10549 ( .A(n36497), .B(n36131), .Z(n36133) );
  XNOR U10550 ( .A(n36134), .B(n35762), .Z(n35764) );
  XNOR U10551 ( .A(n35765), .B(n35387), .Z(n35389) );
  XNOR U10552 ( .A(n35390), .B(n35006), .Z(n35008) );
  XNOR U10553 ( .A(n35009), .B(n34619), .Z(n34621) );
  XNOR U10554 ( .A(n34622), .B(n34226), .Z(n34228) );
  XNOR U10555 ( .A(n34229), .B(n33827), .Z(n33829) );
  XNOR U10556 ( .A(n33830), .B(n33422), .Z(n33424) );
  XNOR U10557 ( .A(n33425), .B(n33011), .Z(n33013) );
  XNOR U10558 ( .A(n33014), .B(n32594), .Z(n32596) );
  XNOR U10559 ( .A(n32597), .B(n32171), .Z(n32173) );
  XNOR U10560 ( .A(n32174), .B(n31742), .Z(n31744) );
  XNOR U10561 ( .A(n31745), .B(n31307), .Z(n31309) );
  XNOR U10562 ( .A(n31310), .B(n30866), .Z(n30868) );
  XNOR U10563 ( .A(n30869), .B(n30419), .Z(n30421) );
  XNOR U10564 ( .A(n30422), .B(n29966), .Z(n29968) );
  XNOR U10565 ( .A(n29969), .B(n29507), .Z(n29509) );
  XNOR U10566 ( .A(n29510), .B(n29042), .Z(n29044) );
  XNOR U10567 ( .A(n29045), .B(n28571), .Z(n28573) );
  XNOR U10568 ( .A(n28574), .B(n28094), .Z(n28096) );
  XNOR U10569 ( .A(n28097), .B(n27611), .Z(n27613) );
  XNOR U10570 ( .A(n27614), .B(n27122), .Z(n27124) );
  XNOR U10571 ( .A(n27125), .B(n26625), .Z(n26627) );
  XNOR U10572 ( .A(n26628), .B(n26124), .Z(n26126) );
  XNOR U10573 ( .A(n26127), .B(n25616), .Z(n25618) );
  XNOR U10574 ( .A(n25619), .B(n25102), .Z(n25104) );
  XNOR U10575 ( .A(n25105), .B(n24579), .Z(n24581) );
  XNOR U10576 ( .A(n24582), .B(n24054), .Z(n24056) );
  XNOR U10577 ( .A(n24057), .B(n23523), .Z(n23525) );
  XNOR U10578 ( .A(n23526), .B(n22985), .Z(n22987) );
  XNOR U10579 ( .A(n22988), .B(n22441), .Z(n22443) );
  XNOR U10580 ( .A(n22444), .B(n21892), .Z(n21894) );
  XNOR U10581 ( .A(n21895), .B(n21337), .Z(n21339) );
  XNOR U10582 ( .A(n21340), .B(n20775), .Z(n20777) );
  XNOR U10583 ( .A(n20778), .B(n20208), .Z(n20210) );
  XNOR U10584 ( .A(n20211), .B(n19635), .Z(n19637) );
  XNOR U10585 ( .A(n19638), .B(n19056), .Z(n19058) );
  XOR U10586 ( .A(n17772), .B(n18033), .Z(n17776) );
  XOR U10587 ( .A(n9233), .B(n9848), .Z(n9237) );
  XOR U10588 ( .A(n7855), .B(n8494), .Z(n7859) );
  XOR U10589 ( .A(n5723), .B(n6422), .Z(n5727) );
  XOR U10590 ( .A(n15950), .B(n16223), .Z(n15954) );
  XOR U10591 ( .A(n14692), .B(n14989), .Z(n14696) );
  XOR U10592 ( .A(n15279), .B(n15618), .Z(n15283) );
  XOR U10593 ( .A(n14009), .B(n14372), .Z(n14013) );
  XOR U10594 ( .A(n12715), .B(n13102), .Z(n12719) );
  XOR U10595 ( .A(n13320), .B(n13749), .Z(n13324) );
  XOR U10596 ( .A(n12012), .B(n12467), .Z(n12016) );
  XOR U10597 ( .A(n10682), .B(n11159), .Z(n10686) );
  XOR U10598 ( .A(n11305), .B(n11824), .Z(n11309) );
  XOR U10599 ( .A(n9963), .B(n10506), .Z(n9967) );
  XOR U10600 ( .A(n8597), .B(n9164), .Z(n8601) );
  XOR U10601 ( .A(n6458), .B(n7115), .Z(n6462) );
  XOR U10602 ( .A(n7147), .B(n7810), .Z(n7151) );
  XOR U10603 ( .A(n9268), .B(n9841), .Z(n9272) );
  XOR U10604 ( .A(n7890), .B(n8487), .Z(n7894) );
  XOR U10605 ( .A(n6488), .B(n7109), .Z(n6492) );
  XOR U10606 ( .A(n11335), .B(n11818), .Z(n11339) );
  XOR U10607 ( .A(n9993), .B(n10500), .Z(n9997) );
  XOR U10608 ( .A(n8627), .B(n9158), .Z(n8631) );
  XOR U10609 ( .A(n13350), .B(n13743), .Z(n13354) );
  XOR U10610 ( .A(n12042), .B(n12461), .Z(n12046) );
  XOR U10611 ( .A(n10712), .B(n11153), .Z(n10716) );
  XOR U10612 ( .A(n15309), .B(n15612), .Z(n15313) );
  XOR U10613 ( .A(n14039), .B(n14366), .Z(n14043) );
  XOR U10614 ( .A(n12745), .B(n13096), .Z(n12749) );
  XOR U10615 ( .A(n14722), .B(n14983), .Z(n14726) );
  XNOR U10616 ( .A(n42512), .B(n42266), .Z(n42268) );
  XNOR U10617 ( .A(n42269), .B(n42017), .Z(n42019) );
  XNOR U10618 ( .A(n42020), .B(n41762), .Z(n41764) );
  XNOR U10619 ( .A(n41765), .B(n41501), .Z(n41503) );
  XNOR U10620 ( .A(n41504), .B(n41234), .Z(n41236) );
  XNOR U10621 ( .A(n41237), .B(n40961), .Z(n40963) );
  XNOR U10622 ( .A(n40964), .B(n40682), .Z(n40684) );
  XNOR U10623 ( .A(n40685), .B(n40397), .Z(n40399) );
  XNOR U10624 ( .A(n40400), .B(n40106), .Z(n40108) );
  XNOR U10625 ( .A(n40109), .B(n39809), .Z(n39811) );
  XNOR U10626 ( .A(n39812), .B(n39506), .Z(n39508) );
  XNOR U10627 ( .A(n39509), .B(n39197), .Z(n39199) );
  XNOR U10628 ( .A(n39200), .B(n38882), .Z(n38884) );
  XNOR U10629 ( .A(n38885), .B(n38561), .Z(n38563) );
  XNOR U10630 ( .A(n38564), .B(n38234), .Z(n38236) );
  XNOR U10631 ( .A(n38237), .B(n37901), .Z(n37903) );
  XNOR U10632 ( .A(n37904), .B(n37562), .Z(n37564) );
  XNOR U10633 ( .A(n37565), .B(n37217), .Z(n37219) );
  XNOR U10634 ( .A(n37220), .B(n36866), .Z(n36868) );
  XNOR U10635 ( .A(n36869), .B(n36509), .Z(n36511) );
  XNOR U10636 ( .A(n36512), .B(n36146), .Z(n36148) );
  XNOR U10637 ( .A(n36149), .B(n35777), .Z(n35779) );
  XNOR U10638 ( .A(n35780), .B(n35402), .Z(n35404) );
  XNOR U10639 ( .A(n35405), .B(n35021), .Z(n35023) );
  XNOR U10640 ( .A(n35024), .B(n34634), .Z(n34636) );
  XNOR U10641 ( .A(n34637), .B(n34241), .Z(n34243) );
  XNOR U10642 ( .A(n34244), .B(n33842), .Z(n33844) );
  XNOR U10643 ( .A(n33845), .B(n33437), .Z(n33439) );
  XNOR U10644 ( .A(n33440), .B(n33026), .Z(n33028) );
  XNOR U10645 ( .A(n33029), .B(n32609), .Z(n32611) );
  XNOR U10646 ( .A(n32612), .B(n32186), .Z(n32188) );
  XNOR U10647 ( .A(n32189), .B(n31757), .Z(n31759) );
  XNOR U10648 ( .A(n31760), .B(n31322), .Z(n31324) );
  XNOR U10649 ( .A(n31325), .B(n30881), .Z(n30883) );
  XNOR U10650 ( .A(n30884), .B(n30434), .Z(n30436) );
  XNOR U10651 ( .A(n30437), .B(n29981), .Z(n29983) );
  XNOR U10652 ( .A(n29984), .B(n29522), .Z(n29524) );
  XNOR U10653 ( .A(n29525), .B(n29057), .Z(n29059) );
  XNOR U10654 ( .A(n29060), .B(n28586), .Z(n28588) );
  XNOR U10655 ( .A(n28589), .B(n28109), .Z(n28111) );
  XNOR U10656 ( .A(n28112), .B(n27626), .Z(n27628) );
  XNOR U10657 ( .A(n27629), .B(n27137), .Z(n27139) );
  XNOR U10658 ( .A(n27140), .B(n26640), .Z(n26642) );
  XNOR U10659 ( .A(n26643), .B(n26139), .Z(n26141) );
  XNOR U10660 ( .A(n26142), .B(n25631), .Z(n25633) );
  XNOR U10661 ( .A(n25634), .B(n25117), .Z(n25119) );
  XNOR U10662 ( .A(n25120), .B(n24594), .Z(n24596) );
  XNOR U10663 ( .A(n24597), .B(n24069), .Z(n24071) );
  XNOR U10664 ( .A(n24072), .B(n23538), .Z(n23540) );
  XNOR U10665 ( .A(n23541), .B(n23000), .Z(n23002) );
  XNOR U10666 ( .A(n23003), .B(n22456), .Z(n22458) );
  XNOR U10667 ( .A(n22459), .B(n21907), .Z(n21909) );
  XNOR U10668 ( .A(n21910), .B(n21352), .Z(n21354) );
  XNOR U10669 ( .A(n21355), .B(n20790), .Z(n20792) );
  XNOR U10670 ( .A(n20793), .B(n20223), .Z(n20225) );
  XNOR U10671 ( .A(n20226), .B(n19650), .Z(n19652) );
  XNOR U10672 ( .A(n19653), .B(n19071), .Z(n19073) );
  XOR U10673 ( .A(n18379), .B(n18667), .Z(n18383) );
  XOR U10674 ( .A(n17189), .B(n17432), .Z(n17193) );
  XOR U10675 ( .A(n15975), .B(n16218), .Z(n15979) );
  XOR U10676 ( .A(n7870), .B(n8491), .Z(n7874) );
  XOR U10677 ( .A(n5738), .B(n6419), .Z(n5742) );
  XOR U10678 ( .A(n4298), .B(n5003), .Z(n4302) );
  XOR U10679 ( .A(n15339), .B(n15606), .Z(n15343) );
  XOR U10680 ( .A(n14069), .B(n14360), .Z(n14073) );
  XOR U10681 ( .A(n12775), .B(n13090), .Z(n12779) );
  XOR U10682 ( .A(n13380), .B(n13737), .Z(n13384) );
  XOR U10683 ( .A(n12072), .B(n12455), .Z(n12076) );
  XOR U10684 ( .A(n10742), .B(n11147), .Z(n10746) );
  XOR U10685 ( .A(n11365), .B(n11812), .Z(n11369) );
  XOR U10686 ( .A(n10023), .B(n10494), .Z(n10027) );
  XOR U10687 ( .A(n8657), .B(n9152), .Z(n8661) );
  XOR U10688 ( .A(n9298), .B(n9835), .Z(n9302) );
  XOR U10689 ( .A(n7920), .B(n8481), .Z(n7924) );
  XOR U10690 ( .A(n6518), .B(n7103), .Z(n6522) );
  XOR U10691 ( .A(n6473), .B(n7112), .Z(n6477) );
  XOR U10692 ( .A(n5045), .B(n5710), .Z(n5049) );
  XOR U10693 ( .A(n2841), .B(n3564), .Z(n2845) );
  XOR U10694 ( .A(n7207), .B(n7798), .Z(n7211) );
  XOR U10695 ( .A(n5793), .B(n6408), .Z(n5797) );
  XOR U10696 ( .A(n4353), .B(n4992), .Z(n4357) );
  XOR U10697 ( .A(n9328), .B(n9829), .Z(n9332) );
  XOR U10698 ( .A(n7950), .B(n8475), .Z(n7954) );
  XOR U10699 ( .A(n6548), .B(n7097), .Z(n6552) );
  XOR U10700 ( .A(n11395), .B(n11806), .Z(n11399) );
  XOR U10701 ( .A(n10053), .B(n10488), .Z(n10057) );
  XOR U10702 ( .A(n8687), .B(n9146), .Z(n8691) );
  XOR U10703 ( .A(n13410), .B(n13731), .Z(n13414) );
  XOR U10704 ( .A(n12102), .B(n12449), .Z(n12106) );
  XOR U10705 ( .A(n10772), .B(n11141), .Z(n10776) );
  XOR U10706 ( .A(n14099), .B(n14354), .Z(n14103) );
  XOR U10707 ( .A(n12805), .B(n13084), .Z(n12809) );
  XNOR U10708 ( .A(n43220), .B(n42992), .Z(n42994) );
  XNOR U10709 ( .A(n42995), .B(n42761), .Z(n42763) );
  XNOR U10710 ( .A(n42764), .B(n42524), .Z(n42526) );
  XNOR U10711 ( .A(n42527), .B(n42281), .Z(n42283) );
  XNOR U10712 ( .A(n42284), .B(n42032), .Z(n42034) );
  XNOR U10713 ( .A(n42035), .B(n41777), .Z(n41779) );
  XNOR U10714 ( .A(n41780), .B(n41516), .Z(n41518) );
  XNOR U10715 ( .A(n41519), .B(n41249), .Z(n41251) );
  XNOR U10716 ( .A(n41252), .B(n40976), .Z(n40978) );
  XNOR U10717 ( .A(n40979), .B(n40697), .Z(n40699) );
  XNOR U10718 ( .A(n40700), .B(n40412), .Z(n40414) );
  XNOR U10719 ( .A(n40415), .B(n40121), .Z(n40123) );
  XNOR U10720 ( .A(n40124), .B(n39824), .Z(n39826) );
  XNOR U10721 ( .A(n39827), .B(n39521), .Z(n39523) );
  XNOR U10722 ( .A(n39524), .B(n39212), .Z(n39214) );
  XNOR U10723 ( .A(n39215), .B(n38897), .Z(n38899) );
  XNOR U10724 ( .A(n38900), .B(n38576), .Z(n38578) );
  XNOR U10725 ( .A(n38579), .B(n38249), .Z(n38251) );
  XNOR U10726 ( .A(n38252), .B(n37916), .Z(n37918) );
  XNOR U10727 ( .A(n37919), .B(n37577), .Z(n37579) );
  XNOR U10728 ( .A(n37580), .B(n37232), .Z(n37234) );
  XNOR U10729 ( .A(n37235), .B(n36881), .Z(n36883) );
  XNOR U10730 ( .A(n36884), .B(n36524), .Z(n36526) );
  XNOR U10731 ( .A(n36527), .B(n36161), .Z(n36163) );
  XNOR U10732 ( .A(n36164), .B(n35792), .Z(n35794) );
  XNOR U10733 ( .A(n35795), .B(n35417), .Z(n35419) );
  XNOR U10734 ( .A(n35420), .B(n35036), .Z(n35038) );
  XNOR U10735 ( .A(n35039), .B(n34649), .Z(n34651) );
  XNOR U10736 ( .A(n34652), .B(n34256), .Z(n34258) );
  XNOR U10737 ( .A(n34259), .B(n33857), .Z(n33859) );
  XNOR U10738 ( .A(n33860), .B(n33452), .Z(n33454) );
  XNOR U10739 ( .A(n33455), .B(n33041), .Z(n33043) );
  XNOR U10740 ( .A(n33044), .B(n32624), .Z(n32626) );
  XNOR U10741 ( .A(n32627), .B(n32201), .Z(n32203) );
  XNOR U10742 ( .A(n32204), .B(n31772), .Z(n31774) );
  XNOR U10743 ( .A(n31775), .B(n31337), .Z(n31339) );
  XNOR U10744 ( .A(n31340), .B(n30896), .Z(n30898) );
  XNOR U10745 ( .A(n30899), .B(n30449), .Z(n30451) );
  XNOR U10746 ( .A(n30452), .B(n29996), .Z(n29998) );
  XNOR U10747 ( .A(n29999), .B(n29537), .Z(n29539) );
  XNOR U10748 ( .A(n29540), .B(n29072), .Z(n29074) );
  XNOR U10749 ( .A(n29075), .B(n28601), .Z(n28603) );
  XNOR U10750 ( .A(n28604), .B(n28124), .Z(n28126) );
  XNOR U10751 ( .A(n28127), .B(n27641), .Z(n27643) );
  XNOR U10752 ( .A(n27644), .B(n27152), .Z(n27154) );
  XNOR U10753 ( .A(n27155), .B(n26655), .Z(n26657) );
  XNOR U10754 ( .A(n26658), .B(n26154), .Z(n26156) );
  XNOR U10755 ( .A(n26157), .B(n25646), .Z(n25648) );
  XNOR U10756 ( .A(n25649), .B(n25132), .Z(n25134) );
  XNOR U10757 ( .A(n25135), .B(n24609), .Z(n24611) );
  XNOR U10758 ( .A(n24612), .B(n24084), .Z(n24086) );
  XNOR U10759 ( .A(n24087), .B(n23553), .Z(n23555) );
  XNOR U10760 ( .A(n23556), .B(n23015), .Z(n23017) );
  XNOR U10761 ( .A(n23018), .B(n22471), .Z(n22473) );
  XNOR U10762 ( .A(n22474), .B(n21922), .Z(n21924) );
  XNOR U10763 ( .A(n21925), .B(n21367), .Z(n21369) );
  XNOR U10764 ( .A(n21370), .B(n20805), .Z(n20807) );
  XNOR U10765 ( .A(n20808), .B(n20238), .Z(n20240) );
  XNOR U10766 ( .A(n20241), .B(n19665), .Z(n19667) );
  XNOR U10767 ( .A(n19668), .B(n19086), .Z(n19088) );
  XOR U10768 ( .A(n17802), .B(n18027), .Z(n17806) );
  XOR U10769 ( .A(n16600), .B(n16825), .Z(n16604) );
  XOR U10770 ( .A(n15374), .B(n15599), .Z(n15378) );
  XOR U10771 ( .A(n14124), .B(n14349), .Z(n14128) );
  XOR U10772 ( .A(n4313), .B(n5000), .Z(n4317) );
  XOR U10773 ( .A(n12835), .B(n13078), .Z(n12839) );
  XOR U10774 ( .A(n13440), .B(n13725), .Z(n13444) );
  XOR U10775 ( .A(n12132), .B(n12443), .Z(n12136) );
  XOR U10776 ( .A(n10802), .B(n11135), .Z(n10806) );
  XOR U10777 ( .A(n11425), .B(n11800), .Z(n11429) );
  XOR U10778 ( .A(n10083), .B(n10482), .Z(n10087) );
  XOR U10779 ( .A(n8717), .B(n9140), .Z(n8721) );
  XOR U10780 ( .A(n9358), .B(n9823), .Z(n9362) );
  XOR U10781 ( .A(n7980), .B(n8469), .Z(n7984) );
  XOR U10782 ( .A(n6578), .B(n7091), .Z(n6582) );
  XOR U10783 ( .A(n7237), .B(n7792), .Z(n7241) );
  XOR U10784 ( .A(n5823), .B(n6402), .Z(n5827) );
  XOR U10785 ( .A(n4383), .B(n4986), .Z(n4387) );
  XOR U10786 ( .A(n5060), .B(n5707), .Z(n5064) );
  XOR U10787 ( .A(n3610), .B(n4279), .Z(n3614) );
  XOR U10788 ( .A(n2136), .B(n2829), .Z(n2140) );
  XOR U10789 ( .A(n2856), .B(n3561), .Z(n2860) );
  XOR U10790 ( .A(n1370), .B(n2099), .Z(n1374) );
  XOR U10791 ( .A(n5090), .B(n5701), .Z(n5094) );
  XOR U10792 ( .A(n3640), .B(n4273), .Z(n3644) );
  XOR U10793 ( .A(n2166), .B(n2823), .Z(n2170) );
  XOR U10794 ( .A(n7267), .B(n7786), .Z(n7271) );
  XOR U10795 ( .A(n5853), .B(n6396), .Z(n5857) );
  XOR U10796 ( .A(n4413), .B(n4980), .Z(n4417) );
  XOR U10797 ( .A(n9388), .B(n9817), .Z(n9392) );
  XOR U10798 ( .A(n8010), .B(n8463), .Z(n8014) );
  XOR U10799 ( .A(n6608), .B(n7085), .Z(n6612) );
  XOR U10800 ( .A(n11455), .B(n11794), .Z(n11459) );
  XOR U10801 ( .A(n10113), .B(n10476), .Z(n10117) );
  XOR U10802 ( .A(n8747), .B(n9134), .Z(n8751) );
  XOR U10803 ( .A(n13470), .B(n13719), .Z(n13474) );
  XOR U10804 ( .A(n12162), .B(n12437), .Z(n12166) );
  XOR U10805 ( .A(n10832), .B(n11129), .Z(n10836) );
  XNOR U10806 ( .A(n43874), .B(n43664), .Z(n43666) );
  XNOR U10807 ( .A(n43667), .B(n43451), .Z(n43453) );
  XNOR U10808 ( .A(n43454), .B(n43232), .Z(n43234) );
  XNOR U10809 ( .A(n43235), .B(n43007), .Z(n43009) );
  XNOR U10810 ( .A(n43010), .B(n42776), .Z(n42778) );
  XNOR U10811 ( .A(n42779), .B(n42539), .Z(n42541) );
  XNOR U10812 ( .A(n42542), .B(n42296), .Z(n42298) );
  XNOR U10813 ( .A(n42299), .B(n42047), .Z(n42049) );
  XNOR U10814 ( .A(n42050), .B(n41792), .Z(n41794) );
  XNOR U10815 ( .A(n41795), .B(n41531), .Z(n41533) );
  XNOR U10816 ( .A(n41534), .B(n41264), .Z(n41266) );
  XNOR U10817 ( .A(n41267), .B(n40991), .Z(n40993) );
  XNOR U10818 ( .A(n40994), .B(n40712), .Z(n40714) );
  XNOR U10819 ( .A(n40715), .B(n40427), .Z(n40429) );
  XNOR U10820 ( .A(n40430), .B(n40136), .Z(n40138) );
  XNOR U10821 ( .A(n40139), .B(n39839), .Z(n39841) );
  XNOR U10822 ( .A(n39842), .B(n39536), .Z(n39538) );
  XNOR U10823 ( .A(n39539), .B(n39227), .Z(n39229) );
  XNOR U10824 ( .A(n39230), .B(n38912), .Z(n38914) );
  XNOR U10825 ( .A(n38915), .B(n38591), .Z(n38593) );
  XNOR U10826 ( .A(n38594), .B(n38264), .Z(n38266) );
  XNOR U10827 ( .A(n38267), .B(n37931), .Z(n37933) );
  XNOR U10828 ( .A(n37934), .B(n37592), .Z(n37594) );
  XNOR U10829 ( .A(n37595), .B(n37247), .Z(n37249) );
  XNOR U10830 ( .A(n37250), .B(n36896), .Z(n36898) );
  XNOR U10831 ( .A(n36899), .B(n36539), .Z(n36541) );
  XNOR U10832 ( .A(n36542), .B(n36176), .Z(n36178) );
  XNOR U10833 ( .A(n36179), .B(n35807), .Z(n35809) );
  XNOR U10834 ( .A(n35810), .B(n35432), .Z(n35434) );
  XNOR U10835 ( .A(n35435), .B(n35051), .Z(n35053) );
  XNOR U10836 ( .A(n35054), .B(n34664), .Z(n34666) );
  XNOR U10837 ( .A(n34667), .B(n34271), .Z(n34273) );
  XNOR U10838 ( .A(n34274), .B(n33872), .Z(n33874) );
  XNOR U10839 ( .A(n33875), .B(n33467), .Z(n33469) );
  XNOR U10840 ( .A(n33470), .B(n33056), .Z(n33058) );
  XNOR U10841 ( .A(n33059), .B(n32639), .Z(n32641) );
  XNOR U10842 ( .A(n32642), .B(n32216), .Z(n32218) );
  XNOR U10843 ( .A(n32219), .B(n31787), .Z(n31789) );
  XNOR U10844 ( .A(n31790), .B(n31352), .Z(n31354) );
  XNOR U10845 ( .A(n31355), .B(n30911), .Z(n30913) );
  XNOR U10846 ( .A(n30914), .B(n30464), .Z(n30466) );
  XNOR U10847 ( .A(n30467), .B(n30011), .Z(n30013) );
  XNOR U10848 ( .A(n30014), .B(n29552), .Z(n29554) );
  XNOR U10849 ( .A(n29555), .B(n29087), .Z(n29089) );
  XNOR U10850 ( .A(n29090), .B(n28616), .Z(n28618) );
  XNOR U10851 ( .A(n28619), .B(n28139), .Z(n28141) );
  XNOR U10852 ( .A(n28142), .B(n27656), .Z(n27658) );
  XNOR U10853 ( .A(n27659), .B(n27167), .Z(n27169) );
  XNOR U10854 ( .A(n27170), .B(n26670), .Z(n26672) );
  XNOR U10855 ( .A(n26673), .B(n26169), .Z(n26171) );
  XNOR U10856 ( .A(n26172), .B(n25661), .Z(n25663) );
  XNOR U10857 ( .A(n25664), .B(n25147), .Z(n25149) );
  XNOR U10858 ( .A(n25150), .B(n24624), .Z(n24626) );
  XNOR U10859 ( .A(n24627), .B(n24099), .Z(n24101) );
  XNOR U10860 ( .A(n24102), .B(n23568), .Z(n23570) );
  XNOR U10861 ( .A(n23571), .B(n23030), .Z(n23032) );
  XNOR U10862 ( .A(n23033), .B(n22486), .Z(n22488) );
  XNOR U10863 ( .A(n22489), .B(n21937), .Z(n21939) );
  XNOR U10864 ( .A(n21940), .B(n21382), .Z(n21384) );
  XNOR U10865 ( .A(n21385), .B(n20820), .Z(n20822) );
  XNOR U10866 ( .A(n20823), .B(n20253), .Z(n20255) );
  XNOR U10867 ( .A(n20256), .B(n19680), .Z(n19682) );
  XNOR U10868 ( .A(n19683), .B(n19101), .Z(n19103) );
  XOR U10869 ( .A(n18409), .B(n18655), .Z(n18413) );
  XOR U10870 ( .A(n17219), .B(n17426), .Z(n17223) );
  XOR U10871 ( .A(n16005), .B(n16212), .Z(n16009) );
  XOR U10872 ( .A(n14767), .B(n14974), .Z(n14771) );
  XOR U10873 ( .A(n13500), .B(n13713), .Z(n13504) );
  XOR U10874 ( .A(n12192), .B(n12431), .Z(n12196) );
  XOR U10875 ( .A(n10862), .B(n11123), .Z(n10866) );
  XOR U10876 ( .A(n11485), .B(n11788), .Z(n11489) );
  XOR U10877 ( .A(n10143), .B(n10470), .Z(n10147) );
  XOR U10878 ( .A(n8777), .B(n9128), .Z(n8781) );
  XOR U10879 ( .A(n9418), .B(n9811), .Z(n9422) );
  XOR U10880 ( .A(n8040), .B(n8457), .Z(n8044) );
  XOR U10881 ( .A(n6638), .B(n7079), .Z(n6642) );
  XOR U10882 ( .A(n7297), .B(n7780), .Z(n7301) );
  XOR U10883 ( .A(n5883), .B(n6390), .Z(n5887) );
  XOR U10884 ( .A(n4443), .B(n4974), .Z(n4447) );
  XOR U10885 ( .A(n5120), .B(n5695), .Z(n5124) );
  XOR U10886 ( .A(n3670), .B(n4267), .Z(n3674) );
  XOR U10887 ( .A(n2196), .B(n2817), .Z(n2200) );
  XOR U10888 ( .A(n2891), .B(n3554), .Z(n2895) );
  XOR U10889 ( .A(n1405), .B(n2092), .Z(n1409) );
  XOR U10890 ( .A(n1385), .B(n2096), .Z(n1389) );
  XOR U10891 ( .A(n12217), .B(n12426), .Z(n12221) );
  XOR U10892 ( .A(n2921), .B(n3548), .Z(n2925) );
  XOR U10893 ( .A(n1435), .B(n2086), .Z(n1439) );
  XOR U10894 ( .A(n5150), .B(n5689), .Z(n5154) );
  XOR U10895 ( .A(n3700), .B(n4261), .Z(n3704) );
  XOR U10896 ( .A(n2226), .B(n2811), .Z(n2230) );
  XOR U10897 ( .A(n7327), .B(n7774), .Z(n7331) );
  XOR U10898 ( .A(n5913), .B(n6384), .Z(n5917) );
  XOR U10899 ( .A(n4473), .B(n4968), .Z(n4477) );
  XOR U10900 ( .A(n9448), .B(n9805), .Z(n9452) );
  XOR U10901 ( .A(n8070), .B(n8451), .Z(n8074) );
  XOR U10902 ( .A(n6668), .B(n7073), .Z(n6672) );
  XOR U10903 ( .A(n11515), .B(n11782), .Z(n11519) );
  XOR U10904 ( .A(n10173), .B(n10464), .Z(n10177) );
  XOR U10905 ( .A(n8807), .B(n9122), .Z(n8811) );
  XOR U10906 ( .A(n10892), .B(n11117), .Z(n10896) );
  XNOR U10907 ( .A(n44474), .B(n44282), .Z(n44284) );
  XNOR U10908 ( .A(n44285), .B(n44087), .Z(n44089) );
  XNOR U10909 ( .A(n44090), .B(n43886), .Z(n43888) );
  XNOR U10910 ( .A(n43889), .B(n43679), .Z(n43681) );
  XNOR U10911 ( .A(n43682), .B(n43466), .Z(n43468) );
  XNOR U10912 ( .A(n43469), .B(n43247), .Z(n43249) );
  XNOR U10913 ( .A(n43250), .B(n43022), .Z(n43024) );
  XNOR U10914 ( .A(n43025), .B(n42791), .Z(n42793) );
  XNOR U10915 ( .A(n42794), .B(n42554), .Z(n42556) );
  XNOR U10916 ( .A(n42557), .B(n42311), .Z(n42313) );
  XNOR U10917 ( .A(n42314), .B(n42062), .Z(n42064) );
  XNOR U10918 ( .A(n42065), .B(n41807), .Z(n41809) );
  XNOR U10919 ( .A(n41810), .B(n41546), .Z(n41548) );
  XNOR U10920 ( .A(n41549), .B(n41279), .Z(n41281) );
  XNOR U10921 ( .A(n41282), .B(n41006), .Z(n41008) );
  XNOR U10922 ( .A(n41009), .B(n40727), .Z(n40729) );
  XNOR U10923 ( .A(n40730), .B(n40442), .Z(n40444) );
  XNOR U10924 ( .A(n40445), .B(n40151), .Z(n40153) );
  XNOR U10925 ( .A(n40154), .B(n39854), .Z(n39856) );
  XNOR U10926 ( .A(n39857), .B(n39551), .Z(n39553) );
  XNOR U10927 ( .A(n39554), .B(n39242), .Z(n39244) );
  XNOR U10928 ( .A(n39245), .B(n38927), .Z(n38929) );
  XNOR U10929 ( .A(n38930), .B(n38606), .Z(n38608) );
  XNOR U10930 ( .A(n38609), .B(n38279), .Z(n38281) );
  XNOR U10931 ( .A(n38282), .B(n37946), .Z(n37948) );
  XNOR U10932 ( .A(n37949), .B(n37607), .Z(n37609) );
  XNOR U10933 ( .A(n37610), .B(n37262), .Z(n37264) );
  XNOR U10934 ( .A(n37265), .B(n36911), .Z(n36913) );
  XNOR U10935 ( .A(n36914), .B(n36554), .Z(n36556) );
  XNOR U10936 ( .A(n36557), .B(n36191), .Z(n36193) );
  XNOR U10937 ( .A(n36194), .B(n35822), .Z(n35824) );
  XNOR U10938 ( .A(n35825), .B(n35447), .Z(n35449) );
  XNOR U10939 ( .A(n35450), .B(n35066), .Z(n35068) );
  XNOR U10940 ( .A(n35069), .B(n34679), .Z(n34681) );
  XNOR U10941 ( .A(n34682), .B(n34286), .Z(n34288) );
  XNOR U10942 ( .A(n34289), .B(n33887), .Z(n33889) );
  XNOR U10943 ( .A(n33890), .B(n33482), .Z(n33484) );
  XNOR U10944 ( .A(n33485), .B(n33071), .Z(n33073) );
  XNOR U10945 ( .A(n33074), .B(n32654), .Z(n32656) );
  XNOR U10946 ( .A(n32657), .B(n32231), .Z(n32233) );
  XNOR U10947 ( .A(n32234), .B(n31802), .Z(n31804) );
  XNOR U10948 ( .A(n31805), .B(n31367), .Z(n31369) );
  XNOR U10949 ( .A(n31370), .B(n30926), .Z(n30928) );
  XNOR U10950 ( .A(n30929), .B(n30479), .Z(n30481) );
  XNOR U10951 ( .A(n30482), .B(n30026), .Z(n30028) );
  XNOR U10952 ( .A(n30029), .B(n29567), .Z(n29569) );
  XNOR U10953 ( .A(n29570), .B(n29102), .Z(n29104) );
  XNOR U10954 ( .A(n29105), .B(n28631), .Z(n28633) );
  XNOR U10955 ( .A(n28634), .B(n28154), .Z(n28156) );
  XNOR U10956 ( .A(n28157), .B(n27671), .Z(n27673) );
  XNOR U10957 ( .A(n27674), .B(n27182), .Z(n27184) );
  XNOR U10958 ( .A(n27185), .B(n26685), .Z(n26687) );
  XNOR U10959 ( .A(n26688), .B(n26184), .Z(n26186) );
  XNOR U10960 ( .A(n26187), .B(n25676), .Z(n25678) );
  XNOR U10961 ( .A(n25679), .B(n25162), .Z(n25164) );
  XNOR U10962 ( .A(n25165), .B(n24639), .Z(n24641) );
  XNOR U10963 ( .A(n24642), .B(n24114), .Z(n24116) );
  XNOR U10964 ( .A(n24117), .B(n23583), .Z(n23585) );
  XNOR U10965 ( .A(n23586), .B(n23045), .Z(n23047) );
  XNOR U10966 ( .A(n23048), .B(n22501), .Z(n22503) );
  XNOR U10967 ( .A(n22504), .B(n21952), .Z(n21954) );
  XNOR U10968 ( .A(n21955), .B(n21397), .Z(n21399) );
  XNOR U10969 ( .A(n21400), .B(n20835), .Z(n20837) );
  XNOR U10970 ( .A(n20838), .B(n20268), .Z(n20270) );
  XNOR U10971 ( .A(n20271), .B(n19695), .Z(n19697) );
  XNOR U10972 ( .A(n19698), .B(n19116), .Z(n19118) );
  XOR U10973 ( .A(n17832), .B(n18021), .Z(n17836) );
  XOR U10974 ( .A(n16630), .B(n16819), .Z(n16634) );
  XOR U10975 ( .A(n15404), .B(n15593), .Z(n15408) );
  XOR U10976 ( .A(n14154), .B(n14343), .Z(n14158) );
  XOR U10977 ( .A(n12880), .B(n13069), .Z(n12884) );
  XOR U10978 ( .A(n10922), .B(n11111), .Z(n10926) );
  XOR U10979 ( .A(n11545), .B(n11776), .Z(n11549) );
  XOR U10980 ( .A(n10203), .B(n10458), .Z(n10207) );
  XOR U10981 ( .A(n8837), .B(n9116), .Z(n8841) );
  XOR U10982 ( .A(n9478), .B(n9799), .Z(n9482) );
  XOR U10983 ( .A(n8100), .B(n8445), .Z(n8104) );
  XOR U10984 ( .A(n6698), .B(n7067), .Z(n6702) );
  XOR U10985 ( .A(n7357), .B(n7768), .Z(n7361) );
  XOR U10986 ( .A(n5943), .B(n6378), .Z(n5947) );
  XOR U10987 ( .A(n4503), .B(n4962), .Z(n4507) );
  XOR U10988 ( .A(n5180), .B(n5683), .Z(n5184) );
  XOR U10989 ( .A(n3730), .B(n4255), .Z(n3734) );
  XOR U10990 ( .A(n2256), .B(n2805), .Z(n2260) );
  XOR U10991 ( .A(n2951), .B(n3542), .Z(n2955) );
  XOR U10992 ( .A(n1465), .B(n2080), .Z(n1469) );
  XOR U10993 ( .A(n703), .B(n1322), .Z(n713) );
  XOR U10994 ( .A(n717), .B(n1304), .Z(n727) );
  XOR U10995 ( .A(n2981), .B(n3536), .Z(n2985) );
  XOR U10996 ( .A(n1495), .B(n2074), .Z(n1499) );
  XOR U10997 ( .A(n5210), .B(n5677), .Z(n5214) );
  XOR U10998 ( .A(n3760), .B(n4249), .Z(n3764) );
  XOR U10999 ( .A(n2286), .B(n2799), .Z(n2290) );
  XOR U11000 ( .A(n7387), .B(n7762), .Z(n7391) );
  XOR U11001 ( .A(n5973), .B(n6372), .Z(n5977) );
  XOR U11002 ( .A(n4533), .B(n4956), .Z(n4537) );
  XOR U11003 ( .A(n9508), .B(n9793), .Z(n9512) );
  XOR U11004 ( .A(n8130), .B(n8439), .Z(n8134) );
  XOR U11005 ( .A(n6728), .B(n7061), .Z(n6732) );
  XOR U11006 ( .A(n11575), .B(n11770), .Z(n11579) );
  XOR U11007 ( .A(n10233), .B(n10452), .Z(n10237) );
  XOR U11008 ( .A(n8867), .B(n9110), .Z(n8871) );
  XNOR U11009 ( .A(n45020), .B(n44846), .Z(n44848) );
  XNOR U11010 ( .A(n44849), .B(n44669), .Z(n44671) );
  XNOR U11011 ( .A(n44672), .B(n44486), .Z(n44488) );
  XNOR U11012 ( .A(n44489), .B(n44297), .Z(n44299) );
  XNOR U11013 ( .A(n44300), .B(n44102), .Z(n44104) );
  XNOR U11014 ( .A(n44105), .B(n43901), .Z(n43903) );
  XNOR U11015 ( .A(n43904), .B(n43694), .Z(n43696) );
  XNOR U11016 ( .A(n43697), .B(n43481), .Z(n43483) );
  XNOR U11017 ( .A(n43484), .B(n43262), .Z(n43264) );
  XNOR U11018 ( .A(n43265), .B(n43037), .Z(n43039) );
  XNOR U11019 ( .A(n43040), .B(n42806), .Z(n42808) );
  XNOR U11020 ( .A(n42809), .B(n42569), .Z(n42571) );
  XNOR U11021 ( .A(n42572), .B(n42326), .Z(n42328) );
  XNOR U11022 ( .A(n42329), .B(n42077), .Z(n42079) );
  XNOR U11023 ( .A(n42080), .B(n41822), .Z(n41824) );
  XNOR U11024 ( .A(n41825), .B(n41561), .Z(n41563) );
  XNOR U11025 ( .A(n41564), .B(n41294), .Z(n41296) );
  XNOR U11026 ( .A(n41297), .B(n41021), .Z(n41023) );
  XNOR U11027 ( .A(n41024), .B(n40742), .Z(n40744) );
  XNOR U11028 ( .A(n40745), .B(n40457), .Z(n40459) );
  XNOR U11029 ( .A(n40460), .B(n40166), .Z(n40168) );
  XNOR U11030 ( .A(n40169), .B(n39869), .Z(n39871) );
  XNOR U11031 ( .A(n39872), .B(n39566), .Z(n39568) );
  XNOR U11032 ( .A(n39569), .B(n39257), .Z(n39259) );
  XNOR U11033 ( .A(n39260), .B(n38942), .Z(n38944) );
  XNOR U11034 ( .A(n38945), .B(n38621), .Z(n38623) );
  XNOR U11035 ( .A(n38624), .B(n38294), .Z(n38296) );
  XNOR U11036 ( .A(n38297), .B(n37961), .Z(n37963) );
  XNOR U11037 ( .A(n37964), .B(n37622), .Z(n37624) );
  XNOR U11038 ( .A(n37625), .B(n37277), .Z(n37279) );
  XNOR U11039 ( .A(n37280), .B(n36926), .Z(n36928) );
  XNOR U11040 ( .A(n36929), .B(n36569), .Z(n36571) );
  XNOR U11041 ( .A(n36572), .B(n36206), .Z(n36208) );
  XNOR U11042 ( .A(n36209), .B(n35837), .Z(n35839) );
  XNOR U11043 ( .A(n35840), .B(n35462), .Z(n35464) );
  XNOR U11044 ( .A(n35465), .B(n35081), .Z(n35083) );
  XNOR U11045 ( .A(n35084), .B(n34694), .Z(n34696) );
  XNOR U11046 ( .A(n34697), .B(n34301), .Z(n34303) );
  XNOR U11047 ( .A(n34304), .B(n33902), .Z(n33904) );
  XNOR U11048 ( .A(n33905), .B(n33497), .Z(n33499) );
  XNOR U11049 ( .A(n33500), .B(n33086), .Z(n33088) );
  XNOR U11050 ( .A(n33089), .B(n32669), .Z(n32671) );
  XNOR U11051 ( .A(n32672), .B(n32246), .Z(n32248) );
  XNOR U11052 ( .A(n32249), .B(n31817), .Z(n31819) );
  XNOR U11053 ( .A(n31820), .B(n31382), .Z(n31384) );
  XNOR U11054 ( .A(n31385), .B(n30941), .Z(n30943) );
  XNOR U11055 ( .A(n30944), .B(n30494), .Z(n30496) );
  XNOR U11056 ( .A(n30497), .B(n30041), .Z(n30043) );
  XNOR U11057 ( .A(n30044), .B(n29582), .Z(n29584) );
  XNOR U11058 ( .A(n29585), .B(n29117), .Z(n29119) );
  XNOR U11059 ( .A(n29120), .B(n28646), .Z(n28648) );
  XNOR U11060 ( .A(n28649), .B(n28169), .Z(n28171) );
  XNOR U11061 ( .A(n28172), .B(n27686), .Z(n27688) );
  XNOR U11062 ( .A(n27689), .B(n27197), .Z(n27199) );
  XNOR U11063 ( .A(n27200), .B(n26700), .Z(n26702) );
  XNOR U11064 ( .A(n26703), .B(n26199), .Z(n26201) );
  XNOR U11065 ( .A(n26202), .B(n25691), .Z(n25693) );
  XNOR U11066 ( .A(n25694), .B(n25177), .Z(n25179) );
  XNOR U11067 ( .A(n25180), .B(n24654), .Z(n24656) );
  XNOR U11068 ( .A(n24657), .B(n24129), .Z(n24131) );
  XNOR U11069 ( .A(n24132), .B(n23598), .Z(n23600) );
  XNOR U11070 ( .A(n23601), .B(n23060), .Z(n23062) );
  XNOR U11071 ( .A(n23063), .B(n22516), .Z(n22518) );
  XNOR U11072 ( .A(n22519), .B(n21967), .Z(n21969) );
  XNOR U11073 ( .A(n21970), .B(n21412), .Z(n21414) );
  XNOR U11074 ( .A(n21415), .B(n20850), .Z(n20852) );
  XNOR U11075 ( .A(n20853), .B(n20283), .Z(n20285) );
  XNOR U11076 ( .A(n20286), .B(n19710), .Z(n19712) );
  XNOR U11077 ( .A(n19713), .B(n19131), .Z(n19133) );
  XOR U11078 ( .A(n18439), .B(n18643), .Z(n18443) );
  XOR U11079 ( .A(n17249), .B(n17420), .Z(n17253) );
  XOR U11080 ( .A(n16035), .B(n16206), .Z(n16039) );
  XOR U11081 ( .A(n14797), .B(n14968), .Z(n14801) );
  XOR U11082 ( .A(n13535), .B(n13706), .Z(n13539) );
  XOR U11083 ( .A(n12247), .B(n12420), .Z(n12251) );
  XOR U11084 ( .A(n10263), .B(n10446), .Z(n10267) );
  XOR U11085 ( .A(n8897), .B(n9104), .Z(n8901) );
  XOR U11086 ( .A(n9538), .B(n9787), .Z(n9542) );
  XOR U11087 ( .A(n8160), .B(n8433), .Z(n8164) );
  XOR U11088 ( .A(n6758), .B(n7055), .Z(n6762) );
  XOR U11089 ( .A(n7417), .B(n7756), .Z(n7421) );
  XOR U11090 ( .A(n6003), .B(n6366), .Z(n6007) );
  XOR U11091 ( .A(n4563), .B(n4950), .Z(n4567) );
  XOR U11092 ( .A(n5240), .B(n5671), .Z(n5244) );
  XOR U11093 ( .A(n3790), .B(n4243), .Z(n3794) );
  XOR U11094 ( .A(n2316), .B(n2793), .Z(n2320) );
  XOR U11095 ( .A(n3011), .B(n3530), .Z(n3015) );
  XOR U11096 ( .A(n1525), .B(n2068), .Z(n1529) );
  XOR U11097 ( .A(n731), .B(n1286), .Z(n741) );
  XOR U11098 ( .A(n745), .B(n1268), .Z(n755) );
  XOR U11099 ( .A(n3041), .B(n3524), .Z(n3045) );
  XOR U11100 ( .A(n1555), .B(n2062), .Z(n1559) );
  XOR U11101 ( .A(n5270), .B(n5665), .Z(n5274) );
  XOR U11102 ( .A(n3820), .B(n4237), .Z(n3824) );
  XOR U11103 ( .A(n2346), .B(n2787), .Z(n2350) );
  XOR U11104 ( .A(n7447), .B(n7750), .Z(n7451) );
  XOR U11105 ( .A(n6033), .B(n6360), .Z(n6037) );
  XOR U11106 ( .A(n4593), .B(n4944), .Z(n4597) );
  XOR U11107 ( .A(n9568), .B(n9781), .Z(n9572) );
  XOR U11108 ( .A(n8190), .B(n8427), .Z(n8194) );
  XOR U11109 ( .A(n6788), .B(n7049), .Z(n6792) );
  XOR U11110 ( .A(n8927), .B(n9098), .Z(n8931) );
  XNOR U11111 ( .A(n45512), .B(n45356), .Z(n45358) );
  XNOR U11112 ( .A(n45359), .B(n45197), .Z(n45199) );
  XNOR U11113 ( .A(n45200), .B(n45032), .Z(n45034) );
  XNOR U11114 ( .A(n45035), .B(n44861), .Z(n44863) );
  XNOR U11115 ( .A(n44864), .B(n44684), .Z(n44686) );
  XNOR U11116 ( .A(n44687), .B(n44501), .Z(n44503) );
  XNOR U11117 ( .A(n44504), .B(n44312), .Z(n44314) );
  XNOR U11118 ( .A(n44315), .B(n44117), .Z(n44119) );
  XNOR U11119 ( .A(n44120), .B(n43916), .Z(n43918) );
  XNOR U11120 ( .A(n43919), .B(n43709), .Z(n43711) );
  XNOR U11121 ( .A(n43712), .B(n43496), .Z(n43498) );
  XNOR U11122 ( .A(n43499), .B(n43277), .Z(n43279) );
  XNOR U11123 ( .A(n43280), .B(n43052), .Z(n43054) );
  XNOR U11124 ( .A(n43055), .B(n42821), .Z(n42823) );
  XNOR U11125 ( .A(n42824), .B(n42584), .Z(n42586) );
  XNOR U11126 ( .A(n42587), .B(n42341), .Z(n42343) );
  XNOR U11127 ( .A(n42344), .B(n42092), .Z(n42094) );
  XNOR U11128 ( .A(n42095), .B(n41837), .Z(n41839) );
  XNOR U11129 ( .A(n41840), .B(n41576), .Z(n41578) );
  XNOR U11130 ( .A(n41579), .B(n41309), .Z(n41311) );
  XNOR U11131 ( .A(n41312), .B(n41036), .Z(n41038) );
  XNOR U11132 ( .A(n41039), .B(n40757), .Z(n40759) );
  XNOR U11133 ( .A(n40760), .B(n40472), .Z(n40474) );
  XNOR U11134 ( .A(n40475), .B(n40181), .Z(n40183) );
  XNOR U11135 ( .A(n40184), .B(n39884), .Z(n39886) );
  XNOR U11136 ( .A(n39887), .B(n39581), .Z(n39583) );
  XNOR U11137 ( .A(n39584), .B(n39272), .Z(n39274) );
  XNOR U11138 ( .A(n39275), .B(n38957), .Z(n38959) );
  XNOR U11139 ( .A(n38960), .B(n38636), .Z(n38638) );
  XNOR U11140 ( .A(n38639), .B(n38309), .Z(n38311) );
  XNOR U11141 ( .A(n38312), .B(n37976), .Z(n37978) );
  XNOR U11142 ( .A(n37979), .B(n37637), .Z(n37639) );
  XNOR U11143 ( .A(n37640), .B(n37292), .Z(n37294) );
  XNOR U11144 ( .A(n37295), .B(n36941), .Z(n36943) );
  XNOR U11145 ( .A(n36944), .B(n36584), .Z(n36586) );
  XNOR U11146 ( .A(n36587), .B(n36221), .Z(n36223) );
  XNOR U11147 ( .A(n36224), .B(n35852), .Z(n35854) );
  XNOR U11148 ( .A(n35855), .B(n35477), .Z(n35479) );
  XNOR U11149 ( .A(n35480), .B(n35096), .Z(n35098) );
  XNOR U11150 ( .A(n35099), .B(n34709), .Z(n34711) );
  XNOR U11151 ( .A(n34712), .B(n34316), .Z(n34318) );
  XNOR U11152 ( .A(n34319), .B(n33917), .Z(n33919) );
  XNOR U11153 ( .A(n33920), .B(n33512), .Z(n33514) );
  XNOR U11154 ( .A(n33515), .B(n33101), .Z(n33103) );
  XNOR U11155 ( .A(n33104), .B(n32684), .Z(n32686) );
  XNOR U11156 ( .A(n32687), .B(n32261), .Z(n32263) );
  XNOR U11157 ( .A(n32264), .B(n31832), .Z(n31834) );
  XNOR U11158 ( .A(n31835), .B(n31397), .Z(n31399) );
  XNOR U11159 ( .A(n31400), .B(n30956), .Z(n30958) );
  XNOR U11160 ( .A(n30959), .B(n30509), .Z(n30511) );
  XNOR U11161 ( .A(n30512), .B(n30056), .Z(n30058) );
  XNOR U11162 ( .A(n30059), .B(n29597), .Z(n29599) );
  XNOR U11163 ( .A(n29600), .B(n29132), .Z(n29134) );
  XNOR U11164 ( .A(n29135), .B(n28661), .Z(n28663) );
  XNOR U11165 ( .A(n28664), .B(n28184), .Z(n28186) );
  XNOR U11166 ( .A(n28187), .B(n27701), .Z(n27703) );
  XNOR U11167 ( .A(n27704), .B(n27212), .Z(n27214) );
  XNOR U11168 ( .A(n27215), .B(n26715), .Z(n26717) );
  XNOR U11169 ( .A(n26718), .B(n26214), .Z(n26216) );
  XNOR U11170 ( .A(n26217), .B(n25706), .Z(n25708) );
  XNOR U11171 ( .A(n25709), .B(n25192), .Z(n25194) );
  XNOR U11172 ( .A(n25195), .B(n24669), .Z(n24671) );
  XNOR U11173 ( .A(n24672), .B(n24144), .Z(n24146) );
  XNOR U11174 ( .A(n24147), .B(n23613), .Z(n23615) );
  XNOR U11175 ( .A(n23616), .B(n23075), .Z(n23077) );
  XNOR U11176 ( .A(n23078), .B(n22531), .Z(n22533) );
  XNOR U11177 ( .A(n22534), .B(n21982), .Z(n21984) );
  XNOR U11178 ( .A(n21985), .B(n21427), .Z(n21429) );
  XNOR U11179 ( .A(n21430), .B(n20865), .Z(n20867) );
  XNOR U11180 ( .A(n20868), .B(n20298), .Z(n20300) );
  XNOR U11181 ( .A(n20301), .B(n19725), .Z(n19727) );
  XNOR U11182 ( .A(n19728), .B(n19146), .Z(n19148) );
  XOR U11183 ( .A(n17862), .B(n18015), .Z(n17866) );
  XOR U11184 ( .A(n16660), .B(n16813), .Z(n16664) );
  XOR U11185 ( .A(n15434), .B(n15587), .Z(n15438) );
  XOR U11186 ( .A(n14184), .B(n14337), .Z(n14188) );
  XOR U11187 ( .A(n12910), .B(n13063), .Z(n12914) );
  XOR U11188 ( .A(n11610), .B(n11763), .Z(n11614) );
  XOR U11189 ( .A(n10288), .B(n10441), .Z(n10292) );
  XOR U11190 ( .A(n9598), .B(n9775), .Z(n9602) );
  XOR U11191 ( .A(n8220), .B(n8421), .Z(n8224) );
  XOR U11192 ( .A(n6818), .B(n7043), .Z(n6822) );
  XOR U11193 ( .A(n7477), .B(n7744), .Z(n7481) );
  XOR U11194 ( .A(n6063), .B(n6354), .Z(n6067) );
  XOR U11195 ( .A(n4623), .B(n4938), .Z(n4627) );
  XOR U11196 ( .A(n5300), .B(n5659), .Z(n5304) );
  XOR U11197 ( .A(n3850), .B(n4231), .Z(n3854) );
  XOR U11198 ( .A(n2376), .B(n2781), .Z(n2380) );
  XOR U11199 ( .A(n3071), .B(n3518), .Z(n3075) );
  XOR U11200 ( .A(n1585), .B(n2056), .Z(n1589) );
  XOR U11201 ( .A(n759), .B(n1250), .Z(n769) );
  XOR U11202 ( .A(n773), .B(n1232), .Z(n783) );
  XOR U11203 ( .A(n3101), .B(n3512), .Z(n3105) );
  XOR U11204 ( .A(n1615), .B(n2050), .Z(n1619) );
  XOR U11205 ( .A(n5330), .B(n5653), .Z(n5334) );
  XOR U11206 ( .A(n3880), .B(n4225), .Z(n3884) );
  XOR U11207 ( .A(n2406), .B(n2775), .Z(n2410) );
  XOR U11208 ( .A(n7507), .B(n7738), .Z(n7511) );
  XOR U11209 ( .A(n6093), .B(n6348), .Z(n6097) );
  XOR U11210 ( .A(n4653), .B(n4932), .Z(n4657) );
  XOR U11211 ( .A(n9628), .B(n9769), .Z(n9632) );
  XOR U11212 ( .A(n8250), .B(n8415), .Z(n8254) );
  XOR U11213 ( .A(n6848), .B(n7037), .Z(n6852) );
  XNOR U11214 ( .A(n45950), .B(n45812), .Z(n45814) );
  XNOR U11215 ( .A(n45815), .B(n45671), .Z(n45673) );
  XNOR U11216 ( .A(n45674), .B(n45524), .Z(n45526) );
  XNOR U11217 ( .A(n45527), .B(n45371), .Z(n45373) );
  XNOR U11218 ( .A(n45374), .B(n45212), .Z(n45214) );
  XNOR U11219 ( .A(n45215), .B(n45047), .Z(n45049) );
  XNOR U11220 ( .A(n45050), .B(n44876), .Z(n44878) );
  XNOR U11221 ( .A(n44879), .B(n44699), .Z(n44701) );
  XNOR U11222 ( .A(n44702), .B(n44516), .Z(n44518) );
  XNOR U11223 ( .A(n44519), .B(n44327), .Z(n44329) );
  XNOR U11224 ( .A(n44330), .B(n44132), .Z(n44134) );
  XNOR U11225 ( .A(n44135), .B(n43931), .Z(n43933) );
  XNOR U11226 ( .A(n43934), .B(n43724), .Z(n43726) );
  XNOR U11227 ( .A(n43727), .B(n43511), .Z(n43513) );
  XNOR U11228 ( .A(n43514), .B(n43292), .Z(n43294) );
  XNOR U11229 ( .A(n43295), .B(n43067), .Z(n43069) );
  XNOR U11230 ( .A(n43070), .B(n42836), .Z(n42838) );
  XNOR U11231 ( .A(n42839), .B(n42599), .Z(n42601) );
  XNOR U11232 ( .A(n42602), .B(n42356), .Z(n42358) );
  XNOR U11233 ( .A(n42359), .B(n42107), .Z(n42109) );
  XNOR U11234 ( .A(n42110), .B(n41852), .Z(n41854) );
  XNOR U11235 ( .A(n41855), .B(n41591), .Z(n41593) );
  XNOR U11236 ( .A(n41594), .B(n41324), .Z(n41326) );
  XNOR U11237 ( .A(n41327), .B(n41051), .Z(n41053) );
  XNOR U11238 ( .A(n41054), .B(n40772), .Z(n40774) );
  XNOR U11239 ( .A(n40775), .B(n40487), .Z(n40489) );
  XNOR U11240 ( .A(n40490), .B(n40196), .Z(n40198) );
  XNOR U11241 ( .A(n40199), .B(n39899), .Z(n39901) );
  XNOR U11242 ( .A(n39902), .B(n39596), .Z(n39598) );
  XNOR U11243 ( .A(n39599), .B(n39287), .Z(n39289) );
  XNOR U11244 ( .A(n39290), .B(n38972), .Z(n38974) );
  XNOR U11245 ( .A(n38975), .B(n38651), .Z(n38653) );
  XNOR U11246 ( .A(n38654), .B(n38324), .Z(n38326) );
  XNOR U11247 ( .A(n38327), .B(n37991), .Z(n37993) );
  XNOR U11248 ( .A(n37994), .B(n37652), .Z(n37654) );
  XNOR U11249 ( .A(n37655), .B(n37307), .Z(n37309) );
  XNOR U11250 ( .A(n37310), .B(n36956), .Z(n36958) );
  XNOR U11251 ( .A(n36959), .B(n36599), .Z(n36601) );
  XNOR U11252 ( .A(n36602), .B(n36236), .Z(n36238) );
  XNOR U11253 ( .A(n36239), .B(n35867), .Z(n35869) );
  XNOR U11254 ( .A(n35870), .B(n35492), .Z(n35494) );
  XNOR U11255 ( .A(n35495), .B(n35111), .Z(n35113) );
  XNOR U11256 ( .A(n35114), .B(n34724), .Z(n34726) );
  XNOR U11257 ( .A(n34727), .B(n34331), .Z(n34333) );
  XNOR U11258 ( .A(n34334), .B(n33932), .Z(n33934) );
  XNOR U11259 ( .A(n33935), .B(n33527), .Z(n33529) );
  XNOR U11260 ( .A(n33530), .B(n33116), .Z(n33118) );
  XNOR U11261 ( .A(n33119), .B(n32699), .Z(n32701) );
  XNOR U11262 ( .A(n32702), .B(n32276), .Z(n32278) );
  XNOR U11263 ( .A(n32279), .B(n31847), .Z(n31849) );
  XNOR U11264 ( .A(n31850), .B(n31412), .Z(n31414) );
  XNOR U11265 ( .A(n31415), .B(n30971), .Z(n30973) );
  XNOR U11266 ( .A(n30974), .B(n30524), .Z(n30526) );
  XNOR U11267 ( .A(n30527), .B(n30071), .Z(n30073) );
  XNOR U11268 ( .A(n30074), .B(n29612), .Z(n29614) );
  XNOR U11269 ( .A(n29615), .B(n29147), .Z(n29149) );
  XNOR U11270 ( .A(n29150), .B(n28676), .Z(n28678) );
  XNOR U11271 ( .A(n28679), .B(n28199), .Z(n28201) );
  XNOR U11272 ( .A(n28202), .B(n27716), .Z(n27718) );
  XNOR U11273 ( .A(n27719), .B(n27227), .Z(n27229) );
  XNOR U11274 ( .A(n27230), .B(n26730), .Z(n26732) );
  XNOR U11275 ( .A(n26733), .B(n26229), .Z(n26231) );
  XNOR U11276 ( .A(n26232), .B(n25721), .Z(n25723) );
  XNOR U11277 ( .A(n25724), .B(n25207), .Z(n25209) );
  XNOR U11278 ( .A(n25210), .B(n24684), .Z(n24686) );
  XNOR U11279 ( .A(n24687), .B(n24159), .Z(n24161) );
  XNOR U11280 ( .A(n24162), .B(n23628), .Z(n23630) );
  XNOR U11281 ( .A(n23631), .B(n23090), .Z(n23092) );
  XNOR U11282 ( .A(n23093), .B(n22546), .Z(n22548) );
  XNOR U11283 ( .A(n22549), .B(n21997), .Z(n21999) );
  XNOR U11284 ( .A(n22000), .B(n21442), .Z(n21444) );
  XNOR U11285 ( .A(n21445), .B(n20880), .Z(n20882) );
  XNOR U11286 ( .A(n20883), .B(n20313), .Z(n20315) );
  XNOR U11287 ( .A(n20316), .B(n19740), .Z(n19742) );
  XNOR U11288 ( .A(n19743), .B(n19161), .Z(n19163) );
  XOR U11289 ( .A(n18469), .B(n18631), .Z(n18473) );
  XOR U11290 ( .A(n17279), .B(n17414), .Z(n17283) );
  XOR U11291 ( .A(n16065), .B(n16200), .Z(n16069) );
  XOR U11292 ( .A(n14827), .B(n14962), .Z(n14831) );
  XOR U11293 ( .A(n13565), .B(n13700), .Z(n13569) );
  XOR U11294 ( .A(n12277), .B(n12414), .Z(n12281) );
  XOR U11295 ( .A(n10967), .B(n11102), .Z(n10971) );
  XOR U11296 ( .A(n6878), .B(n7031), .Z(n6882) );
  XOR U11297 ( .A(n7537), .B(n7732), .Z(n7541) );
  XOR U11298 ( .A(n6123), .B(n6342), .Z(n6127) );
  XOR U11299 ( .A(n4683), .B(n4926), .Z(n4687) );
  XOR U11300 ( .A(n5360), .B(n5647), .Z(n5364) );
  XOR U11301 ( .A(n3910), .B(n4219), .Z(n3914) );
  XOR U11302 ( .A(n2436), .B(n2769), .Z(n2440) );
  XOR U11303 ( .A(n3131), .B(n3506), .Z(n3135) );
  XOR U11304 ( .A(n1645), .B(n2044), .Z(n1649) );
  XOR U11305 ( .A(n787), .B(n1214), .Z(n797) );
  XOR U11306 ( .A(n10313), .B(n10436), .Z(n10317) );
  XOR U11307 ( .A(n8967), .B(n9090), .Z(n8971) );
  XOR U11308 ( .A(n801), .B(n1196), .Z(n811) );
  XOR U11309 ( .A(n3161), .B(n3500), .Z(n3165) );
  XOR U11310 ( .A(n1675), .B(n2038), .Z(n1679) );
  XOR U11311 ( .A(n5390), .B(n5641), .Z(n5394) );
  XOR U11312 ( .A(n3940), .B(n4213), .Z(n3944) );
  XOR U11313 ( .A(n2466), .B(n2763), .Z(n2470) );
  XOR U11314 ( .A(n7567), .B(n7726), .Z(n7571) );
  XOR U11315 ( .A(n6153), .B(n6336), .Z(n6157) );
  XOR U11316 ( .A(n4713), .B(n4920), .Z(n4717) );
  XNOR U11317 ( .A(n46334), .B(n46214), .Z(n46216) );
  XNOR U11318 ( .A(n46217), .B(n46091), .Z(n46093) );
  XNOR U11319 ( .A(n46094), .B(n45962), .Z(n45964) );
  XNOR U11320 ( .A(n45965), .B(n45827), .Z(n45829) );
  XNOR U11321 ( .A(n45830), .B(n45686), .Z(n45688) );
  XNOR U11322 ( .A(n45689), .B(n45539), .Z(n45541) );
  XNOR U11323 ( .A(n45542), .B(n45386), .Z(n45388) );
  XNOR U11324 ( .A(n45389), .B(n45227), .Z(n45229) );
  XNOR U11325 ( .A(n45230), .B(n45062), .Z(n45064) );
  XNOR U11326 ( .A(n45065), .B(n44891), .Z(n44893) );
  XNOR U11327 ( .A(n44894), .B(n44714), .Z(n44716) );
  XNOR U11328 ( .A(n44717), .B(n44531), .Z(n44533) );
  XNOR U11329 ( .A(n44534), .B(n44342), .Z(n44344) );
  XNOR U11330 ( .A(n44345), .B(n44147), .Z(n44149) );
  XNOR U11331 ( .A(n44150), .B(n43946), .Z(n43948) );
  XNOR U11332 ( .A(n43949), .B(n43739), .Z(n43741) );
  XNOR U11333 ( .A(n43742), .B(n43526), .Z(n43528) );
  XNOR U11334 ( .A(n43529), .B(n43307), .Z(n43309) );
  XNOR U11335 ( .A(n43310), .B(n43082), .Z(n43084) );
  XNOR U11336 ( .A(n43085), .B(n42851), .Z(n42853) );
  XNOR U11337 ( .A(n42854), .B(n42614), .Z(n42616) );
  XNOR U11338 ( .A(n42617), .B(n42371), .Z(n42373) );
  XNOR U11339 ( .A(n42374), .B(n42122), .Z(n42124) );
  XNOR U11340 ( .A(n42125), .B(n41867), .Z(n41869) );
  XNOR U11341 ( .A(n41870), .B(n41606), .Z(n41608) );
  XNOR U11342 ( .A(n41609), .B(n41339), .Z(n41341) );
  XNOR U11343 ( .A(n41342), .B(n41066), .Z(n41068) );
  XNOR U11344 ( .A(n41069), .B(n40787), .Z(n40789) );
  XNOR U11345 ( .A(n40790), .B(n40502), .Z(n40504) );
  XNOR U11346 ( .A(n40505), .B(n40211), .Z(n40213) );
  XNOR U11347 ( .A(n40214), .B(n39914), .Z(n39916) );
  XNOR U11348 ( .A(n39917), .B(n39611), .Z(n39613) );
  XNOR U11349 ( .A(n39614), .B(n39302), .Z(n39304) );
  XNOR U11350 ( .A(n39305), .B(n38987), .Z(n38989) );
  XNOR U11351 ( .A(n38990), .B(n38666), .Z(n38668) );
  XNOR U11352 ( .A(n38669), .B(n38339), .Z(n38341) );
  XNOR U11353 ( .A(n38342), .B(n38006), .Z(n38008) );
  XNOR U11354 ( .A(n38009), .B(n37667), .Z(n37669) );
  XNOR U11355 ( .A(n37670), .B(n37322), .Z(n37324) );
  XNOR U11356 ( .A(n37325), .B(n36971), .Z(n36973) );
  XNOR U11357 ( .A(n36974), .B(n36614), .Z(n36616) );
  XNOR U11358 ( .A(n36617), .B(n36251), .Z(n36253) );
  XNOR U11359 ( .A(n36254), .B(n35882), .Z(n35884) );
  XNOR U11360 ( .A(n35885), .B(n35507), .Z(n35509) );
  XNOR U11361 ( .A(n35510), .B(n35126), .Z(n35128) );
  XNOR U11362 ( .A(n35129), .B(n34739), .Z(n34741) );
  XNOR U11363 ( .A(n34742), .B(n34346), .Z(n34348) );
  XNOR U11364 ( .A(n34349), .B(n33947), .Z(n33949) );
  XNOR U11365 ( .A(n33950), .B(n33542), .Z(n33544) );
  XNOR U11366 ( .A(n33545), .B(n33131), .Z(n33133) );
  XNOR U11367 ( .A(n33134), .B(n32714), .Z(n32716) );
  XNOR U11368 ( .A(n32717), .B(n32291), .Z(n32293) );
  XNOR U11369 ( .A(n32294), .B(n31862), .Z(n31864) );
  XNOR U11370 ( .A(n31865), .B(n31427), .Z(n31429) );
  XNOR U11371 ( .A(n31430), .B(n30986), .Z(n30988) );
  XNOR U11372 ( .A(n30989), .B(n30539), .Z(n30541) );
  XNOR U11373 ( .A(n30542), .B(n30086), .Z(n30088) );
  XNOR U11374 ( .A(n30089), .B(n29627), .Z(n29629) );
  XNOR U11375 ( .A(n29630), .B(n29162), .Z(n29164) );
  XNOR U11376 ( .A(n29165), .B(n28691), .Z(n28693) );
  XNOR U11377 ( .A(n28694), .B(n28214), .Z(n28216) );
  XNOR U11378 ( .A(n28217), .B(n27731), .Z(n27733) );
  XNOR U11379 ( .A(n27734), .B(n27242), .Z(n27244) );
  XNOR U11380 ( .A(n27245), .B(n26745), .Z(n26747) );
  XNOR U11381 ( .A(n26748), .B(n26244), .Z(n26246) );
  XNOR U11382 ( .A(n26247), .B(n25736), .Z(n25738) );
  XNOR U11383 ( .A(n25739), .B(n25222), .Z(n25224) );
  XNOR U11384 ( .A(n25225), .B(n24699), .Z(n24701) );
  XNOR U11385 ( .A(n24702), .B(n24174), .Z(n24176) );
  XNOR U11386 ( .A(n24177), .B(n23643), .Z(n23645) );
  XNOR U11387 ( .A(n23646), .B(n23105), .Z(n23107) );
  XNOR U11388 ( .A(n23108), .B(n22561), .Z(n22563) );
  XNOR U11389 ( .A(n22564), .B(n22012), .Z(n22014) );
  XNOR U11390 ( .A(n22015), .B(n21457), .Z(n21459) );
  XNOR U11391 ( .A(n21460), .B(n20895), .Z(n20897) );
  XNOR U11392 ( .A(n20898), .B(n20328), .Z(n20330) );
  XNOR U11393 ( .A(n20331), .B(n19755), .Z(n19757) );
  XNOR U11394 ( .A(n19758), .B(n19176), .Z(n19178) );
  XOR U11395 ( .A(n18484), .B(n18625), .Z(n18488) );
  XOR U11396 ( .A(n17294), .B(n17411), .Z(n17298) );
  XOR U11397 ( .A(n16080), .B(n16197), .Z(n16084) );
  XOR U11398 ( .A(n14842), .B(n14959), .Z(n14846) );
  XOR U11399 ( .A(n13580), .B(n13697), .Z(n13584) );
  XOR U11400 ( .A(n12292), .B(n12411), .Z(n12296) );
  XOR U11401 ( .A(n7597), .B(n7720), .Z(n7601) );
  XOR U11402 ( .A(n6183), .B(n6330), .Z(n6187) );
  XOR U11403 ( .A(n4743), .B(n4914), .Z(n4747) );
  XOR U11404 ( .A(n5420), .B(n5635), .Z(n5424) );
  XOR U11405 ( .A(n3970), .B(n4207), .Z(n3974) );
  XOR U11406 ( .A(n2496), .B(n2757), .Z(n2500) );
  XOR U11407 ( .A(n3191), .B(n3494), .Z(n3195) );
  XOR U11408 ( .A(n1705), .B(n2032), .Z(n1709) );
  XOR U11409 ( .A(n815), .B(n1178), .Z(n825) );
  XOR U11410 ( .A(n11650), .B(n11755), .Z(n11654) );
  XOR U11411 ( .A(n10328), .B(n10433), .Z(n10332) );
  XOR U11412 ( .A(n8982), .B(n9087), .Z(n8986) );
  XOR U11413 ( .A(n7612), .B(n7717), .Z(n7616) );
  XOR U11414 ( .A(n829), .B(n1160), .Z(n839) );
  XOR U11415 ( .A(n3221), .B(n3488), .Z(n3225) );
  XOR U11416 ( .A(n1735), .B(n2026), .Z(n1739) );
  XOR U11417 ( .A(n5450), .B(n5629), .Z(n5454) );
  XOR U11418 ( .A(n4000), .B(n4201), .Z(n4004) );
  XOR U11419 ( .A(n2526), .B(n2751), .Z(n2530) );
  XOR U11420 ( .A(n6213), .B(n6324), .Z(n6217) );
  XOR U11421 ( .A(n4773), .B(n4908), .Z(n4777) );
  XNOR U11422 ( .A(n46664), .B(n46562), .Z(n46564) );
  XNOR U11423 ( .A(n46565), .B(n46457), .Z(n46459) );
  XNOR U11424 ( .A(n46460), .B(n46346), .Z(n46348) );
  XNOR U11425 ( .A(n46349), .B(n46229), .Z(n46231) );
  XNOR U11426 ( .A(n46232), .B(n46106), .Z(n46108) );
  XNOR U11427 ( .A(n46109), .B(n45977), .Z(n45979) );
  XNOR U11428 ( .A(n45980), .B(n45842), .Z(n45844) );
  XNOR U11429 ( .A(n45845), .B(n45701), .Z(n45703) );
  XNOR U11430 ( .A(n45704), .B(n45554), .Z(n45556) );
  XNOR U11431 ( .A(n45557), .B(n45401), .Z(n45403) );
  XNOR U11432 ( .A(n45404), .B(n45242), .Z(n45244) );
  XNOR U11433 ( .A(n45245), .B(n45077), .Z(n45079) );
  XNOR U11434 ( .A(n45080), .B(n44906), .Z(n44908) );
  XNOR U11435 ( .A(n44909), .B(n44729), .Z(n44731) );
  XNOR U11436 ( .A(n44732), .B(n44546), .Z(n44548) );
  XNOR U11437 ( .A(n44549), .B(n44357), .Z(n44359) );
  XNOR U11438 ( .A(n44360), .B(n44162), .Z(n44164) );
  XNOR U11439 ( .A(n44165), .B(n43961), .Z(n43963) );
  XNOR U11440 ( .A(n43964), .B(n43754), .Z(n43756) );
  XNOR U11441 ( .A(n43757), .B(n43541), .Z(n43543) );
  XNOR U11442 ( .A(n43544), .B(n43322), .Z(n43324) );
  XNOR U11443 ( .A(n43325), .B(n43097), .Z(n43099) );
  XNOR U11444 ( .A(n43100), .B(n42866), .Z(n42868) );
  XNOR U11445 ( .A(n42869), .B(n42629), .Z(n42631) );
  XNOR U11446 ( .A(n42632), .B(n42386), .Z(n42388) );
  XNOR U11447 ( .A(n42389), .B(n42137), .Z(n42139) );
  XNOR U11448 ( .A(n42140), .B(n41882), .Z(n41884) );
  XNOR U11449 ( .A(n41885), .B(n41621), .Z(n41623) );
  XNOR U11450 ( .A(n41624), .B(n41354), .Z(n41356) );
  XNOR U11451 ( .A(n41357), .B(n41081), .Z(n41083) );
  XNOR U11452 ( .A(n41084), .B(n40802), .Z(n40804) );
  XNOR U11453 ( .A(n40805), .B(n40517), .Z(n40519) );
  XNOR U11454 ( .A(n40520), .B(n40226), .Z(n40228) );
  XNOR U11455 ( .A(n40229), .B(n39929), .Z(n39931) );
  XNOR U11456 ( .A(n39932), .B(n39626), .Z(n39628) );
  XNOR U11457 ( .A(n39629), .B(n39317), .Z(n39319) );
  XNOR U11458 ( .A(n39320), .B(n39002), .Z(n39004) );
  XNOR U11459 ( .A(n39005), .B(n38681), .Z(n38683) );
  XNOR U11460 ( .A(n38684), .B(n38354), .Z(n38356) );
  XNOR U11461 ( .A(n38357), .B(n38021), .Z(n38023) );
  XNOR U11462 ( .A(n38024), .B(n37682), .Z(n37684) );
  XNOR U11463 ( .A(n37685), .B(n37337), .Z(n37339) );
  XNOR U11464 ( .A(n37340), .B(n36986), .Z(n36988) );
  XNOR U11465 ( .A(n36989), .B(n36629), .Z(n36631) );
  XNOR U11466 ( .A(n36632), .B(n36266), .Z(n36268) );
  XNOR U11467 ( .A(n36269), .B(n35897), .Z(n35899) );
  XNOR U11468 ( .A(n35900), .B(n35522), .Z(n35524) );
  XNOR U11469 ( .A(n35525), .B(n35141), .Z(n35143) );
  XNOR U11470 ( .A(n35144), .B(n34754), .Z(n34756) );
  XNOR U11471 ( .A(n34757), .B(n34361), .Z(n34363) );
  XNOR U11472 ( .A(n34364), .B(n33962), .Z(n33964) );
  XNOR U11473 ( .A(n33965), .B(n33557), .Z(n33559) );
  XNOR U11474 ( .A(n33560), .B(n33146), .Z(n33148) );
  XNOR U11475 ( .A(n33149), .B(n32729), .Z(n32731) );
  XNOR U11476 ( .A(n32732), .B(n32306), .Z(n32308) );
  XNOR U11477 ( .A(n32309), .B(n31877), .Z(n31879) );
  XNOR U11478 ( .A(n31880), .B(n31442), .Z(n31444) );
  XNOR U11479 ( .A(n31445), .B(n31001), .Z(n31003) );
  XNOR U11480 ( .A(n31004), .B(n30554), .Z(n30556) );
  XNOR U11481 ( .A(n30557), .B(n30101), .Z(n30103) );
  XNOR U11482 ( .A(n30104), .B(n29642), .Z(n29644) );
  XNOR U11483 ( .A(n29645), .B(n29177), .Z(n29179) );
  XNOR U11484 ( .A(n29180), .B(n28706), .Z(n28708) );
  XNOR U11485 ( .A(n28709), .B(n28229), .Z(n28231) );
  XNOR U11486 ( .A(n28232), .B(n27746), .Z(n27748) );
  XNOR U11487 ( .A(n27749), .B(n27257), .Z(n27259) );
  XNOR U11488 ( .A(n27260), .B(n26760), .Z(n26762) );
  XNOR U11489 ( .A(n26763), .B(n26259), .Z(n26261) );
  XNOR U11490 ( .A(n26262), .B(n25751), .Z(n25753) );
  XNOR U11491 ( .A(n25754), .B(n25237), .Z(n25239) );
  XNOR U11492 ( .A(n25240), .B(n24714), .Z(n24716) );
  XNOR U11493 ( .A(n24717), .B(n24189), .Z(n24191) );
  XNOR U11494 ( .A(n24192), .B(n23658), .Z(n23660) );
  XNOR U11495 ( .A(n23661), .B(n23120), .Z(n23122) );
  XNOR U11496 ( .A(n23123), .B(n22576), .Z(n22578) );
  XNOR U11497 ( .A(n22579), .B(n22027), .Z(n22029) );
  XNOR U11498 ( .A(n22030), .B(n21472), .Z(n21474) );
  XNOR U11499 ( .A(n21475), .B(n20910), .Z(n20912) );
  XNOR U11500 ( .A(n20913), .B(n20343), .Z(n20345) );
  XNOR U11501 ( .A(n20346), .B(n19770), .Z(n19772) );
  XNOR U11502 ( .A(n19773), .B(n19191), .Z(n19193) );
  XOR U11503 ( .A(n17907), .B(n18006), .Z(n17911) );
  XOR U11504 ( .A(n16705), .B(n16804), .Z(n16709) );
  XOR U11505 ( .A(n15479), .B(n15578), .Z(n15483) );
  XOR U11506 ( .A(n14229), .B(n14328), .Z(n14233) );
  XOR U11507 ( .A(n12955), .B(n13054), .Z(n12959) );
  XOR U11508 ( .A(n5480), .B(n5623), .Z(n5484) );
  XOR U11509 ( .A(n4030), .B(n4195), .Z(n4034) );
  XOR U11510 ( .A(n2556), .B(n2745), .Z(n2560) );
  XOR U11511 ( .A(n3251), .B(n3482), .Z(n3255) );
  XOR U11512 ( .A(n1765), .B(n2020), .Z(n1769) );
  XOR U11513 ( .A(n843), .B(n1142), .Z(n853) );
  XOR U11514 ( .A(n12317), .B(n12406), .Z(n12321) );
  XOR U11515 ( .A(n11007), .B(n11094), .Z(n11011) );
  XOR U11516 ( .A(n9673), .B(n9760), .Z(n9677) );
  XOR U11517 ( .A(n8315), .B(n8402), .Z(n8319) );
  XOR U11518 ( .A(n6933), .B(n7020), .Z(n6937) );
  XOR U11519 ( .A(n5525), .B(n5614), .Z(n5529) );
  XOR U11520 ( .A(n857), .B(n1124), .Z(n867) );
  XOR U11521 ( .A(n3281), .B(n3476), .Z(n3285) );
  XOR U11522 ( .A(n1795), .B(n2014), .Z(n1799) );
  XOR U11523 ( .A(n5510), .B(n5617), .Z(n5514) );
  XOR U11524 ( .A(n4060), .B(n4189), .Z(n4064) );
  XOR U11525 ( .A(n2586), .B(n2739), .Z(n2590) );
  XNOR U11526 ( .A(n46940), .B(n46856), .Z(n46858) );
  XNOR U11527 ( .A(n46859), .B(n46769), .Z(n46771) );
  XNOR U11528 ( .A(n46772), .B(n46676), .Z(n46678) );
  XNOR U11529 ( .A(n46679), .B(n46577), .Z(n46579) );
  XNOR U11530 ( .A(n46580), .B(n46472), .Z(n46474) );
  XNOR U11531 ( .A(n46475), .B(n46361), .Z(n46363) );
  XNOR U11532 ( .A(n46364), .B(n46244), .Z(n46246) );
  XNOR U11533 ( .A(n46247), .B(n46121), .Z(n46123) );
  XNOR U11534 ( .A(n46124), .B(n45992), .Z(n45994) );
  XNOR U11535 ( .A(n45995), .B(n45857), .Z(n45859) );
  XNOR U11536 ( .A(n45860), .B(n45716), .Z(n45718) );
  XNOR U11537 ( .A(n45719), .B(n45569), .Z(n45571) );
  XNOR U11538 ( .A(n45572), .B(n45416), .Z(n45418) );
  XNOR U11539 ( .A(n45419), .B(n45257), .Z(n45259) );
  XNOR U11540 ( .A(n45260), .B(n45092), .Z(n45094) );
  XNOR U11541 ( .A(n45095), .B(n44921), .Z(n44923) );
  XNOR U11542 ( .A(n44924), .B(n44744), .Z(n44746) );
  XNOR U11543 ( .A(n44747), .B(n44561), .Z(n44563) );
  XNOR U11544 ( .A(n44564), .B(n44372), .Z(n44374) );
  XNOR U11545 ( .A(n44375), .B(n44177), .Z(n44179) );
  XNOR U11546 ( .A(n44180), .B(n43976), .Z(n43978) );
  XNOR U11547 ( .A(n43979), .B(n43769), .Z(n43771) );
  XNOR U11548 ( .A(n43772), .B(n43556), .Z(n43558) );
  XNOR U11549 ( .A(n43559), .B(n43337), .Z(n43339) );
  XNOR U11550 ( .A(n43340), .B(n43112), .Z(n43114) );
  XNOR U11551 ( .A(n43115), .B(n42881), .Z(n42883) );
  XNOR U11552 ( .A(n42884), .B(n42644), .Z(n42646) );
  XNOR U11553 ( .A(n42647), .B(n42401), .Z(n42403) );
  XNOR U11554 ( .A(n42404), .B(n42152), .Z(n42154) );
  XNOR U11555 ( .A(n42155), .B(n41897), .Z(n41899) );
  XNOR U11556 ( .A(n41900), .B(n41636), .Z(n41638) );
  XNOR U11557 ( .A(n41639), .B(n41369), .Z(n41371) );
  XNOR U11558 ( .A(n41372), .B(n41096), .Z(n41098) );
  XNOR U11559 ( .A(n41099), .B(n40817), .Z(n40819) );
  XNOR U11560 ( .A(n40820), .B(n40532), .Z(n40534) );
  XNOR U11561 ( .A(n40535), .B(n40241), .Z(n40243) );
  XNOR U11562 ( .A(n40244), .B(n39944), .Z(n39946) );
  XNOR U11563 ( .A(n39947), .B(n39641), .Z(n39643) );
  XNOR U11564 ( .A(n39644), .B(n39332), .Z(n39334) );
  XNOR U11565 ( .A(n39335), .B(n39017), .Z(n39019) );
  XNOR U11566 ( .A(n39020), .B(n38696), .Z(n38698) );
  XNOR U11567 ( .A(n38699), .B(n38369), .Z(n38371) );
  XNOR U11568 ( .A(n38372), .B(n38036), .Z(n38038) );
  XNOR U11569 ( .A(n38039), .B(n37697), .Z(n37699) );
  XNOR U11570 ( .A(n37700), .B(n37352), .Z(n37354) );
  XNOR U11571 ( .A(n37355), .B(n37001), .Z(n37003) );
  XNOR U11572 ( .A(n37004), .B(n36644), .Z(n36646) );
  XNOR U11573 ( .A(n36647), .B(n36281), .Z(n36283) );
  XNOR U11574 ( .A(n36284), .B(n35912), .Z(n35914) );
  XNOR U11575 ( .A(n35915), .B(n35537), .Z(n35539) );
  XNOR U11576 ( .A(n35540), .B(n35156), .Z(n35158) );
  XNOR U11577 ( .A(n35159), .B(n34769), .Z(n34771) );
  XNOR U11578 ( .A(n34772), .B(n34376), .Z(n34378) );
  XNOR U11579 ( .A(n34379), .B(n33977), .Z(n33979) );
  XNOR U11580 ( .A(n33980), .B(n33572), .Z(n33574) );
  XNOR U11581 ( .A(n33575), .B(n33161), .Z(n33163) );
  XNOR U11582 ( .A(n33164), .B(n32744), .Z(n32746) );
  XNOR U11583 ( .A(n32747), .B(n32321), .Z(n32323) );
  XNOR U11584 ( .A(n32324), .B(n31892), .Z(n31894) );
  XNOR U11585 ( .A(n31895), .B(n31457), .Z(n31459) );
  XNOR U11586 ( .A(n31460), .B(n31016), .Z(n31018) );
  XNOR U11587 ( .A(n31019), .B(n30569), .Z(n30571) );
  XNOR U11588 ( .A(n30572), .B(n30116), .Z(n30118) );
  XNOR U11589 ( .A(n30119), .B(n29657), .Z(n29659) );
  XNOR U11590 ( .A(n29660), .B(n29192), .Z(n29194) );
  XNOR U11591 ( .A(n29195), .B(n28721), .Z(n28723) );
  XNOR U11592 ( .A(n28724), .B(n28244), .Z(n28246) );
  XNOR U11593 ( .A(n28247), .B(n27761), .Z(n27763) );
  XNOR U11594 ( .A(n27764), .B(n27272), .Z(n27274) );
  XNOR U11595 ( .A(n27275), .B(n26775), .Z(n26777) );
  XNOR U11596 ( .A(n26778), .B(n26274), .Z(n26276) );
  XNOR U11597 ( .A(n26277), .B(n25766), .Z(n25768) );
  XNOR U11598 ( .A(n25769), .B(n25252), .Z(n25254) );
  XNOR U11599 ( .A(n25255), .B(n24729), .Z(n24731) );
  XNOR U11600 ( .A(n24732), .B(n24204), .Z(n24206) );
  XNOR U11601 ( .A(n24207), .B(n23673), .Z(n23675) );
  XNOR U11602 ( .A(n23676), .B(n23135), .Z(n23137) );
  XNOR U11603 ( .A(n23138), .B(n22591), .Z(n22593) );
  XNOR U11604 ( .A(n22594), .B(n22042), .Z(n22044) );
  XNOR U11605 ( .A(n22045), .B(n21487), .Z(n21489) );
  XNOR U11606 ( .A(n21490), .B(n20925), .Z(n20927) );
  XNOR U11607 ( .A(n20928), .B(n20358), .Z(n20360) );
  XNOR U11608 ( .A(n20361), .B(n19785), .Z(n19787) );
  XNOR U11609 ( .A(n19788), .B(n19206), .Z(n19208) );
  XOR U11610 ( .A(n18514), .B(n18613), .Z(n18518) );
  XOR U11611 ( .A(n17324), .B(n17405), .Z(n17328) );
  XOR U11612 ( .A(n16110), .B(n16191), .Z(n16114) );
  XOR U11613 ( .A(n14872), .B(n14953), .Z(n14876) );
  XOR U11614 ( .A(n13610), .B(n13691), .Z(n13614) );
  XOR U11615 ( .A(n4090), .B(n4183), .Z(n4094) );
  XOR U11616 ( .A(n2616), .B(n2733), .Z(n2620) );
  XOR U11617 ( .A(n3311), .B(n3470), .Z(n3315) );
  XOR U11618 ( .A(n1825), .B(n2008), .Z(n1829) );
  XOR U11619 ( .A(n871), .B(n1106), .Z(n881) );
  XOR U11620 ( .A(n12980), .B(n13049), .Z(n12984) );
  XOR U11621 ( .A(n11680), .B(n11749), .Z(n11684) );
  XOR U11622 ( .A(n10358), .B(n10427), .Z(n10362) );
  XOR U11623 ( .A(n9012), .B(n9081), .Z(n9016) );
  XOR U11624 ( .A(n7642), .B(n7711), .Z(n7646) );
  XOR U11625 ( .A(n6248), .B(n6317), .Z(n6252) );
  XOR U11626 ( .A(n4828), .B(n4897), .Z(n4832) );
  XOR U11627 ( .A(n885), .B(n1088), .Z(n895) );
  XOR U11628 ( .A(n3341), .B(n3464), .Z(n3345) );
  XOR U11629 ( .A(n1855), .B(n2002), .Z(n1859) );
  XOR U11630 ( .A(n3386), .B(n3455), .Z(n3390) );
  XNOR U11631 ( .A(n47162), .B(n47096), .Z(n47098) );
  XNOR U11632 ( .A(n47099), .B(n47027), .Z(n47029) );
  XNOR U11633 ( .A(n47030), .B(n46952), .Z(n46954) );
  XNOR U11634 ( .A(n46955), .B(n46871), .Z(n46873) );
  XNOR U11635 ( .A(n46874), .B(n46784), .Z(n46786) );
  XNOR U11636 ( .A(n46787), .B(n46691), .Z(n46693) );
  XNOR U11637 ( .A(n46694), .B(n46592), .Z(n46594) );
  XNOR U11638 ( .A(n46595), .B(n46487), .Z(n46489) );
  XNOR U11639 ( .A(n46490), .B(n46376), .Z(n46378) );
  XNOR U11640 ( .A(n46379), .B(n46259), .Z(n46261) );
  XNOR U11641 ( .A(n46262), .B(n46136), .Z(n46138) );
  XNOR U11642 ( .A(n46139), .B(n46007), .Z(n46009) );
  XNOR U11643 ( .A(n46010), .B(n45872), .Z(n45874) );
  XNOR U11644 ( .A(n45875), .B(n45731), .Z(n45733) );
  XNOR U11645 ( .A(n45734), .B(n45584), .Z(n45586) );
  XNOR U11646 ( .A(n45587), .B(n45431), .Z(n45433) );
  XNOR U11647 ( .A(n45434), .B(n45272), .Z(n45274) );
  XNOR U11648 ( .A(n45275), .B(n45107), .Z(n45109) );
  XNOR U11649 ( .A(n45110), .B(n44936), .Z(n44938) );
  XNOR U11650 ( .A(n44939), .B(n44759), .Z(n44761) );
  XNOR U11651 ( .A(n44762), .B(n44576), .Z(n44578) );
  XNOR U11652 ( .A(n44579), .B(n44387), .Z(n44389) );
  XNOR U11653 ( .A(n44390), .B(n44192), .Z(n44194) );
  XNOR U11654 ( .A(n44195), .B(n43991), .Z(n43993) );
  XNOR U11655 ( .A(n43994), .B(n43784), .Z(n43786) );
  XNOR U11656 ( .A(n43787), .B(n43571), .Z(n43573) );
  XNOR U11657 ( .A(n43574), .B(n43352), .Z(n43354) );
  XNOR U11658 ( .A(n43355), .B(n43127), .Z(n43129) );
  XNOR U11659 ( .A(n43130), .B(n42896), .Z(n42898) );
  XNOR U11660 ( .A(n42899), .B(n42659), .Z(n42661) );
  XNOR U11661 ( .A(n42662), .B(n42416), .Z(n42418) );
  XNOR U11662 ( .A(n42419), .B(n42167), .Z(n42169) );
  XNOR U11663 ( .A(n42170), .B(n41912), .Z(n41914) );
  XNOR U11664 ( .A(n41915), .B(n41651), .Z(n41653) );
  XNOR U11665 ( .A(n41654), .B(n41384), .Z(n41386) );
  XNOR U11666 ( .A(n41387), .B(n41111), .Z(n41113) );
  XNOR U11667 ( .A(n41114), .B(n40832), .Z(n40834) );
  XNOR U11668 ( .A(n40835), .B(n40547), .Z(n40549) );
  XNOR U11669 ( .A(n40550), .B(n40256), .Z(n40258) );
  XNOR U11670 ( .A(n40259), .B(n39959), .Z(n39961) );
  XNOR U11671 ( .A(n39962), .B(n39656), .Z(n39658) );
  XNOR U11672 ( .A(n39659), .B(n39347), .Z(n39349) );
  XNOR U11673 ( .A(n39350), .B(n39032), .Z(n39034) );
  XNOR U11674 ( .A(n39035), .B(n38711), .Z(n38713) );
  XNOR U11675 ( .A(n38714), .B(n38384), .Z(n38386) );
  XNOR U11676 ( .A(n38387), .B(n38051), .Z(n38053) );
  XNOR U11677 ( .A(n38054), .B(n37712), .Z(n37714) );
  XNOR U11678 ( .A(n37715), .B(n37367), .Z(n37369) );
  XNOR U11679 ( .A(n37370), .B(n37016), .Z(n37018) );
  XNOR U11680 ( .A(n37019), .B(n36659), .Z(n36661) );
  XNOR U11681 ( .A(n36662), .B(n36296), .Z(n36298) );
  XNOR U11682 ( .A(n36299), .B(n35927), .Z(n35929) );
  XNOR U11683 ( .A(n35930), .B(n35552), .Z(n35554) );
  XNOR U11684 ( .A(n35555), .B(n35171), .Z(n35173) );
  XNOR U11685 ( .A(n35174), .B(n34784), .Z(n34786) );
  XNOR U11686 ( .A(n34787), .B(n34391), .Z(n34393) );
  XNOR U11687 ( .A(n34394), .B(n33992), .Z(n33994) );
  XNOR U11688 ( .A(n33995), .B(n33587), .Z(n33589) );
  XNOR U11689 ( .A(n33590), .B(n33176), .Z(n33178) );
  XNOR U11690 ( .A(n33179), .B(n32759), .Z(n32761) );
  XNOR U11691 ( .A(n32762), .B(n32336), .Z(n32338) );
  XNOR U11692 ( .A(n32339), .B(n31907), .Z(n31909) );
  XNOR U11693 ( .A(n31910), .B(n31472), .Z(n31474) );
  XNOR U11694 ( .A(n31475), .B(n31031), .Z(n31033) );
  XNOR U11695 ( .A(n31034), .B(n30584), .Z(n30586) );
  XNOR U11696 ( .A(n30587), .B(n30131), .Z(n30133) );
  XNOR U11697 ( .A(n30134), .B(n29672), .Z(n29674) );
  XNOR U11698 ( .A(n29675), .B(n29207), .Z(n29209) );
  XNOR U11699 ( .A(n29210), .B(n28736), .Z(n28738) );
  XNOR U11700 ( .A(n28739), .B(n28259), .Z(n28261) );
  XNOR U11701 ( .A(n28262), .B(n27776), .Z(n27778) );
  XNOR U11702 ( .A(n27779), .B(n27287), .Z(n27289) );
  XNOR U11703 ( .A(n27290), .B(n26790), .Z(n26792) );
  XNOR U11704 ( .A(n26793), .B(n26289), .Z(n26291) );
  XNOR U11705 ( .A(n26292), .B(n25781), .Z(n25783) );
  XNOR U11706 ( .A(n25784), .B(n25267), .Z(n25269) );
  XNOR U11707 ( .A(n25270), .B(n24744), .Z(n24746) );
  XNOR U11708 ( .A(n24747), .B(n24219), .Z(n24221) );
  XNOR U11709 ( .A(n24222), .B(n23688), .Z(n23690) );
  XNOR U11710 ( .A(n23691), .B(n23150), .Z(n23152) );
  XNOR U11711 ( .A(n23153), .B(n22606), .Z(n22608) );
  XNOR U11712 ( .A(n22609), .B(n22057), .Z(n22059) );
  XNOR U11713 ( .A(n22060), .B(n21502), .Z(n21504) );
  XNOR U11714 ( .A(n21505), .B(n20940), .Z(n20942) );
  XNOR U11715 ( .A(n20943), .B(n20373), .Z(n20375) );
  XNOR U11716 ( .A(n20376), .B(n19800), .Z(n19802) );
  XNOR U11717 ( .A(n19803), .B(n19221), .Z(n19223) );
  XOR U11718 ( .A(n18529), .B(n18607), .Z(n18533) );
  XOR U11719 ( .A(n17339), .B(n17402), .Z(n17343) );
  XOR U11720 ( .A(n16125), .B(n16188), .Z(n16129) );
  XOR U11721 ( .A(n14887), .B(n14950), .Z(n14891) );
  XOR U11722 ( .A(n1905), .B(n1992), .Z(n1909) );
  XOR U11723 ( .A(n3371), .B(n3458), .Z(n3375) );
  XOR U11724 ( .A(n1885), .B(n1996), .Z(n1889) );
  XOR U11725 ( .A(n899), .B(n1070), .Z(n909) );
  XOR U11726 ( .A(n14269), .B(n14320), .Z(n14273) );
  XOR U11727 ( .A(n12995), .B(n13046), .Z(n12999) );
  XOR U11728 ( .A(n11695), .B(n11746), .Z(n11699) );
  XOR U11729 ( .A(n10373), .B(n10424), .Z(n10377) );
  XOR U11730 ( .A(n9027), .B(n9078), .Z(n9031) );
  XOR U11731 ( .A(n7657), .B(n7708), .Z(n7661) );
  XOR U11732 ( .A(n6263), .B(n6314), .Z(n6267) );
  XOR U11733 ( .A(n4843), .B(n4894), .Z(n4847) );
  XOR U11734 ( .A(n3401), .B(n3452), .Z(n3405) );
  XOR U11735 ( .A(n1935), .B(n1986), .Z(n1939) );
  XOR U11736 ( .A(n913), .B(n1052), .Z(n923) );
  XNOR U11737 ( .A(n47329), .B(n47281), .Z(n47283) );
  XNOR U11738 ( .A(n47284), .B(n47230), .Z(n47232) );
  XNOR U11739 ( .A(n47233), .B(n47174), .Z(n47176) );
  XNOR U11740 ( .A(n47177), .B(n47111), .Z(n47113) );
  XNOR U11741 ( .A(n47114), .B(n47042), .Z(n47044) );
  XNOR U11742 ( .A(n47045), .B(n46967), .Z(n46969) );
  XNOR U11743 ( .A(n46970), .B(n46886), .Z(n46888) );
  XNOR U11744 ( .A(n46889), .B(n46799), .Z(n46801) );
  XNOR U11745 ( .A(n46802), .B(n46706), .Z(n46708) );
  XNOR U11746 ( .A(n46709), .B(n46607), .Z(n46609) );
  XNOR U11747 ( .A(n46610), .B(n46502), .Z(n46504) );
  XNOR U11748 ( .A(n46505), .B(n46391), .Z(n46393) );
  XNOR U11749 ( .A(n46394), .B(n46274), .Z(n46276) );
  XNOR U11750 ( .A(n46277), .B(n46151), .Z(n46153) );
  XNOR U11751 ( .A(n46154), .B(n46022), .Z(n46024) );
  XNOR U11752 ( .A(n46025), .B(n45887), .Z(n45889) );
  XNOR U11753 ( .A(n45890), .B(n45746), .Z(n45748) );
  XNOR U11754 ( .A(n45749), .B(n45599), .Z(n45601) );
  XNOR U11755 ( .A(n45602), .B(n45446), .Z(n45448) );
  XNOR U11756 ( .A(n45449), .B(n45287), .Z(n45289) );
  XNOR U11757 ( .A(n45290), .B(n45122), .Z(n45124) );
  XNOR U11758 ( .A(n45125), .B(n44951), .Z(n44953) );
  XNOR U11759 ( .A(n44954), .B(n44774), .Z(n44776) );
  XNOR U11760 ( .A(n44777), .B(n44591), .Z(n44593) );
  XNOR U11761 ( .A(n44594), .B(n44402), .Z(n44404) );
  XNOR U11762 ( .A(n44405), .B(n44207), .Z(n44209) );
  XNOR U11763 ( .A(n44210), .B(n44006), .Z(n44008) );
  XNOR U11764 ( .A(n44009), .B(n43799), .Z(n43801) );
  XNOR U11765 ( .A(n43802), .B(n43586), .Z(n43588) );
  XNOR U11766 ( .A(n43589), .B(n43367), .Z(n43369) );
  XNOR U11767 ( .A(n43370), .B(n43142), .Z(n43144) );
  XNOR U11768 ( .A(n43145), .B(n42911), .Z(n42913) );
  XNOR U11769 ( .A(n42914), .B(n42674), .Z(n42676) );
  XNOR U11770 ( .A(n42677), .B(n42431), .Z(n42433) );
  XNOR U11771 ( .A(n42434), .B(n42182), .Z(n42184) );
  XNOR U11772 ( .A(n42185), .B(n41927), .Z(n41929) );
  XNOR U11773 ( .A(n41930), .B(n41666), .Z(n41668) );
  XNOR U11774 ( .A(n41669), .B(n41399), .Z(n41401) );
  XNOR U11775 ( .A(n41402), .B(n41126), .Z(n41128) );
  XNOR U11776 ( .A(n41129), .B(n40847), .Z(n40849) );
  XNOR U11777 ( .A(n40850), .B(n40562), .Z(n40564) );
  XNOR U11778 ( .A(n40565), .B(n40271), .Z(n40273) );
  XNOR U11779 ( .A(n40274), .B(n39974), .Z(n39976) );
  XNOR U11780 ( .A(n39977), .B(n39671), .Z(n39673) );
  XNOR U11781 ( .A(n39674), .B(n39362), .Z(n39364) );
  XNOR U11782 ( .A(n39365), .B(n39047), .Z(n39049) );
  XNOR U11783 ( .A(n39050), .B(n38726), .Z(n38728) );
  XNOR U11784 ( .A(n38729), .B(n38399), .Z(n38401) );
  XNOR U11785 ( .A(n38402), .B(n38066), .Z(n38068) );
  XNOR U11786 ( .A(n38069), .B(n37727), .Z(n37729) );
  XNOR U11787 ( .A(n37730), .B(n37382), .Z(n37384) );
  XNOR U11788 ( .A(n37385), .B(n37031), .Z(n37033) );
  XNOR U11789 ( .A(n37034), .B(n36674), .Z(n36676) );
  XNOR U11790 ( .A(n36677), .B(n36311), .Z(n36313) );
  XNOR U11791 ( .A(n36314), .B(n35942), .Z(n35944) );
  XNOR U11792 ( .A(n35945), .B(n35567), .Z(n35569) );
  XNOR U11793 ( .A(n35570), .B(n35186), .Z(n35188) );
  XNOR U11794 ( .A(n35189), .B(n34799), .Z(n34801) );
  XNOR U11795 ( .A(n34802), .B(n34406), .Z(n34408) );
  XNOR U11796 ( .A(n34409), .B(n34007), .Z(n34009) );
  XNOR U11797 ( .A(n34010), .B(n33602), .Z(n33604) );
  XNOR U11798 ( .A(n33605), .B(n33191), .Z(n33193) );
  XNOR U11799 ( .A(n33194), .B(n32774), .Z(n32776) );
  XNOR U11800 ( .A(n32777), .B(n32351), .Z(n32353) );
  XNOR U11801 ( .A(n32354), .B(n31922), .Z(n31924) );
  XNOR U11802 ( .A(n31925), .B(n31487), .Z(n31489) );
  XNOR U11803 ( .A(n31490), .B(n31046), .Z(n31048) );
  XNOR U11804 ( .A(n31049), .B(n30599), .Z(n30601) );
  XNOR U11805 ( .A(n30602), .B(n30146), .Z(n30148) );
  XNOR U11806 ( .A(n30149), .B(n29687), .Z(n29689) );
  XNOR U11807 ( .A(n29690), .B(n29222), .Z(n29224) );
  XNOR U11808 ( .A(n29225), .B(n28751), .Z(n28753) );
  XNOR U11809 ( .A(n28754), .B(n28274), .Z(n28276) );
  XNOR U11810 ( .A(n28277), .B(n27791), .Z(n27793) );
  XNOR U11811 ( .A(n27794), .B(n27302), .Z(n27304) );
  XNOR U11812 ( .A(n27305), .B(n26805), .Z(n26807) );
  XNOR U11813 ( .A(n26808), .B(n26304), .Z(n26306) );
  XNOR U11814 ( .A(n26307), .B(n25796), .Z(n25798) );
  XNOR U11815 ( .A(n25799), .B(n25282), .Z(n25284) );
  XNOR U11816 ( .A(n25285), .B(n24759), .Z(n24761) );
  XNOR U11817 ( .A(n24762), .B(n24234), .Z(n24236) );
  XNOR U11818 ( .A(n24237), .B(n23703), .Z(n23705) );
  XNOR U11819 ( .A(n23706), .B(n23165), .Z(n23167) );
  XNOR U11820 ( .A(n23168), .B(n22621), .Z(n22623) );
  XNOR U11821 ( .A(n22624), .B(n22072), .Z(n22074) );
  XNOR U11822 ( .A(n22075), .B(n21517), .Z(n21519) );
  XNOR U11823 ( .A(n21520), .B(n20955), .Z(n20957) );
  XNOR U11824 ( .A(n20958), .B(n20388), .Z(n20390) );
  XNOR U11825 ( .A(n20391), .B(n19815), .Z(n19817) );
  XNOR U11826 ( .A(n19818), .B(n19236), .Z(n19238) );
  XOR U11827 ( .A(n18544), .B(n18601), .Z(n18548) );
  XOR U11828 ( .A(n17354), .B(n17399), .Z(n17358) );
  XOR U11829 ( .A(n16140), .B(n16185), .Z(n16144) );
  XOR U11830 ( .A(n1920), .B(n1989), .Z(n1924) );
  XOR U11831 ( .A(n927), .B(n1034), .Z(n937) );
  XOR U11832 ( .A(n15534), .B(n15567), .Z(n15538) );
  XOR U11833 ( .A(n14284), .B(n14317), .Z(n14288) );
  XOR U11834 ( .A(n13010), .B(n13043), .Z(n13014) );
  XOR U11835 ( .A(n11710), .B(n11743), .Z(n11714) );
  XOR U11836 ( .A(n10388), .B(n10421), .Z(n10392) );
  XOR U11837 ( .A(n9042), .B(n9075), .Z(n9046) );
  XOR U11838 ( .A(n7672), .B(n7705), .Z(n7676) );
  XOR U11839 ( .A(n6278), .B(n6311), .Z(n6282) );
  XOR U11840 ( .A(n4858), .B(n4891), .Z(n4862) );
  XOR U11841 ( .A(n3416), .B(n3449), .Z(n3420) );
  XOR U11842 ( .A(n1950), .B(n1983), .Z(n1954) );
  XNOR U11843 ( .A(n47443), .B(n47413), .Z(n47415) );
  XNOR U11844 ( .A(n47416), .B(n47380), .Z(n47382) );
  XNOR U11845 ( .A(n47383), .B(n47341), .Z(n47343) );
  XNOR U11846 ( .A(n47344), .B(n47296), .Z(n47298) );
  XNOR U11847 ( .A(n47299), .B(n47245), .Z(n47247) );
  XNOR U11848 ( .A(n47248), .B(n47189), .Z(n47191) );
  XNOR U11849 ( .A(n47192), .B(n47126), .Z(n47128) );
  XNOR U11850 ( .A(n47129), .B(n47057), .Z(n47059) );
  XNOR U11851 ( .A(n47060), .B(n46982), .Z(n46984) );
  XNOR U11852 ( .A(n46985), .B(n46901), .Z(n46903) );
  XNOR U11853 ( .A(n46904), .B(n46814), .Z(n46816) );
  XNOR U11854 ( .A(n46817), .B(n46721), .Z(n46723) );
  XNOR U11855 ( .A(n46724), .B(n46622), .Z(n46624) );
  XNOR U11856 ( .A(n46625), .B(n46517), .Z(n46519) );
  XNOR U11857 ( .A(n46520), .B(n46406), .Z(n46408) );
  XNOR U11858 ( .A(n46409), .B(n46289), .Z(n46291) );
  XNOR U11859 ( .A(n46292), .B(n46166), .Z(n46168) );
  XNOR U11860 ( .A(n46169), .B(n46037), .Z(n46039) );
  XNOR U11861 ( .A(n46040), .B(n45902), .Z(n45904) );
  XNOR U11862 ( .A(n45905), .B(n45761), .Z(n45763) );
  XNOR U11863 ( .A(n45764), .B(n45614), .Z(n45616) );
  XNOR U11864 ( .A(n45617), .B(n45461), .Z(n45463) );
  XNOR U11865 ( .A(n45464), .B(n45302), .Z(n45304) );
  XNOR U11866 ( .A(n45305), .B(n45137), .Z(n45139) );
  XNOR U11867 ( .A(n45140), .B(n44966), .Z(n44968) );
  XNOR U11868 ( .A(n44969), .B(n44789), .Z(n44791) );
  XNOR U11869 ( .A(n44792), .B(n44606), .Z(n44608) );
  XNOR U11870 ( .A(n44609), .B(n44417), .Z(n44419) );
  XNOR U11871 ( .A(n44420), .B(n44222), .Z(n44224) );
  XNOR U11872 ( .A(n44225), .B(n44021), .Z(n44023) );
  XNOR U11873 ( .A(n44024), .B(n43814), .Z(n43816) );
  XNOR U11874 ( .A(n43817), .B(n43601), .Z(n43603) );
  XNOR U11875 ( .A(n43604), .B(n43382), .Z(n43384) );
  XNOR U11876 ( .A(n43385), .B(n43157), .Z(n43159) );
  XNOR U11877 ( .A(n43160), .B(n42926), .Z(n42928) );
  XNOR U11878 ( .A(n42929), .B(n42689), .Z(n42691) );
  XNOR U11879 ( .A(n42692), .B(n42446), .Z(n42448) );
  XNOR U11880 ( .A(n42449), .B(n42197), .Z(n42199) );
  XNOR U11881 ( .A(n42200), .B(n41942), .Z(n41944) );
  XNOR U11882 ( .A(n41945), .B(n41681), .Z(n41683) );
  XNOR U11883 ( .A(n41684), .B(n41414), .Z(n41416) );
  XNOR U11884 ( .A(n41417), .B(n41141), .Z(n41143) );
  XNOR U11885 ( .A(n41144), .B(n40862), .Z(n40864) );
  XNOR U11886 ( .A(n40865), .B(n40577), .Z(n40579) );
  XNOR U11887 ( .A(n40580), .B(n40286), .Z(n40288) );
  XNOR U11888 ( .A(n40289), .B(n39989), .Z(n39991) );
  XNOR U11889 ( .A(n39992), .B(n39686), .Z(n39688) );
  XNOR U11890 ( .A(n39689), .B(n39377), .Z(n39379) );
  XNOR U11891 ( .A(n39380), .B(n39062), .Z(n39064) );
  XNOR U11892 ( .A(n39065), .B(n38741), .Z(n38743) );
  XNOR U11893 ( .A(n38744), .B(n38414), .Z(n38416) );
  XNOR U11894 ( .A(n38417), .B(n38081), .Z(n38083) );
  XNOR U11895 ( .A(n38084), .B(n37742), .Z(n37744) );
  XNOR U11896 ( .A(n37745), .B(n37397), .Z(n37399) );
  XNOR U11897 ( .A(n37400), .B(n37046), .Z(n37048) );
  XNOR U11898 ( .A(n37049), .B(n36689), .Z(n36691) );
  XNOR U11899 ( .A(n36692), .B(n36326), .Z(n36328) );
  XNOR U11900 ( .A(n36329), .B(n35957), .Z(n35959) );
  XNOR U11901 ( .A(n35960), .B(n35582), .Z(n35584) );
  XNOR U11902 ( .A(n35585), .B(n35201), .Z(n35203) );
  XNOR U11903 ( .A(n35204), .B(n34814), .Z(n34816) );
  XNOR U11904 ( .A(n34817), .B(n34421), .Z(n34423) );
  XNOR U11905 ( .A(n34424), .B(n34022), .Z(n34024) );
  XNOR U11906 ( .A(n34025), .B(n33617), .Z(n33619) );
  XNOR U11907 ( .A(n33620), .B(n33206), .Z(n33208) );
  XNOR U11908 ( .A(n33209), .B(n32789), .Z(n32791) );
  XNOR U11909 ( .A(n32792), .B(n32366), .Z(n32368) );
  XNOR U11910 ( .A(n32369), .B(n31937), .Z(n31939) );
  XNOR U11911 ( .A(n31940), .B(n31502), .Z(n31504) );
  XNOR U11912 ( .A(n31505), .B(n31061), .Z(n31063) );
  XNOR U11913 ( .A(n31064), .B(n30614), .Z(n30616) );
  XNOR U11914 ( .A(n30617), .B(n30161), .Z(n30163) );
  XNOR U11915 ( .A(n30164), .B(n29702), .Z(n29704) );
  XNOR U11916 ( .A(n29705), .B(n29237), .Z(n29239) );
  XNOR U11917 ( .A(n29240), .B(n28766), .Z(n28768) );
  XNOR U11918 ( .A(n28769), .B(n28289), .Z(n28291) );
  XNOR U11919 ( .A(n28292), .B(n27806), .Z(n27808) );
  XNOR U11920 ( .A(n27809), .B(n27317), .Z(n27319) );
  XNOR U11921 ( .A(n27320), .B(n26820), .Z(n26822) );
  XNOR U11922 ( .A(n26823), .B(n26319), .Z(n26321) );
  XNOR U11923 ( .A(n26322), .B(n25811), .Z(n25813) );
  XNOR U11924 ( .A(n25814), .B(n25297), .Z(n25299) );
  XNOR U11925 ( .A(n25300), .B(n24774), .Z(n24776) );
  XNOR U11926 ( .A(n24777), .B(n24249), .Z(n24251) );
  XNOR U11927 ( .A(n24252), .B(n23718), .Z(n23720) );
  XNOR U11928 ( .A(n23721), .B(n23180), .Z(n23182) );
  XNOR U11929 ( .A(n23183), .B(n22636), .Z(n22638) );
  XNOR U11930 ( .A(n22639), .B(n22087), .Z(n22089) );
  XNOR U11931 ( .A(n22090), .B(n21532), .Z(n21534) );
  XNOR U11932 ( .A(n21535), .B(n20970), .Z(n20972) );
  XNOR U11933 ( .A(n20973), .B(n20403), .Z(n20405) );
  XNOR U11934 ( .A(n20406), .B(n19830), .Z(n19832) );
  XNOR U11935 ( .A(n19833), .B(n19251), .Z(n19253) );
  XOR U11936 ( .A(n18559), .B(n18595), .Z(n18563) );
  XOR U11937 ( .A(n17369), .B(n17396), .Z(n17373) );
  XOR U11938 ( .A(n16775), .B(n16790), .Z(n16784) );
  XOR U11939 ( .A(n15549), .B(n15564), .Z(n15558) );
  XOR U11940 ( .A(n14299), .B(n14314), .Z(n14308) );
  XOR U11941 ( .A(n13025), .B(n13040), .Z(n13034) );
  XOR U11942 ( .A(n11725), .B(n11740), .Z(n11734) );
  XOR U11943 ( .A(n10403), .B(n10418), .Z(n10412) );
  XOR U11944 ( .A(n9057), .B(n9072), .Z(n9066) );
  XOR U11945 ( .A(n7687), .B(n7702), .Z(n7696) );
  XOR U11946 ( .A(n6293), .B(n6308), .Z(n6302) );
  XOR U11947 ( .A(n4873), .B(n4888), .Z(n4882) );
  XOR U11948 ( .A(n3431), .B(n3446), .Z(n3440) );
  XOR U11949 ( .A(n1965), .B(n1980), .Z(n1974) );
  XNOR U11950 ( .A(n47479), .B(n47476), .Z(n47461) );
  XNOR U11951 ( .A(n47458), .B(n47455), .Z(n47434) );
  XNOR U11952 ( .A(n47431), .B(n47428), .Z(n47401) );
  XNOR U11953 ( .A(n47398), .B(n47395), .Z(n47362) );
  XNOR U11954 ( .A(n47359), .B(n47356), .Z(n47317) );
  XNOR U11955 ( .A(n47314), .B(n47311), .Z(n47266) );
  XNOR U11956 ( .A(n47206), .B(n47204), .Z(n47147) );
  XNOR U11957 ( .A(n47144), .B(n47141), .Z(n47078) );
  XNOR U11958 ( .A(n47075), .B(n47072), .Z(n47003) );
  XNOR U11959 ( .A(n47000), .B(n46997), .Z(n46922) );
  XNOR U11960 ( .A(n46919), .B(n46916), .Z(n46835) );
  XNOR U11961 ( .A(n46832), .B(n46829), .Z(n46742) );
  XNOR U11962 ( .A(n46739), .B(n46736), .Z(n46643) );
  XNOR U11963 ( .A(n46640), .B(n46637), .Z(n46538) );
  XNOR U11964 ( .A(n46535), .B(n46532), .Z(n46427) );
  XNOR U11965 ( .A(n46424), .B(n46421), .Z(n46310) );
  XNOR U11966 ( .A(n46307), .B(n46304), .Z(n46187) );
  XNOR U11967 ( .A(n46184), .B(n46181), .Z(n46058) );
  XNOR U11968 ( .A(n46055), .B(n46052), .Z(n45923) );
  XNOR U11969 ( .A(n45920), .B(n45917), .Z(n45782) );
  XNOR U11970 ( .A(n45779), .B(n45776), .Z(n45635) );
  XNOR U11971 ( .A(n45632), .B(n45629), .Z(n45482) );
  XNOR U11972 ( .A(n45479), .B(n45476), .Z(n45323) );
  XNOR U11973 ( .A(n45320), .B(n45317), .Z(n45158) );
  XNOR U11974 ( .A(n45155), .B(n45152), .Z(n44987) );
  XNOR U11975 ( .A(n44984), .B(n44981), .Z(n44810) );
  XNOR U11976 ( .A(n44807), .B(n44804), .Z(n44627) );
  XNOR U11977 ( .A(n44624), .B(n44621), .Z(n44438) );
  XNOR U11978 ( .A(n44435), .B(n44432), .Z(n44243) );
  XNOR U11979 ( .A(n44240), .B(n44237), .Z(n44042) );
  XNOR U11980 ( .A(n44039), .B(n44036), .Z(n43835) );
  XNOR U11981 ( .A(n43832), .B(n43829), .Z(n43622) );
  XNOR U11982 ( .A(n43619), .B(n43616), .Z(n43403) );
  XNOR U11983 ( .A(n43400), .B(n43397), .Z(n43178) );
  XNOR U11984 ( .A(n43175), .B(n43172), .Z(n42947) );
  XNOR U11985 ( .A(n42944), .B(n42941), .Z(n42710) );
  XNOR U11986 ( .A(n42707), .B(n42704), .Z(n42467) );
  XNOR U11987 ( .A(n42464), .B(n42461), .Z(n42218) );
  XNOR U11988 ( .A(n42215), .B(n42212), .Z(n41963) );
  XNOR U11989 ( .A(n41960), .B(n41957), .Z(n41702) );
  XNOR U11990 ( .A(n41699), .B(n41696), .Z(n41435) );
  XNOR U11991 ( .A(n41432), .B(n41429), .Z(n41162) );
  XNOR U11992 ( .A(n41159), .B(n41156), .Z(n40883) );
  XNOR U11993 ( .A(n40880), .B(n40877), .Z(n40598) );
  XNOR U11994 ( .A(n40595), .B(n40592), .Z(n40307) );
  XNOR U11995 ( .A(n40304), .B(n40301), .Z(n40010) );
  XNOR U11996 ( .A(n40007), .B(n40004), .Z(n39707) );
  XNOR U11997 ( .A(n39704), .B(n39701), .Z(n39398) );
  XNOR U11998 ( .A(n39395), .B(n39392), .Z(n39083) );
  XNOR U11999 ( .A(n39080), .B(n39077), .Z(n38762) );
  XNOR U12000 ( .A(n38759), .B(n38756), .Z(n38435) );
  XNOR U12001 ( .A(n38432), .B(n38429), .Z(n38102) );
  XNOR U12002 ( .A(n38099), .B(n38096), .Z(n37763) );
  XNOR U12003 ( .A(n37760), .B(n37757), .Z(n37418) );
  XNOR U12004 ( .A(n37415), .B(n37412), .Z(n37067) );
  XNOR U12005 ( .A(n37064), .B(n37061), .Z(n36710) );
  XNOR U12006 ( .A(n36707), .B(n36704), .Z(n36347) );
  XNOR U12007 ( .A(n36344), .B(n36341), .Z(n35978) );
  XNOR U12008 ( .A(n35975), .B(n35972), .Z(n35603) );
  XNOR U12009 ( .A(n35600), .B(n35597), .Z(n35222) );
  XNOR U12010 ( .A(n35219), .B(n35216), .Z(n34835) );
  XNOR U12011 ( .A(n34832), .B(n34829), .Z(n34442) );
  XNOR U12012 ( .A(n34439), .B(n34436), .Z(n34043) );
  XNOR U12013 ( .A(n34040), .B(n34037), .Z(n33638) );
  XNOR U12014 ( .A(n33635), .B(n33632), .Z(n33227) );
  XNOR U12015 ( .A(n33224), .B(n33221), .Z(n32810) );
  XNOR U12016 ( .A(n32807), .B(n32804), .Z(n32387) );
  XNOR U12017 ( .A(n32384), .B(n32381), .Z(n31958) );
  XNOR U12018 ( .A(n31955), .B(n31952), .Z(n31523) );
  XNOR U12019 ( .A(n31520), .B(n31517), .Z(n31082) );
  XNOR U12020 ( .A(n31079), .B(n31076), .Z(n30635) );
  XNOR U12021 ( .A(n30632), .B(n30629), .Z(n30182) );
  XNOR U12022 ( .A(n30179), .B(n30176), .Z(n29723) );
  XNOR U12023 ( .A(n29720), .B(n29717), .Z(n29258) );
  XNOR U12024 ( .A(n29255), .B(n29252), .Z(n28787) );
  XNOR U12025 ( .A(n28784), .B(n28781), .Z(n28310) );
  XNOR U12026 ( .A(n28307), .B(n28304), .Z(n27827) );
  XNOR U12027 ( .A(n27824), .B(n27821), .Z(n27338) );
  XNOR U12028 ( .A(n27335), .B(n27332), .Z(n26841) );
  XNOR U12029 ( .A(n26838), .B(n26835), .Z(n26340) );
  XNOR U12030 ( .A(n26337), .B(n26334), .Z(n25832) );
  XNOR U12031 ( .A(n25829), .B(n25826), .Z(n25318) );
  XNOR U12032 ( .A(n25315), .B(n25312), .Z(n24795) );
  XNOR U12033 ( .A(n24792), .B(n24789), .Z(n24270) );
  XNOR U12034 ( .A(n24267), .B(n24264), .Z(n23739) );
  XNOR U12035 ( .A(n23736), .B(n23733), .Z(n23201) );
  XNOR U12036 ( .A(n23198), .B(n23195), .Z(n22657) );
  XNOR U12037 ( .A(n22654), .B(n22651), .Z(n22108) );
  XNOR U12038 ( .A(n22105), .B(n22102), .Z(n21553) );
  XNOR U12039 ( .A(n21550), .B(n21547), .Z(n20991) );
  XNOR U12040 ( .A(n20988), .B(n20985), .Z(n20424) );
  XNOR U12041 ( .A(n20421), .B(n20418), .Z(n19851) );
  XNOR U12042 ( .A(n19848), .B(n19845), .Z(n19272) );
  XNOR U12043 ( .A(n19269), .B(n19266), .Z(n18592) );
  XNOR U12044 ( .A(n18575), .B(n18573), .Z(n17991) );
  XOR U12045 ( .A(n1), .B(n2), .Z(c[9]) );
  XOR U12046 ( .A(n3), .B(n4), .Z(c[99]) );
  XNOR U12047 ( .A(n5), .B(n6), .Z(c[98]) );
  XNOR U12048 ( .A(n7), .B(n8), .Z(c[97]) );
  XNOR U12049 ( .A(n9), .B(n10), .Z(c[96]) );
  XNOR U12050 ( .A(n11), .B(n12), .Z(c[95]) );
  XNOR U12051 ( .A(n13), .B(n14), .Z(c[94]) );
  XNOR U12052 ( .A(n15), .B(n16), .Z(c[93]) );
  XNOR U12053 ( .A(n17), .B(n18), .Z(c[92]) );
  XNOR U12054 ( .A(n19), .B(n20), .Z(c[91]) );
  XNOR U12055 ( .A(n21), .B(n22), .Z(c[90]) );
  XNOR U12056 ( .A(n23), .B(n24), .Z(c[8]) );
  XNOR U12057 ( .A(n25), .B(n26), .Z(c[89]) );
  XNOR U12058 ( .A(n27), .B(n28), .Z(c[88]) );
  XNOR U12059 ( .A(n29), .B(n30), .Z(c[87]) );
  XNOR U12060 ( .A(n31), .B(n32), .Z(c[86]) );
  XNOR U12061 ( .A(n33), .B(n34), .Z(c[85]) );
  XNOR U12062 ( .A(n35), .B(n36), .Z(c[84]) );
  XNOR U12063 ( .A(n37), .B(n38), .Z(c[83]) );
  XNOR U12064 ( .A(n39), .B(n40), .Z(c[82]) );
  XNOR U12065 ( .A(n41), .B(n42), .Z(c[81]) );
  XNOR U12066 ( .A(n43), .B(n44), .Z(c[80]) );
  XNOR U12067 ( .A(n45), .B(n46), .Z(c[7]) );
  XNOR U12068 ( .A(n47), .B(n48), .Z(c[79]) );
  XNOR U12069 ( .A(n49), .B(n50), .Z(c[78]) );
  XNOR U12070 ( .A(n51), .B(n52), .Z(c[77]) );
  XNOR U12071 ( .A(n53), .B(n54), .Z(c[76]) );
  XNOR U12072 ( .A(n55), .B(n56), .Z(c[75]) );
  XNOR U12073 ( .A(n57), .B(n58), .Z(c[74]) );
  XNOR U12074 ( .A(n59), .B(n60), .Z(c[73]) );
  XNOR U12075 ( .A(n61), .B(n62), .Z(c[72]) );
  XNOR U12076 ( .A(n63), .B(n64), .Z(c[71]) );
  XNOR U12077 ( .A(n65), .B(n66), .Z(c[70]) );
  XNOR U12078 ( .A(n67), .B(n68), .Z(c[6]) );
  XNOR U12079 ( .A(n69), .B(n70), .Z(c[69]) );
  XNOR U12080 ( .A(n71), .B(n72), .Z(c[68]) );
  XNOR U12081 ( .A(n73), .B(n74), .Z(c[67]) );
  XNOR U12082 ( .A(n75), .B(n76), .Z(c[66]) );
  XNOR U12083 ( .A(n77), .B(n78), .Z(c[65]) );
  XNOR U12084 ( .A(n79), .B(n80), .Z(c[64]) );
  XNOR U12085 ( .A(n81), .B(n82), .Z(c[63]) );
  XNOR U12086 ( .A(n83), .B(n84), .Z(c[62]) );
  XNOR U12087 ( .A(n85), .B(n86), .Z(c[61]) );
  XNOR U12088 ( .A(n87), .B(n88), .Z(c[60]) );
  XNOR U12089 ( .A(n89), .B(n90), .Z(c[5]) );
  XNOR U12090 ( .A(n91), .B(n92), .Z(c[59]) );
  XNOR U12091 ( .A(n93), .B(n94), .Z(c[58]) );
  XNOR U12092 ( .A(n95), .B(n96), .Z(c[57]) );
  XNOR U12093 ( .A(n97), .B(n98), .Z(c[56]) );
  XNOR U12094 ( .A(n99), .B(n100), .Z(c[55]) );
  XNOR U12095 ( .A(n101), .B(n102), .Z(c[54]) );
  XNOR U12096 ( .A(n103), .B(n104), .Z(c[53]) );
  XNOR U12097 ( .A(n105), .B(n106), .Z(c[52]) );
  XNOR U12098 ( .A(n107), .B(n108), .Z(c[51]) );
  XNOR U12099 ( .A(n109), .B(n110), .Z(c[50]) );
  XNOR U12100 ( .A(n111), .B(n112), .Z(c[4]) );
  XNOR U12101 ( .A(n113), .B(n114), .Z(c[49]) );
  XNOR U12102 ( .A(n115), .B(n116), .Z(c[48]) );
  XNOR U12103 ( .A(n117), .B(n118), .Z(c[47]) );
  XNOR U12104 ( .A(n119), .B(n120), .Z(c[46]) );
  XNOR U12105 ( .A(n121), .B(n122), .Z(c[45]) );
  XNOR U12106 ( .A(n123), .B(n124), .Z(c[44]) );
  XNOR U12107 ( .A(n125), .B(n126), .Z(c[43]) );
  XNOR U12108 ( .A(n127), .B(n128), .Z(c[42]) );
  XNOR U12109 ( .A(n129), .B(n130), .Z(c[41]) );
  XNOR U12110 ( .A(n131), .B(n132), .Z(c[40]) );
  XNOR U12111 ( .A(n133), .B(n134), .Z(c[3]) );
  XNOR U12112 ( .A(n135), .B(n136), .Z(c[39]) );
  XNOR U12113 ( .A(n137), .B(n138), .Z(c[38]) );
  XNOR U12114 ( .A(n139), .B(n140), .Z(c[37]) );
  XNOR U12115 ( .A(n141), .B(n142), .Z(c[36]) );
  XNOR U12116 ( .A(n143), .B(n144), .Z(c[35]) );
  XNOR U12117 ( .A(n145), .B(n146), .Z(c[34]) );
  XNOR U12118 ( .A(n147), .B(n148), .Z(c[33]) );
  XNOR U12119 ( .A(n149), .B(n150), .Z(c[32]) );
  XNOR U12120 ( .A(n151), .B(n152), .Z(c[31]) );
  XNOR U12121 ( .A(n153), .B(n154), .Z(c[30]) );
  XNOR U12122 ( .A(n155), .B(n156), .Z(c[2]) );
  XNOR U12123 ( .A(n157), .B(n158), .Z(c[29]) );
  XNOR U12124 ( .A(n159), .B(n160), .Z(c[28]) );
  XNOR U12125 ( .A(n161), .B(n162), .Z(c[27]) );
  XNOR U12126 ( .A(n163), .B(n164), .Z(c[26]) );
  XNOR U12127 ( .A(n165), .B(n166), .Z(c[25]) );
  XNOR U12128 ( .A(n167), .B(n168), .Z(c[24]) );
  XNOR U12129 ( .A(n169), .B(n170), .Z(c[23]) );
  XNOR U12130 ( .A(n171), .B(n172), .Z(c[22]) );
  XNOR U12131 ( .A(n173), .B(n174), .Z(c[21]) );
  XNOR U12132 ( .A(n175), .B(n176), .Z(c[20]) );
  XOR U12133 ( .A(n177), .B(n178), .Z(c[1]) );
  XNOR U12134 ( .A(n179), .B(n180), .Z(c[19]) );
  XNOR U12135 ( .A(n181), .B(n182), .Z(c[18]) );
  XNOR U12136 ( .A(n183), .B(n184), .Z(c[17]) );
  XNOR U12137 ( .A(n185), .B(n186), .Z(c[16]) );
  XNOR U12138 ( .A(n187), .B(n188), .Z(c[15]) );
  XNOR U12139 ( .A(n189), .B(n190), .Z(c[14]) );
  XNOR U12140 ( .A(n191), .B(n192), .Z(c[13]) );
  XNOR U12141 ( .A(n193), .B(n194), .Z(c[12]) );
  XOR U12142 ( .A(n195), .B(n196), .Z(c[127]) );
  XOR U12143 ( .A(n197), .B(n198), .Z(n196) );
  XOR U12144 ( .A(n199), .B(n200), .Z(n198) );
  XOR U12145 ( .A(n201), .B(n202), .Z(n200) );
  XOR U12146 ( .A(n203), .B(n204), .Z(n202) );
  XNOR U12147 ( .A(n205), .B(n206), .Z(n204) );
  AND U12148 ( .A(b[1]), .B(a[126]), .Z(n206) );
  XOR U12149 ( .A(n207), .B(n208), .Z(n203) );
  XOR U12150 ( .A(n209), .B(n210), .Z(n208) );
  XOR U12151 ( .A(n211), .B(n212), .Z(n210) );
  AND U12152 ( .A(b[7]), .B(a[120]), .Z(n212) );
  AND U12153 ( .A(b[8]), .B(a[119]), .Z(n211) );
  XOR U12154 ( .A(n213), .B(n214), .Z(n209) );
  XOR U12155 ( .A(n215), .B(n216), .Z(n214) );
  XOR U12156 ( .A(n217), .B(n218), .Z(n216) );
  AND U12157 ( .A(b[13]), .B(a[114]), .Z(n218) );
  AND U12158 ( .A(b[14]), .B(a[113]), .Z(n217) );
  XOR U12159 ( .A(n219), .B(n220), .Z(n215) );
  XOR U12160 ( .A(n221), .B(n222), .Z(n220) );
  XOR U12161 ( .A(n223), .B(n224), .Z(n222) );
  XOR U12162 ( .A(n225), .B(n226), .Z(n224) );
  XOR U12163 ( .A(n227), .B(n228), .Z(n226) );
  XOR U12164 ( .A(n229), .B(n230), .Z(n228) );
  XOR U12165 ( .A(n231), .B(n232), .Z(n230) );
  XOR U12166 ( .A(n233), .B(n234), .Z(n232) );
  XOR U12167 ( .A(n235), .B(n236), .Z(n234) );
  XOR U12168 ( .A(n237), .B(n238), .Z(n236) );
  XOR U12169 ( .A(n239), .B(n240), .Z(n238) );
  XOR U12170 ( .A(n241), .B(n242), .Z(n240) );
  XOR U12171 ( .A(n243), .B(n244), .Z(n242) );
  XOR U12172 ( .A(n245), .B(n246), .Z(n244) );
  XOR U12173 ( .A(n247), .B(n248), .Z(n246) );
  XOR U12174 ( .A(n249), .B(n250), .Z(n248) );
  XOR U12175 ( .A(n251), .B(n252), .Z(n250) );
  XOR U12176 ( .A(n253), .B(n254), .Z(n252) );
  XOR U12177 ( .A(n255), .B(n256), .Z(n254) );
  XOR U12178 ( .A(n257), .B(n258), .Z(n256) );
  XOR U12179 ( .A(n259), .B(n260), .Z(n258) );
  XOR U12180 ( .A(n261), .B(n262), .Z(n260) );
  XOR U12181 ( .A(n263), .B(n264), .Z(n262) );
  XOR U12182 ( .A(n265), .B(n266), .Z(n264) );
  XOR U12183 ( .A(n267), .B(n268), .Z(n266) );
  XOR U12184 ( .A(n269), .B(n270), .Z(n268) );
  XOR U12185 ( .A(n271), .B(n272), .Z(n270) );
  XOR U12186 ( .A(n273), .B(n274), .Z(n272) );
  XOR U12187 ( .A(n275), .B(n276), .Z(n274) );
  XOR U12188 ( .A(n277), .B(n278), .Z(n276) );
  XOR U12189 ( .A(n279), .B(n280), .Z(n278) );
  XOR U12190 ( .A(n281), .B(n282), .Z(n280) );
  XOR U12191 ( .A(n283), .B(n284), .Z(n282) );
  XOR U12192 ( .A(n285), .B(n286), .Z(n284) );
  XOR U12193 ( .A(n287), .B(n288), .Z(n286) );
  XOR U12194 ( .A(n289), .B(n290), .Z(n288) );
  XOR U12195 ( .A(n291), .B(n292), .Z(n290) );
  XOR U12196 ( .A(n293), .B(n294), .Z(n292) );
  XOR U12197 ( .A(n295), .B(n296), .Z(n294) );
  XOR U12198 ( .A(n297), .B(n298), .Z(n296) );
  XOR U12199 ( .A(n299), .B(n300), .Z(n298) );
  XOR U12200 ( .A(n301), .B(n302), .Z(n300) );
  XOR U12201 ( .A(n303), .B(n304), .Z(n302) );
  XOR U12202 ( .A(n305), .B(n306), .Z(n304) );
  XOR U12203 ( .A(n307), .B(n308), .Z(n306) );
  XOR U12204 ( .A(n309), .B(n310), .Z(n308) );
  XOR U12205 ( .A(n311), .B(n312), .Z(n310) );
  XOR U12206 ( .A(n313), .B(n314), .Z(n312) );
  AND U12207 ( .A(b[109]), .B(a[18]), .Z(n314) );
  AND U12208 ( .A(b[115]), .B(a[12]), .Z(n313) );
  XOR U12209 ( .A(n315), .B(n316), .Z(n311) );
  XOR U12210 ( .A(n317), .B(n318), .Z(n316) );
  XOR U12211 ( .A(n319), .B(n320), .Z(n318) );
  XOR U12212 ( .A(n321), .B(n322), .Z(n320) );
  AND U12213 ( .A(b[116]), .B(a[11]), .Z(n322) );
  AND U12214 ( .A(b[121]), .B(a[6]), .Z(n321) );
  XOR U12215 ( .A(n323), .B(n324), .Z(n319) );
  AND U12216 ( .A(b[122]), .B(a[5]), .Z(n324) );
  AND U12217 ( .A(b[123]), .B(a[4]), .Z(n323) );
  XOR U12218 ( .A(n325), .B(n326), .Z(n317) );
  XOR U12219 ( .A(n327), .B(n328), .Z(n326) );
  AND U12220 ( .A(b[124]), .B(a[3]), .Z(n328) );
  AND U12221 ( .A(b[125]), .B(a[2]), .Z(n327) );
  XOR U12222 ( .A(n329), .B(n330), .Z(n325) );
  AND U12223 ( .A(b[126]), .B(a[1]), .Z(n330) );
  AND U12224 ( .A(b[127]), .B(a[0]), .Z(n329) );
  AND U12225 ( .A(b[110]), .B(a[17]), .Z(n315) );
  XOR U12226 ( .A(n331), .B(n332), .Z(n309) );
  XOR U12227 ( .A(n333), .B(n334), .Z(n332) );
  AND U12228 ( .A(b[117]), .B(a[10]), .Z(n334) );
  AND U12229 ( .A(b[118]), .B(a[9]), .Z(n333) );
  XOR U12230 ( .A(n335), .B(n336), .Z(n331) );
  AND U12231 ( .A(b[119]), .B(a[8]), .Z(n336) );
  AND U12232 ( .A(b[120]), .B(a[7]), .Z(n335) );
  AND U12233 ( .A(b[104]), .B(a[23]), .Z(n307) );
  AND U12234 ( .A(b[103]), .B(a[24]), .Z(n305) );
  XOR U12235 ( .A(n337), .B(n338), .Z(n303) );
  XOR U12236 ( .A(n339), .B(n340), .Z(n338) );
  AND U12237 ( .A(b[111]), .B(a[16]), .Z(n340) );
  AND U12238 ( .A(b[112]), .B(a[15]), .Z(n339) );
  XOR U12239 ( .A(n341), .B(n342), .Z(n337) );
  AND U12240 ( .A(b[113]), .B(a[14]), .Z(n342) );
  AND U12241 ( .A(b[114]), .B(a[13]), .Z(n341) );
  AND U12242 ( .A(b[98]), .B(a[29]), .Z(n301) );
  AND U12243 ( .A(b[97]), .B(a[30]), .Z(n299) );
  XOR U12244 ( .A(n343), .B(n344), .Z(n297) );
  XOR U12245 ( .A(n345), .B(n346), .Z(n344) );
  AND U12246 ( .A(b[105]), .B(a[22]), .Z(n346) );
  AND U12247 ( .A(b[106]), .B(a[21]), .Z(n345) );
  XOR U12248 ( .A(n347), .B(n348), .Z(n343) );
  AND U12249 ( .A(b[107]), .B(a[20]), .Z(n348) );
  AND U12250 ( .A(b[108]), .B(a[19]), .Z(n347) );
  AND U12251 ( .A(b[92]), .B(a[35]), .Z(n295) );
  AND U12252 ( .A(b[91]), .B(a[36]), .Z(n293) );
  XOR U12253 ( .A(n349), .B(n350), .Z(n291) );
  XOR U12254 ( .A(n351), .B(n352), .Z(n350) );
  AND U12255 ( .A(b[99]), .B(a[28]), .Z(n352) );
  AND U12256 ( .A(b[100]), .B(a[27]), .Z(n351) );
  XOR U12257 ( .A(n353), .B(n354), .Z(n349) );
  AND U12258 ( .A(b[101]), .B(a[26]), .Z(n354) );
  AND U12259 ( .A(b[102]), .B(a[25]), .Z(n353) );
  AND U12260 ( .A(b[86]), .B(a[41]), .Z(n289) );
  AND U12261 ( .A(b[85]), .B(a[42]), .Z(n287) );
  XOR U12262 ( .A(n355), .B(n356), .Z(n285) );
  XOR U12263 ( .A(n357), .B(n358), .Z(n356) );
  AND U12264 ( .A(b[93]), .B(a[34]), .Z(n358) );
  AND U12265 ( .A(b[94]), .B(a[33]), .Z(n357) );
  XOR U12266 ( .A(n359), .B(n360), .Z(n355) );
  AND U12267 ( .A(b[95]), .B(a[32]), .Z(n360) );
  AND U12268 ( .A(b[96]), .B(a[31]), .Z(n359) );
  AND U12269 ( .A(b[80]), .B(a[47]), .Z(n283) );
  AND U12270 ( .A(b[79]), .B(a[48]), .Z(n281) );
  XOR U12271 ( .A(n361), .B(n362), .Z(n279) );
  XOR U12272 ( .A(n363), .B(n364), .Z(n362) );
  AND U12273 ( .A(b[87]), .B(a[40]), .Z(n364) );
  AND U12274 ( .A(b[88]), .B(a[39]), .Z(n363) );
  XOR U12275 ( .A(n365), .B(n366), .Z(n361) );
  AND U12276 ( .A(b[89]), .B(a[38]), .Z(n366) );
  AND U12277 ( .A(b[90]), .B(a[37]), .Z(n365) );
  AND U12278 ( .A(b[74]), .B(a[53]), .Z(n277) );
  AND U12279 ( .A(b[73]), .B(a[54]), .Z(n275) );
  XOR U12280 ( .A(n367), .B(n368), .Z(n273) );
  XOR U12281 ( .A(n369), .B(n370), .Z(n368) );
  AND U12282 ( .A(b[81]), .B(a[46]), .Z(n370) );
  AND U12283 ( .A(b[82]), .B(a[45]), .Z(n369) );
  XOR U12284 ( .A(n371), .B(n372), .Z(n367) );
  AND U12285 ( .A(b[83]), .B(a[44]), .Z(n372) );
  AND U12286 ( .A(b[84]), .B(a[43]), .Z(n371) );
  AND U12287 ( .A(b[68]), .B(a[59]), .Z(n271) );
  AND U12288 ( .A(b[67]), .B(a[60]), .Z(n269) );
  XOR U12289 ( .A(n373), .B(n374), .Z(n267) );
  XOR U12290 ( .A(n375), .B(n376), .Z(n374) );
  AND U12291 ( .A(b[75]), .B(a[52]), .Z(n376) );
  AND U12292 ( .A(b[76]), .B(a[51]), .Z(n375) );
  XOR U12293 ( .A(n377), .B(n378), .Z(n373) );
  AND U12294 ( .A(b[77]), .B(a[50]), .Z(n378) );
  AND U12295 ( .A(b[78]), .B(a[49]), .Z(n377) );
  AND U12296 ( .A(b[62]), .B(a[65]), .Z(n265) );
  AND U12297 ( .A(b[61]), .B(a[66]), .Z(n263) );
  XOR U12298 ( .A(n379), .B(n380), .Z(n261) );
  XOR U12299 ( .A(n381), .B(n382), .Z(n380) );
  AND U12300 ( .A(b[69]), .B(a[58]), .Z(n382) );
  AND U12301 ( .A(b[70]), .B(a[57]), .Z(n381) );
  XOR U12302 ( .A(n383), .B(n384), .Z(n379) );
  AND U12303 ( .A(b[71]), .B(a[56]), .Z(n384) );
  AND U12304 ( .A(b[72]), .B(a[55]), .Z(n383) );
  AND U12305 ( .A(b[56]), .B(a[71]), .Z(n259) );
  AND U12306 ( .A(b[55]), .B(a[72]), .Z(n257) );
  XOR U12307 ( .A(n385), .B(n386), .Z(n255) );
  XOR U12308 ( .A(n387), .B(n388), .Z(n386) );
  AND U12309 ( .A(b[63]), .B(a[64]), .Z(n388) );
  AND U12310 ( .A(b[64]), .B(a[63]), .Z(n387) );
  XOR U12311 ( .A(n389), .B(n390), .Z(n385) );
  AND U12312 ( .A(b[65]), .B(a[62]), .Z(n390) );
  AND U12313 ( .A(b[66]), .B(a[61]), .Z(n389) );
  AND U12314 ( .A(b[50]), .B(a[77]), .Z(n253) );
  AND U12315 ( .A(b[49]), .B(a[78]), .Z(n251) );
  XOR U12316 ( .A(n391), .B(n392), .Z(n249) );
  XOR U12317 ( .A(n393), .B(n394), .Z(n392) );
  AND U12318 ( .A(b[57]), .B(a[70]), .Z(n394) );
  AND U12319 ( .A(b[58]), .B(a[69]), .Z(n393) );
  XOR U12320 ( .A(n395), .B(n396), .Z(n391) );
  AND U12321 ( .A(b[59]), .B(a[68]), .Z(n396) );
  AND U12322 ( .A(b[60]), .B(a[67]), .Z(n395) );
  AND U12323 ( .A(b[44]), .B(a[83]), .Z(n247) );
  AND U12324 ( .A(b[43]), .B(a[84]), .Z(n245) );
  XOR U12325 ( .A(n397), .B(n398), .Z(n243) );
  XOR U12326 ( .A(n399), .B(n400), .Z(n398) );
  AND U12327 ( .A(b[51]), .B(a[76]), .Z(n400) );
  AND U12328 ( .A(b[52]), .B(a[75]), .Z(n399) );
  XOR U12329 ( .A(n401), .B(n402), .Z(n397) );
  AND U12330 ( .A(b[53]), .B(a[74]), .Z(n402) );
  AND U12331 ( .A(b[54]), .B(a[73]), .Z(n401) );
  AND U12332 ( .A(b[38]), .B(a[89]), .Z(n241) );
  AND U12333 ( .A(b[37]), .B(a[90]), .Z(n239) );
  XOR U12334 ( .A(n403), .B(n404), .Z(n237) );
  XOR U12335 ( .A(n405), .B(n406), .Z(n404) );
  AND U12336 ( .A(b[45]), .B(a[82]), .Z(n406) );
  AND U12337 ( .A(b[46]), .B(a[81]), .Z(n405) );
  XOR U12338 ( .A(n407), .B(n408), .Z(n403) );
  AND U12339 ( .A(b[47]), .B(a[80]), .Z(n408) );
  AND U12340 ( .A(b[48]), .B(a[79]), .Z(n407) );
  AND U12341 ( .A(b[32]), .B(a[95]), .Z(n235) );
  AND U12342 ( .A(b[31]), .B(a[96]), .Z(n233) );
  XOR U12343 ( .A(n409), .B(n410), .Z(n231) );
  XOR U12344 ( .A(n411), .B(n412), .Z(n410) );
  AND U12345 ( .A(b[39]), .B(a[88]), .Z(n412) );
  AND U12346 ( .A(b[40]), .B(a[87]), .Z(n411) );
  XOR U12347 ( .A(n413), .B(n414), .Z(n409) );
  AND U12348 ( .A(b[41]), .B(a[86]), .Z(n414) );
  AND U12349 ( .A(b[42]), .B(a[85]), .Z(n413) );
  AND U12350 ( .A(b[26]), .B(a[101]), .Z(n229) );
  AND U12351 ( .A(b[25]), .B(a[102]), .Z(n227) );
  XOR U12352 ( .A(n415), .B(n416), .Z(n225) );
  XOR U12353 ( .A(n417), .B(n418), .Z(n416) );
  AND U12354 ( .A(b[33]), .B(a[94]), .Z(n418) );
  AND U12355 ( .A(b[34]), .B(a[93]), .Z(n417) );
  XOR U12356 ( .A(n419), .B(n420), .Z(n415) );
  AND U12357 ( .A(b[35]), .B(a[92]), .Z(n420) );
  AND U12358 ( .A(b[36]), .B(a[91]), .Z(n419) );
  AND U12359 ( .A(b[20]), .B(a[107]), .Z(n223) );
  AND U12360 ( .A(b[19]), .B(a[108]), .Z(n221) );
  XOR U12361 ( .A(n421), .B(n422), .Z(n219) );
  XOR U12362 ( .A(n423), .B(n424), .Z(n422) );
  AND U12363 ( .A(b[27]), .B(a[100]), .Z(n424) );
  AND U12364 ( .A(b[28]), .B(a[99]), .Z(n423) );
  XOR U12365 ( .A(n425), .B(n426), .Z(n421) );
  AND U12366 ( .A(b[29]), .B(a[98]), .Z(n426) );
  AND U12367 ( .A(b[30]), .B(a[97]), .Z(n425) );
  XOR U12368 ( .A(n427), .B(n428), .Z(n213) );
  XOR U12369 ( .A(n429), .B(n430), .Z(n428) );
  AND U12370 ( .A(b[21]), .B(a[106]), .Z(n430) );
  AND U12371 ( .A(b[22]), .B(a[105]), .Z(n429) );
  XOR U12372 ( .A(n431), .B(n432), .Z(n427) );
  AND U12373 ( .A(b[23]), .B(a[104]), .Z(n432) );
  AND U12374 ( .A(b[24]), .B(a[103]), .Z(n431) );
  XOR U12375 ( .A(n433), .B(n434), .Z(n207) );
  XOR U12376 ( .A(n435), .B(n436), .Z(n434) );
  AND U12377 ( .A(b[15]), .B(a[112]), .Z(n436) );
  AND U12378 ( .A(b[16]), .B(a[111]), .Z(n435) );
  XOR U12379 ( .A(n437), .B(n438), .Z(n433) );
  AND U12380 ( .A(b[17]), .B(a[110]), .Z(n438) );
  AND U12381 ( .A(b[18]), .B(a[109]), .Z(n437) );
  XOR U12382 ( .A(n439), .B(n440), .Z(n201) );
  XOR U12383 ( .A(n441), .B(n442), .Z(n440) );
  AND U12384 ( .A(b[9]), .B(a[118]), .Z(n442) );
  AND U12385 ( .A(b[10]), .B(a[117]), .Z(n441) );
  XOR U12386 ( .A(n443), .B(n444), .Z(n439) );
  AND U12387 ( .A(b[11]), .B(a[116]), .Z(n444) );
  AND U12388 ( .A(b[12]), .B(a[115]), .Z(n443) );
  AND U12389 ( .A(a[127]), .B(b[0]), .Z(n199) );
  XNOR U12390 ( .A(n445), .B(n205), .Z(n197) );
  OR U12391 ( .A(n446), .B(n447), .Z(n205) );
  AND U12392 ( .A(b[2]), .B(a[125]), .Z(n445) );
  XOR U12393 ( .A(n448), .B(n449), .Z(n195) );
  XOR U12394 ( .A(n450), .B(n451), .Z(n449) );
  AND U12395 ( .A(b[3]), .B(a[124]), .Z(n451) );
  AND U12396 ( .A(b[4]), .B(a[123]), .Z(n450) );
  XOR U12397 ( .A(n452), .B(n453), .Z(n448) );
  AND U12398 ( .A(b[5]), .B(a[122]), .Z(n453) );
  AND U12399 ( .A(b[6]), .B(a[121]), .Z(n452) );
  XOR U12400 ( .A(n446), .B(n447), .Z(c[126]) );
  XOR U12401 ( .A(n454), .B(n455), .Z(n447) );
  XNOR U12402 ( .A(n456), .B(n457), .Z(n455) );
  XOR U12403 ( .A(n458), .B(n459), .Z(n457) );
  XOR U12404 ( .A(n460), .B(n461), .Z(n459) );
  XNOR U12405 ( .A(n462), .B(n456), .Z(n461) );
  XOR U12406 ( .A(n463), .B(n464), .Z(n460) );
  XOR U12407 ( .A(n465), .B(n466), .Z(n464) );
  XOR U12408 ( .A(n467), .B(n468), .Z(n466) );
  XOR U12409 ( .A(n469), .B(n470), .Z(n468) );
  AND U12410 ( .A(b[7]), .B(a[119]), .Z(n469) );
  XOR U12411 ( .A(n471), .B(n472), .Z(n467) );
  XOR U12412 ( .A(n473), .B(n474), .Z(n472) );
  XOR U12413 ( .A(n475), .B(n476), .Z(n474) );
  XOR U12414 ( .A(n477), .B(n478), .Z(n476) );
  AND U12415 ( .A(b[13]), .B(a[113]), .Z(n477) );
  XOR U12416 ( .A(n479), .B(n480), .Z(n475) );
  AND U12417 ( .A(b[18]), .B(a[108]), .Z(n479) );
  XOR U12418 ( .A(n478), .B(n481), .Z(n473) );
  XOR U12419 ( .A(n480), .B(n482), .Z(n481) );
  XOR U12420 ( .A(n483), .B(n484), .Z(n482) );
  XOR U12421 ( .A(n485), .B(n486), .Z(n484) );
  XOR U12422 ( .A(n487), .B(n488), .Z(n486) );
  XOR U12423 ( .A(n489), .B(n490), .Z(n488) );
  AND U12424 ( .A(b[19]), .B(a[107]), .Z(n489) );
  XOR U12425 ( .A(n491), .B(n492), .Z(n487) );
  AND U12426 ( .A(b[24]), .B(a[102]), .Z(n491) );
  XOR U12427 ( .A(n490), .B(n493), .Z(n485) );
  XOR U12428 ( .A(n492), .B(n494), .Z(n493) );
  XOR U12429 ( .A(n495), .B(n496), .Z(n494) );
  XOR U12430 ( .A(n497), .B(n498), .Z(n496) );
  XOR U12431 ( .A(n499), .B(n500), .Z(n498) );
  XOR U12432 ( .A(n501), .B(n502), .Z(n500) );
  AND U12433 ( .A(b[25]), .B(a[101]), .Z(n501) );
  XOR U12434 ( .A(n503), .B(n504), .Z(n499) );
  AND U12435 ( .A(a[96]), .B(b[30]), .Z(n503) );
  XOR U12436 ( .A(n502), .B(n505), .Z(n497) );
  XOR U12437 ( .A(n504), .B(n506), .Z(n505) );
  XOR U12438 ( .A(n507), .B(n508), .Z(n506) );
  XOR U12439 ( .A(n509), .B(n510), .Z(n508) );
  XOR U12440 ( .A(n511), .B(n512), .Z(n510) );
  XOR U12441 ( .A(n513), .B(n514), .Z(n512) );
  AND U12442 ( .A(a[95]), .B(b[31]), .Z(n513) );
  XOR U12443 ( .A(n515), .B(n516), .Z(n511) );
  AND U12444 ( .A(a[90]), .B(b[36]), .Z(n515) );
  XOR U12445 ( .A(n514), .B(n517), .Z(n509) );
  XOR U12446 ( .A(n516), .B(n518), .Z(n517) );
  XOR U12447 ( .A(n519), .B(n520), .Z(n518) );
  XOR U12448 ( .A(n521), .B(n522), .Z(n520) );
  XOR U12449 ( .A(n523), .B(n524), .Z(n522) );
  XOR U12450 ( .A(n525), .B(n526), .Z(n524) );
  AND U12451 ( .A(a[89]), .B(b[37]), .Z(n525) );
  XOR U12452 ( .A(n527), .B(n528), .Z(n523) );
  AND U12453 ( .A(a[84]), .B(b[42]), .Z(n527) );
  XOR U12454 ( .A(n526), .B(n529), .Z(n521) );
  XOR U12455 ( .A(n528), .B(n530), .Z(n529) );
  XOR U12456 ( .A(n531), .B(n532), .Z(n530) );
  XOR U12457 ( .A(n533), .B(n534), .Z(n532) );
  XOR U12458 ( .A(n535), .B(n536), .Z(n534) );
  XOR U12459 ( .A(n537), .B(n538), .Z(n536) );
  AND U12460 ( .A(a[83]), .B(b[43]), .Z(n537) );
  XOR U12461 ( .A(n539), .B(n540), .Z(n535) );
  AND U12462 ( .A(a[78]), .B(b[48]), .Z(n539) );
  XOR U12463 ( .A(n538), .B(n541), .Z(n533) );
  XOR U12464 ( .A(n540), .B(n542), .Z(n541) );
  XOR U12465 ( .A(n543), .B(n544), .Z(n542) );
  XOR U12466 ( .A(n545), .B(n546), .Z(n544) );
  XOR U12467 ( .A(n547), .B(n548), .Z(n546) );
  XOR U12468 ( .A(n549), .B(n550), .Z(n548) );
  AND U12469 ( .A(a[77]), .B(b[49]), .Z(n549) );
  XOR U12470 ( .A(n551), .B(n552), .Z(n547) );
  AND U12471 ( .A(a[72]), .B(b[54]), .Z(n551) );
  XOR U12472 ( .A(n550), .B(n553), .Z(n545) );
  XOR U12473 ( .A(n552), .B(n554), .Z(n553) );
  XOR U12474 ( .A(n555), .B(n556), .Z(n554) );
  XOR U12475 ( .A(n557), .B(n558), .Z(n556) );
  XOR U12476 ( .A(n559), .B(n560), .Z(n558) );
  XOR U12477 ( .A(n561), .B(n562), .Z(n560) );
  AND U12478 ( .A(a[71]), .B(b[55]), .Z(n561) );
  XOR U12479 ( .A(n563), .B(n564), .Z(n559) );
  AND U12480 ( .A(a[66]), .B(b[60]), .Z(n563) );
  XOR U12481 ( .A(n562), .B(n565), .Z(n557) );
  XOR U12482 ( .A(n564), .B(n566), .Z(n565) );
  XOR U12483 ( .A(n567), .B(n568), .Z(n566) );
  XOR U12484 ( .A(n569), .B(n570), .Z(n568) );
  XOR U12485 ( .A(n571), .B(n572), .Z(n570) );
  XOR U12486 ( .A(n573), .B(n574), .Z(n572) );
  AND U12487 ( .A(a[65]), .B(b[61]), .Z(n573) );
  XOR U12488 ( .A(n575), .B(n576), .Z(n571) );
  AND U12489 ( .A(a[60]), .B(b[66]), .Z(n575) );
  XOR U12490 ( .A(n574), .B(n577), .Z(n569) );
  XOR U12491 ( .A(n576), .B(n578), .Z(n577) );
  XOR U12492 ( .A(n579), .B(n580), .Z(n578) );
  XOR U12493 ( .A(n581), .B(n582), .Z(n580) );
  XOR U12494 ( .A(n583), .B(n584), .Z(n582) );
  XOR U12495 ( .A(n585), .B(n586), .Z(n584) );
  AND U12496 ( .A(a[59]), .B(b[67]), .Z(n585) );
  XOR U12497 ( .A(n587), .B(n588), .Z(n583) );
  AND U12498 ( .A(a[54]), .B(b[72]), .Z(n587) );
  XOR U12499 ( .A(n586), .B(n589), .Z(n581) );
  XOR U12500 ( .A(n588), .B(n590), .Z(n589) );
  XOR U12501 ( .A(n591), .B(n592), .Z(n590) );
  XOR U12502 ( .A(n593), .B(n594), .Z(n592) );
  XOR U12503 ( .A(n595), .B(n596), .Z(n594) );
  XOR U12504 ( .A(n597), .B(n598), .Z(n596) );
  AND U12505 ( .A(a[53]), .B(b[73]), .Z(n597) );
  XOR U12506 ( .A(n599), .B(n600), .Z(n595) );
  AND U12507 ( .A(a[48]), .B(b[78]), .Z(n599) );
  XOR U12508 ( .A(n598), .B(n601), .Z(n593) );
  XOR U12509 ( .A(n600), .B(n602), .Z(n601) );
  XOR U12510 ( .A(n603), .B(n604), .Z(n602) );
  XOR U12511 ( .A(n605), .B(n606), .Z(n604) );
  XOR U12512 ( .A(n607), .B(n608), .Z(n606) );
  XOR U12513 ( .A(n609), .B(n610), .Z(n608) );
  AND U12514 ( .A(a[47]), .B(b[79]), .Z(n609) );
  XOR U12515 ( .A(n611), .B(n612), .Z(n607) );
  AND U12516 ( .A(a[42]), .B(b[84]), .Z(n611) );
  XOR U12517 ( .A(n610), .B(n613), .Z(n605) );
  XOR U12518 ( .A(n612), .B(n614), .Z(n613) );
  XOR U12519 ( .A(n615), .B(n616), .Z(n614) );
  XOR U12520 ( .A(n617), .B(n618), .Z(n616) );
  XOR U12521 ( .A(n619), .B(n620), .Z(n618) );
  XOR U12522 ( .A(n621), .B(n622), .Z(n620) );
  AND U12523 ( .A(a[41]), .B(b[85]), .Z(n621) );
  XOR U12524 ( .A(n623), .B(n624), .Z(n619) );
  AND U12525 ( .A(a[36]), .B(b[90]), .Z(n623) );
  XOR U12526 ( .A(n622), .B(n625), .Z(n617) );
  XOR U12527 ( .A(n624), .B(n626), .Z(n625) );
  XOR U12528 ( .A(n627), .B(n628), .Z(n626) );
  XOR U12529 ( .A(n629), .B(n630), .Z(n628) );
  XOR U12530 ( .A(n631), .B(n632), .Z(n630) );
  XOR U12531 ( .A(n633), .B(n634), .Z(n632) );
  AND U12532 ( .A(a[35]), .B(b[91]), .Z(n633) );
  XOR U12533 ( .A(n635), .B(n636), .Z(n631) );
  AND U12534 ( .A(a[30]), .B(b[96]), .Z(n635) );
  XOR U12535 ( .A(n634), .B(n637), .Z(n629) );
  XOR U12536 ( .A(n636), .B(n638), .Z(n637) );
  XOR U12537 ( .A(n639), .B(n640), .Z(n638) );
  XOR U12538 ( .A(n641), .B(n642), .Z(n640) );
  XOR U12539 ( .A(n643), .B(n644), .Z(n642) );
  XOR U12540 ( .A(n645), .B(n646), .Z(n644) );
  AND U12541 ( .A(a[29]), .B(b[97]), .Z(n645) );
  XOR U12542 ( .A(n647), .B(n648), .Z(n643) );
  AND U12543 ( .A(a[24]), .B(b[102]), .Z(n647) );
  XOR U12544 ( .A(n646), .B(n649), .Z(n641) );
  XOR U12545 ( .A(n648), .B(n650), .Z(n649) );
  XOR U12546 ( .A(n651), .B(n652), .Z(n650) );
  XOR U12547 ( .A(n653), .B(n654), .Z(n652) );
  XOR U12548 ( .A(n655), .B(n656), .Z(n654) );
  XOR U12549 ( .A(n657), .B(n658), .Z(n656) );
  AND U12550 ( .A(a[23]), .B(b[103]), .Z(n657) );
  XOR U12551 ( .A(n659), .B(n660), .Z(n655) );
  AND U12552 ( .A(a[18]), .B(b[108]), .Z(n659) );
  XOR U12553 ( .A(n658), .B(n661), .Z(n653) );
  XOR U12554 ( .A(n660), .B(n662), .Z(n661) );
  XOR U12555 ( .A(n663), .B(n664), .Z(n662) );
  XOR U12556 ( .A(n665), .B(n666), .Z(n664) );
  XOR U12557 ( .A(n667), .B(n668), .Z(n666) );
  XOR U12558 ( .A(n669), .B(n670), .Z(n668) );
  AND U12559 ( .A(a[17]), .B(b[109]), .Z(n669) );
  XOR U12560 ( .A(n671), .B(n672), .Z(n667) );
  AND U12561 ( .A(a[12]), .B(b[114]), .Z(n671) );
  XOR U12562 ( .A(n670), .B(n673), .Z(n665) );
  XOR U12563 ( .A(n672), .B(n674), .Z(n673) );
  XOR U12564 ( .A(n675), .B(n676), .Z(n674) );
  XOR U12565 ( .A(n677), .B(n678), .Z(n676) );
  XOR U12566 ( .A(n679), .B(n680), .Z(n678) );
  XOR U12567 ( .A(n681), .B(n682), .Z(n680) );
  AND U12568 ( .A(a[11]), .B(b[115]), .Z(n681) );
  XOR U12569 ( .A(n683), .B(n684), .Z(n679) );
  AND U12570 ( .A(a[6]), .B(b[120]), .Z(n683) );
  XOR U12571 ( .A(n682), .B(n685), .Z(n677) );
  XOR U12572 ( .A(n686), .B(n687), .Z(n685) );
  XOR U12573 ( .A(n684), .B(n688), .Z(n687) );
  XOR U12574 ( .A(n689), .B(n690), .Z(n688) );
  AND U12575 ( .A(a[5]), .B(b[121]), .Z(n690) );
  AND U12576 ( .A(a[4]), .B(b[122]), .Z(n689) );
  XOR U12577 ( .A(n691), .B(n692), .Z(n684) );
  ANDN U12578 ( .B(n693), .A(n694), .Z(n691) );
  XOR U12579 ( .A(n695), .B(n696), .Z(n686) );
  XOR U12580 ( .A(n697), .B(n698), .Z(n696) );
  AND U12581 ( .A(a[3]), .B(b[123]), .Z(n698) );
  AND U12582 ( .A(a[2]), .B(b[124]), .Z(n697) );
  XOR U12583 ( .A(n699), .B(n700), .Z(n695) );
  AND U12584 ( .A(a[1]), .B(b[125]), .Z(n700) );
  AND U12585 ( .A(a[0]), .B(b[126]), .Z(n699) );
  XOR U12586 ( .A(n701), .B(n702), .Z(n682) );
  NOR U12587 ( .A(n703), .B(n704), .Z(n701) );
  XOR U12588 ( .A(n705), .B(n706), .Z(n675) );
  XOR U12589 ( .A(n707), .B(n708), .Z(n706) );
  AND U12590 ( .A(a[10]), .B(b[116]), .Z(n708) );
  AND U12591 ( .A(a[9]), .B(b[117]), .Z(n707) );
  XOR U12592 ( .A(n709), .B(n710), .Z(n705) );
  AND U12593 ( .A(a[8]), .B(b[118]), .Z(n710) );
  AND U12594 ( .A(a[7]), .B(b[119]), .Z(n709) );
  XOR U12595 ( .A(n711), .B(n712), .Z(n672) );
  AND U12596 ( .A(n713), .B(n714), .Z(n711) );
  XOR U12597 ( .A(n715), .B(n716), .Z(n670) );
  NOR U12598 ( .A(n717), .B(n718), .Z(n715) );
  XOR U12599 ( .A(n719), .B(n720), .Z(n663) );
  XOR U12600 ( .A(n721), .B(n722), .Z(n720) );
  AND U12601 ( .A(a[16]), .B(b[110]), .Z(n722) );
  AND U12602 ( .A(a[15]), .B(b[111]), .Z(n721) );
  XOR U12603 ( .A(n723), .B(n724), .Z(n719) );
  AND U12604 ( .A(a[14]), .B(b[112]), .Z(n724) );
  AND U12605 ( .A(a[13]), .B(b[113]), .Z(n723) );
  XOR U12606 ( .A(n725), .B(n726), .Z(n660) );
  AND U12607 ( .A(n727), .B(n728), .Z(n725) );
  XOR U12608 ( .A(n729), .B(n730), .Z(n658) );
  NOR U12609 ( .A(n731), .B(n732), .Z(n729) );
  XOR U12610 ( .A(n733), .B(n734), .Z(n651) );
  XOR U12611 ( .A(n735), .B(n736), .Z(n734) );
  AND U12612 ( .A(a[22]), .B(b[104]), .Z(n736) );
  AND U12613 ( .A(a[21]), .B(b[105]), .Z(n735) );
  XOR U12614 ( .A(n737), .B(n738), .Z(n733) );
  AND U12615 ( .A(a[20]), .B(b[106]), .Z(n738) );
  AND U12616 ( .A(a[19]), .B(b[107]), .Z(n737) );
  XOR U12617 ( .A(n739), .B(n740), .Z(n648) );
  AND U12618 ( .A(n741), .B(n742), .Z(n739) );
  XOR U12619 ( .A(n743), .B(n744), .Z(n646) );
  NOR U12620 ( .A(n745), .B(n746), .Z(n743) );
  XOR U12621 ( .A(n747), .B(n748), .Z(n639) );
  XOR U12622 ( .A(n749), .B(n750), .Z(n748) );
  AND U12623 ( .A(a[28]), .B(b[98]), .Z(n750) );
  AND U12624 ( .A(a[27]), .B(b[99]), .Z(n749) );
  XOR U12625 ( .A(n751), .B(n752), .Z(n747) );
  AND U12626 ( .A(a[26]), .B(b[100]), .Z(n752) );
  AND U12627 ( .A(a[25]), .B(b[101]), .Z(n751) );
  XOR U12628 ( .A(n753), .B(n754), .Z(n636) );
  AND U12629 ( .A(n755), .B(n756), .Z(n753) );
  XOR U12630 ( .A(n757), .B(n758), .Z(n634) );
  NOR U12631 ( .A(n759), .B(n760), .Z(n757) );
  XOR U12632 ( .A(n761), .B(n762), .Z(n627) );
  XOR U12633 ( .A(n763), .B(n764), .Z(n762) );
  AND U12634 ( .A(a[34]), .B(b[92]), .Z(n764) );
  AND U12635 ( .A(a[33]), .B(b[93]), .Z(n763) );
  XOR U12636 ( .A(n765), .B(n766), .Z(n761) );
  AND U12637 ( .A(a[32]), .B(b[94]), .Z(n766) );
  AND U12638 ( .A(a[31]), .B(b[95]), .Z(n765) );
  XOR U12639 ( .A(n767), .B(n768), .Z(n624) );
  AND U12640 ( .A(n769), .B(n770), .Z(n767) );
  XOR U12641 ( .A(n771), .B(n772), .Z(n622) );
  NOR U12642 ( .A(n773), .B(n774), .Z(n771) );
  XOR U12643 ( .A(n775), .B(n776), .Z(n615) );
  XOR U12644 ( .A(n777), .B(n778), .Z(n776) );
  AND U12645 ( .A(a[40]), .B(b[86]), .Z(n778) );
  AND U12646 ( .A(a[39]), .B(b[87]), .Z(n777) );
  XOR U12647 ( .A(n779), .B(n780), .Z(n775) );
  AND U12648 ( .A(a[38]), .B(b[88]), .Z(n780) );
  AND U12649 ( .A(a[37]), .B(b[89]), .Z(n779) );
  XOR U12650 ( .A(n781), .B(n782), .Z(n612) );
  AND U12651 ( .A(n783), .B(n784), .Z(n781) );
  XOR U12652 ( .A(n785), .B(n786), .Z(n610) );
  NOR U12653 ( .A(n787), .B(n788), .Z(n785) );
  XOR U12654 ( .A(n789), .B(n790), .Z(n603) );
  XOR U12655 ( .A(n791), .B(n792), .Z(n790) );
  AND U12656 ( .A(a[46]), .B(b[80]), .Z(n792) );
  AND U12657 ( .A(a[45]), .B(b[81]), .Z(n791) );
  XOR U12658 ( .A(n793), .B(n794), .Z(n789) );
  AND U12659 ( .A(a[44]), .B(b[82]), .Z(n794) );
  AND U12660 ( .A(a[43]), .B(b[83]), .Z(n793) );
  XOR U12661 ( .A(n795), .B(n796), .Z(n600) );
  AND U12662 ( .A(n797), .B(n798), .Z(n795) );
  XOR U12663 ( .A(n799), .B(n800), .Z(n598) );
  NOR U12664 ( .A(n801), .B(n802), .Z(n799) );
  XOR U12665 ( .A(n803), .B(n804), .Z(n591) );
  XOR U12666 ( .A(n805), .B(n806), .Z(n804) );
  AND U12667 ( .A(a[52]), .B(b[74]), .Z(n806) );
  AND U12668 ( .A(a[51]), .B(b[75]), .Z(n805) );
  XOR U12669 ( .A(n807), .B(n808), .Z(n803) );
  AND U12670 ( .A(a[50]), .B(b[76]), .Z(n808) );
  AND U12671 ( .A(a[49]), .B(b[77]), .Z(n807) );
  XOR U12672 ( .A(n809), .B(n810), .Z(n588) );
  AND U12673 ( .A(n811), .B(n812), .Z(n809) );
  XOR U12674 ( .A(n813), .B(n814), .Z(n586) );
  NOR U12675 ( .A(n815), .B(n816), .Z(n813) );
  XOR U12676 ( .A(n817), .B(n818), .Z(n579) );
  XOR U12677 ( .A(n819), .B(n820), .Z(n818) );
  AND U12678 ( .A(a[58]), .B(b[68]), .Z(n820) );
  AND U12679 ( .A(a[57]), .B(b[69]), .Z(n819) );
  XOR U12680 ( .A(n821), .B(n822), .Z(n817) );
  AND U12681 ( .A(a[56]), .B(b[70]), .Z(n822) );
  AND U12682 ( .A(a[55]), .B(b[71]), .Z(n821) );
  XOR U12683 ( .A(n823), .B(n824), .Z(n576) );
  AND U12684 ( .A(n825), .B(n826), .Z(n823) );
  XOR U12685 ( .A(n827), .B(n828), .Z(n574) );
  NOR U12686 ( .A(n829), .B(n830), .Z(n827) );
  XOR U12687 ( .A(n831), .B(n832), .Z(n567) );
  XOR U12688 ( .A(n833), .B(n834), .Z(n832) );
  AND U12689 ( .A(a[64]), .B(b[62]), .Z(n834) );
  AND U12690 ( .A(a[63]), .B(b[63]), .Z(n833) );
  XOR U12691 ( .A(n835), .B(n836), .Z(n831) );
  AND U12692 ( .A(a[62]), .B(b[64]), .Z(n836) );
  AND U12693 ( .A(a[61]), .B(b[65]), .Z(n835) );
  XOR U12694 ( .A(n837), .B(n838), .Z(n564) );
  AND U12695 ( .A(n839), .B(n840), .Z(n837) );
  XOR U12696 ( .A(n841), .B(n842), .Z(n562) );
  NOR U12697 ( .A(n843), .B(n844), .Z(n841) );
  XOR U12698 ( .A(n845), .B(n846), .Z(n555) );
  XOR U12699 ( .A(n847), .B(n848), .Z(n846) );
  AND U12700 ( .A(a[70]), .B(b[56]), .Z(n848) );
  AND U12701 ( .A(a[69]), .B(b[57]), .Z(n847) );
  XOR U12702 ( .A(n849), .B(n850), .Z(n845) );
  AND U12703 ( .A(a[68]), .B(b[58]), .Z(n850) );
  AND U12704 ( .A(a[67]), .B(b[59]), .Z(n849) );
  XOR U12705 ( .A(n851), .B(n852), .Z(n552) );
  AND U12706 ( .A(n853), .B(n854), .Z(n851) );
  XOR U12707 ( .A(n855), .B(n856), .Z(n550) );
  NOR U12708 ( .A(n857), .B(n858), .Z(n855) );
  XOR U12709 ( .A(n859), .B(n860), .Z(n543) );
  XOR U12710 ( .A(n861), .B(n862), .Z(n860) );
  AND U12711 ( .A(a[76]), .B(b[50]), .Z(n862) );
  AND U12712 ( .A(a[75]), .B(b[51]), .Z(n861) );
  XOR U12713 ( .A(n863), .B(n864), .Z(n859) );
  AND U12714 ( .A(a[74]), .B(b[52]), .Z(n864) );
  AND U12715 ( .A(a[73]), .B(b[53]), .Z(n863) );
  XOR U12716 ( .A(n865), .B(n866), .Z(n540) );
  AND U12717 ( .A(n867), .B(n868), .Z(n865) );
  XOR U12718 ( .A(n869), .B(n870), .Z(n538) );
  NOR U12719 ( .A(n871), .B(n872), .Z(n869) );
  XOR U12720 ( .A(n873), .B(n874), .Z(n531) );
  XOR U12721 ( .A(n875), .B(n876), .Z(n874) );
  AND U12722 ( .A(a[82]), .B(b[44]), .Z(n876) );
  AND U12723 ( .A(a[81]), .B(b[45]), .Z(n875) );
  XOR U12724 ( .A(n877), .B(n878), .Z(n873) );
  AND U12725 ( .A(a[80]), .B(b[46]), .Z(n878) );
  AND U12726 ( .A(a[79]), .B(b[47]), .Z(n877) );
  XOR U12727 ( .A(n879), .B(n880), .Z(n528) );
  AND U12728 ( .A(n881), .B(n882), .Z(n879) );
  XOR U12729 ( .A(n883), .B(n884), .Z(n526) );
  NOR U12730 ( .A(n885), .B(n886), .Z(n883) );
  XOR U12731 ( .A(n887), .B(n888), .Z(n519) );
  XOR U12732 ( .A(n889), .B(n890), .Z(n888) );
  AND U12733 ( .A(a[88]), .B(b[38]), .Z(n890) );
  AND U12734 ( .A(a[87]), .B(b[39]), .Z(n889) );
  XOR U12735 ( .A(n891), .B(n892), .Z(n887) );
  AND U12736 ( .A(a[86]), .B(b[40]), .Z(n892) );
  AND U12737 ( .A(a[85]), .B(b[41]), .Z(n891) );
  XOR U12738 ( .A(n893), .B(n894), .Z(n516) );
  AND U12739 ( .A(n895), .B(n896), .Z(n893) );
  XOR U12740 ( .A(n897), .B(n898), .Z(n514) );
  NOR U12741 ( .A(n899), .B(n900), .Z(n897) );
  XOR U12742 ( .A(n901), .B(n902), .Z(n507) );
  XOR U12743 ( .A(n903), .B(n904), .Z(n902) );
  AND U12744 ( .A(a[94]), .B(b[32]), .Z(n904) );
  AND U12745 ( .A(a[93]), .B(b[33]), .Z(n903) );
  XOR U12746 ( .A(n905), .B(n906), .Z(n901) );
  AND U12747 ( .A(a[92]), .B(b[34]), .Z(n906) );
  AND U12748 ( .A(a[91]), .B(b[35]), .Z(n905) );
  XOR U12749 ( .A(n907), .B(n908), .Z(n504) );
  AND U12750 ( .A(n909), .B(n910), .Z(n907) );
  XOR U12751 ( .A(n911), .B(n912), .Z(n502) );
  NOR U12752 ( .A(n913), .B(n914), .Z(n911) );
  XOR U12753 ( .A(n915), .B(n916), .Z(n495) );
  XOR U12754 ( .A(n917), .B(n918), .Z(n916) );
  AND U12755 ( .A(b[26]), .B(a[100]), .Z(n918) );
  AND U12756 ( .A(a[99]), .B(b[27]), .Z(n917) );
  XOR U12757 ( .A(n919), .B(n920), .Z(n915) );
  AND U12758 ( .A(a[98]), .B(b[28]), .Z(n920) );
  AND U12759 ( .A(a[97]), .B(b[29]), .Z(n919) );
  XOR U12760 ( .A(n921), .B(n922), .Z(n492) );
  AND U12761 ( .A(n923), .B(n924), .Z(n921) );
  XOR U12762 ( .A(n925), .B(n926), .Z(n490) );
  NOR U12763 ( .A(n927), .B(n928), .Z(n925) );
  XOR U12764 ( .A(n929), .B(n930), .Z(n483) );
  XOR U12765 ( .A(n931), .B(n932), .Z(n930) );
  AND U12766 ( .A(b[20]), .B(a[106]), .Z(n932) );
  AND U12767 ( .A(b[21]), .B(a[105]), .Z(n931) );
  XOR U12768 ( .A(n933), .B(n934), .Z(n929) );
  AND U12769 ( .A(b[22]), .B(a[104]), .Z(n934) );
  AND U12770 ( .A(b[23]), .B(a[103]), .Z(n933) );
  XOR U12771 ( .A(n935), .B(n936), .Z(n480) );
  AND U12772 ( .A(n937), .B(n938), .Z(n935) );
  XOR U12773 ( .A(n939), .B(n940), .Z(n478) );
  ANDN U12774 ( .B(n941), .A(n942), .Z(n939) );
  XOR U12775 ( .A(n943), .B(n944), .Z(n471) );
  XOR U12776 ( .A(n945), .B(n946), .Z(n944) );
  AND U12777 ( .A(b[14]), .B(a[112]), .Z(n946) );
  AND U12778 ( .A(b[15]), .B(a[111]), .Z(n945) );
  XOR U12779 ( .A(n947), .B(n948), .Z(n943) );
  AND U12780 ( .A(b[16]), .B(a[110]), .Z(n948) );
  AND U12781 ( .A(b[17]), .B(a[109]), .Z(n947) );
  XOR U12782 ( .A(n949), .B(n470), .Z(n465) );
  XOR U12783 ( .A(n950), .B(n951), .Z(n470) );
  ANDN U12784 ( .B(n952), .A(n953), .Z(n950) );
  AND U12785 ( .A(b[8]), .B(a[118]), .Z(n949) );
  XOR U12786 ( .A(n954), .B(n955), .Z(n463) );
  XOR U12787 ( .A(n956), .B(n957), .Z(n955) );
  AND U12788 ( .A(b[9]), .B(a[117]), .Z(n957) );
  AND U12789 ( .A(b[10]), .B(a[116]), .Z(n956) );
  XOR U12790 ( .A(n958), .B(n959), .Z(n954) );
  AND U12791 ( .A(b[11]), .B(a[115]), .Z(n959) );
  AND U12792 ( .A(b[12]), .B(a[114]), .Z(n958) );
  XOR U12793 ( .A(n960), .B(n961), .Z(n458) );
  XOR U12794 ( .A(n962), .B(n963), .Z(n961) );
  AND U12795 ( .A(b[3]), .B(a[123]), .Z(n963) );
  AND U12796 ( .A(b[4]), .B(a[122]), .Z(n962) );
  XOR U12797 ( .A(n964), .B(n965), .Z(n960) );
  AND U12798 ( .A(b[5]), .B(a[121]), .Z(n965) );
  AND U12799 ( .A(b[6]), .B(a[120]), .Z(n964) );
  XOR U12800 ( .A(n966), .B(n967), .Z(n456) );
  OR U12801 ( .A(n968), .B(n969), .Z(n967) );
  XOR U12802 ( .A(n970), .B(n971), .Z(n454) );
  XNOR U12803 ( .A(n972), .B(n462), .Z(n971) );
  NANDN U12804 ( .A(n973), .B(n974), .Z(n462) );
  AND U12805 ( .A(b[2]), .B(a[124]), .Z(n972) );
  AND U12806 ( .A(b[1]), .B(a[125]), .Z(n970) );
  NAND U12807 ( .A(a[126]), .B(b[0]), .Z(n446) );
  XNOR U12808 ( .A(n973), .B(n974), .Z(c[125]) );
  XOR U12809 ( .A(n968), .B(n969), .Z(n974) );
  XOR U12810 ( .A(n966), .B(n975), .Z(n969) );
  NAND U12811 ( .A(b[1]), .B(a[124]), .Z(n975) );
  XOR U12812 ( .A(n976), .B(n977), .Z(n968) );
  XOR U12813 ( .A(n966), .B(n978), .Z(n977) );
  XOR U12814 ( .A(n979), .B(n980), .Z(n978) );
  AND U12815 ( .A(b[2]), .B(a[123]), .Z(n979) );
  ANDN U12816 ( .B(n981), .A(n982), .Z(n966) );
  XOR U12817 ( .A(n983), .B(n984), .Z(n976) );
  XNOR U12818 ( .A(n980), .B(n985), .Z(n984) );
  XOR U12819 ( .A(n986), .B(n987), .Z(n985) );
  XOR U12820 ( .A(n988), .B(n989), .Z(n987) );
  XOR U12821 ( .A(n990), .B(n991), .Z(n989) );
  XOR U12822 ( .A(n992), .B(n993), .Z(n991) );
  XOR U12823 ( .A(n952), .B(n994), .Z(n993) );
  XNOR U12824 ( .A(n995), .B(n953), .Z(n994) );
  XOR U12825 ( .A(n996), .B(n997), .Z(n953) );
  XOR U12826 ( .A(n951), .B(n998), .Z(n997) );
  XOR U12827 ( .A(n999), .B(n1000), .Z(n998) );
  XOR U12828 ( .A(n1001), .B(n1002), .Z(n1000) );
  XOR U12829 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR U12830 ( .A(n1005), .B(n1006), .Z(n1004) );
  XOR U12831 ( .A(n1007), .B(n1008), .Z(n1006) );
  XOR U12832 ( .A(n1009), .B(n1010), .Z(n1008) );
  XOR U12833 ( .A(n1011), .B(n1012), .Z(n1010) );
  XOR U12834 ( .A(n1013), .B(n1014), .Z(n1012) );
  XOR U12835 ( .A(n941), .B(n1015), .Z(n1014) );
  XOR U12836 ( .A(n1016), .B(n942), .Z(n1015) );
  XOR U12837 ( .A(n1017), .B(n1018), .Z(n942) );
  XOR U12838 ( .A(n940), .B(n1019), .Z(n1018) );
  XOR U12839 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR U12840 ( .A(n1022), .B(n1023), .Z(n1021) );
  XOR U12841 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U12842 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR U12843 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U12844 ( .A(n1030), .B(n1031), .Z(n1029) );
  XOR U12845 ( .A(n938), .B(n1032), .Z(n1031) );
  XNOR U12846 ( .A(n1033), .B(n937), .Z(n1032) );
  XOR U12847 ( .A(n936), .B(n928), .Z(n1034) );
  XOR U12848 ( .A(n1035), .B(n1036), .Z(n928) );
  XOR U12849 ( .A(n926), .B(n1037), .Z(n1036) );
  XOR U12850 ( .A(n1038), .B(n1039), .Z(n1037) );
  XOR U12851 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U12852 ( .A(n1042), .B(n1043), .Z(n1041) );
  XOR U12853 ( .A(n1044), .B(n1045), .Z(n1043) );
  XOR U12854 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U12855 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U12856 ( .A(n924), .B(n1050), .Z(n1049) );
  XNOR U12857 ( .A(n1051), .B(n923), .Z(n1050) );
  XOR U12858 ( .A(n922), .B(n914), .Z(n1052) );
  XOR U12859 ( .A(n1053), .B(n1054), .Z(n914) );
  XOR U12860 ( .A(n912), .B(n1055), .Z(n1054) );
  XOR U12861 ( .A(n1056), .B(n1057), .Z(n1055) );
  XOR U12862 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U12863 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR U12864 ( .A(n1062), .B(n1063), .Z(n1061) );
  XOR U12865 ( .A(n1064), .B(n1065), .Z(n1063) );
  XOR U12866 ( .A(n1066), .B(n1067), .Z(n1065) );
  XOR U12867 ( .A(n910), .B(n1068), .Z(n1067) );
  XNOR U12868 ( .A(n1069), .B(n909), .Z(n1068) );
  XOR U12869 ( .A(n908), .B(n900), .Z(n1070) );
  XOR U12870 ( .A(n1071), .B(n1072), .Z(n900) );
  XOR U12871 ( .A(n898), .B(n1073), .Z(n1072) );
  XOR U12872 ( .A(n1074), .B(n1075), .Z(n1073) );
  XOR U12873 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U12874 ( .A(n1078), .B(n1079), .Z(n1077) );
  XOR U12875 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U12876 ( .A(n1082), .B(n1083), .Z(n1081) );
  XOR U12877 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U12878 ( .A(n896), .B(n1086), .Z(n1085) );
  XNOR U12879 ( .A(n1087), .B(n895), .Z(n1086) );
  XOR U12880 ( .A(n894), .B(n886), .Z(n1088) );
  XOR U12881 ( .A(n1089), .B(n1090), .Z(n886) );
  XOR U12882 ( .A(n884), .B(n1091), .Z(n1090) );
  XOR U12883 ( .A(n1092), .B(n1093), .Z(n1091) );
  XOR U12884 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U12885 ( .A(n1096), .B(n1097), .Z(n1095) );
  XOR U12886 ( .A(n1098), .B(n1099), .Z(n1097) );
  XOR U12887 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U12888 ( .A(n1102), .B(n1103), .Z(n1101) );
  XOR U12889 ( .A(n882), .B(n1104), .Z(n1103) );
  XNOR U12890 ( .A(n1105), .B(n881), .Z(n1104) );
  XOR U12891 ( .A(n880), .B(n872), .Z(n1106) );
  XOR U12892 ( .A(n1107), .B(n1108), .Z(n872) );
  XOR U12893 ( .A(n870), .B(n1109), .Z(n1108) );
  XOR U12894 ( .A(n1110), .B(n1111), .Z(n1109) );
  XOR U12895 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR U12896 ( .A(n1114), .B(n1115), .Z(n1113) );
  XOR U12897 ( .A(n1116), .B(n1117), .Z(n1115) );
  XOR U12898 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U12899 ( .A(n1120), .B(n1121), .Z(n1119) );
  XOR U12900 ( .A(n868), .B(n1122), .Z(n1121) );
  XNOR U12901 ( .A(n1123), .B(n867), .Z(n1122) );
  XOR U12902 ( .A(n866), .B(n858), .Z(n1124) );
  XOR U12903 ( .A(n1125), .B(n1126), .Z(n858) );
  XOR U12904 ( .A(n856), .B(n1127), .Z(n1126) );
  XOR U12905 ( .A(n1128), .B(n1129), .Z(n1127) );
  XOR U12906 ( .A(n1130), .B(n1131), .Z(n1129) );
  XOR U12907 ( .A(n1132), .B(n1133), .Z(n1131) );
  XOR U12908 ( .A(n1134), .B(n1135), .Z(n1133) );
  XOR U12909 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U12910 ( .A(n1138), .B(n1139), .Z(n1137) );
  XOR U12911 ( .A(n854), .B(n1140), .Z(n1139) );
  XNOR U12912 ( .A(n1141), .B(n853), .Z(n1140) );
  XOR U12913 ( .A(n852), .B(n844), .Z(n1142) );
  XOR U12914 ( .A(n1143), .B(n1144), .Z(n844) );
  XOR U12915 ( .A(n842), .B(n1145), .Z(n1144) );
  XOR U12916 ( .A(n1146), .B(n1147), .Z(n1145) );
  XOR U12917 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U12918 ( .A(n1150), .B(n1151), .Z(n1149) );
  XOR U12919 ( .A(n1152), .B(n1153), .Z(n1151) );
  XOR U12920 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U12921 ( .A(n1156), .B(n1157), .Z(n1155) );
  XOR U12922 ( .A(n840), .B(n1158), .Z(n1157) );
  XNOR U12923 ( .A(n1159), .B(n839), .Z(n1158) );
  XOR U12924 ( .A(n838), .B(n830), .Z(n1160) );
  XOR U12925 ( .A(n1161), .B(n1162), .Z(n830) );
  XOR U12926 ( .A(n828), .B(n1163), .Z(n1162) );
  XOR U12927 ( .A(n1164), .B(n1165), .Z(n1163) );
  XOR U12928 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U12929 ( .A(n1168), .B(n1169), .Z(n1167) );
  XOR U12930 ( .A(n1170), .B(n1171), .Z(n1169) );
  XOR U12931 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U12932 ( .A(n1174), .B(n1175), .Z(n1173) );
  XOR U12933 ( .A(n826), .B(n1176), .Z(n1175) );
  XNOR U12934 ( .A(n1177), .B(n825), .Z(n1176) );
  XOR U12935 ( .A(n824), .B(n816), .Z(n1178) );
  XOR U12936 ( .A(n1179), .B(n1180), .Z(n816) );
  XOR U12937 ( .A(n814), .B(n1181), .Z(n1180) );
  XOR U12938 ( .A(n1182), .B(n1183), .Z(n1181) );
  XOR U12939 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U12940 ( .A(n1186), .B(n1187), .Z(n1185) );
  XOR U12941 ( .A(n1188), .B(n1189), .Z(n1187) );
  XOR U12942 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U12943 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U12944 ( .A(n812), .B(n1194), .Z(n1193) );
  XNOR U12945 ( .A(n1195), .B(n811), .Z(n1194) );
  XOR U12946 ( .A(n810), .B(n802), .Z(n1196) );
  XOR U12947 ( .A(n1197), .B(n1198), .Z(n802) );
  XOR U12948 ( .A(n800), .B(n1199), .Z(n1198) );
  XOR U12949 ( .A(n1200), .B(n1201), .Z(n1199) );
  XOR U12950 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U12951 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U12952 ( .A(n1206), .B(n1207), .Z(n1205) );
  XOR U12953 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U12954 ( .A(n1210), .B(n1211), .Z(n1209) );
  XOR U12955 ( .A(n798), .B(n1212), .Z(n1211) );
  XNOR U12956 ( .A(n1213), .B(n797), .Z(n1212) );
  XOR U12957 ( .A(n796), .B(n788), .Z(n1214) );
  XOR U12958 ( .A(n1215), .B(n1216), .Z(n788) );
  XOR U12959 ( .A(n786), .B(n1217), .Z(n1216) );
  XOR U12960 ( .A(n1218), .B(n1219), .Z(n1217) );
  XOR U12961 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U12962 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U12963 ( .A(n1224), .B(n1225), .Z(n1223) );
  XOR U12964 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U12965 ( .A(n1228), .B(n1229), .Z(n1227) );
  XOR U12966 ( .A(n784), .B(n1230), .Z(n1229) );
  XNOR U12967 ( .A(n1231), .B(n783), .Z(n1230) );
  XOR U12968 ( .A(n782), .B(n774), .Z(n1232) );
  XOR U12969 ( .A(n1233), .B(n1234), .Z(n774) );
  XOR U12970 ( .A(n772), .B(n1235), .Z(n1234) );
  XOR U12971 ( .A(n1236), .B(n1237), .Z(n1235) );
  XOR U12972 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U12973 ( .A(n1240), .B(n1241), .Z(n1239) );
  XOR U12974 ( .A(n1242), .B(n1243), .Z(n1241) );
  XOR U12975 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U12976 ( .A(n1246), .B(n1247), .Z(n1245) );
  XOR U12977 ( .A(n770), .B(n1248), .Z(n1247) );
  XNOR U12978 ( .A(n1249), .B(n769), .Z(n1248) );
  XOR U12979 ( .A(n768), .B(n760), .Z(n1250) );
  XOR U12980 ( .A(n1251), .B(n1252), .Z(n760) );
  XOR U12981 ( .A(n758), .B(n1253), .Z(n1252) );
  XOR U12982 ( .A(n1254), .B(n1255), .Z(n1253) );
  XOR U12983 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U12984 ( .A(n1258), .B(n1259), .Z(n1257) );
  XOR U12985 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR U12986 ( .A(n1262), .B(n1263), .Z(n1261) );
  XOR U12987 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U12988 ( .A(n756), .B(n1266), .Z(n1265) );
  XNOR U12989 ( .A(n1267), .B(n755), .Z(n1266) );
  XOR U12990 ( .A(n754), .B(n746), .Z(n1268) );
  XOR U12991 ( .A(n1269), .B(n1270), .Z(n746) );
  XOR U12992 ( .A(n744), .B(n1271), .Z(n1270) );
  XOR U12993 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U12994 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U12995 ( .A(n1276), .B(n1277), .Z(n1275) );
  XOR U12996 ( .A(n1278), .B(n1279), .Z(n1277) );
  XOR U12997 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U12998 ( .A(n1282), .B(n1283), .Z(n1281) );
  XOR U12999 ( .A(n742), .B(n1284), .Z(n1283) );
  XNOR U13000 ( .A(n1285), .B(n741), .Z(n1284) );
  XOR U13001 ( .A(n740), .B(n732), .Z(n1286) );
  XOR U13002 ( .A(n1287), .B(n1288), .Z(n732) );
  XOR U13003 ( .A(n730), .B(n1289), .Z(n1288) );
  XOR U13004 ( .A(n1290), .B(n1291), .Z(n1289) );
  XOR U13005 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U13006 ( .A(n1294), .B(n1295), .Z(n1293) );
  XOR U13007 ( .A(n1296), .B(n1297), .Z(n1295) );
  XOR U13008 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U13009 ( .A(n1300), .B(n1301), .Z(n1299) );
  XOR U13010 ( .A(n728), .B(n1302), .Z(n1301) );
  XNOR U13011 ( .A(n1303), .B(n727), .Z(n1302) );
  XOR U13012 ( .A(n726), .B(n718), .Z(n1304) );
  XOR U13013 ( .A(n1305), .B(n1306), .Z(n718) );
  XOR U13014 ( .A(n716), .B(n1307), .Z(n1306) );
  XOR U13015 ( .A(n1308), .B(n1309), .Z(n1307) );
  XOR U13016 ( .A(n1310), .B(n1311), .Z(n1309) );
  XOR U13017 ( .A(n1312), .B(n1313), .Z(n1311) );
  XOR U13018 ( .A(n1314), .B(n1315), .Z(n1313) );
  XOR U13019 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U13020 ( .A(n1318), .B(n1319), .Z(n1317) );
  XOR U13021 ( .A(n714), .B(n1320), .Z(n1319) );
  XNOR U13022 ( .A(n1321), .B(n713), .Z(n1320) );
  XOR U13023 ( .A(n712), .B(n704), .Z(n1322) );
  XOR U13024 ( .A(n1323), .B(n1324), .Z(n704) );
  XOR U13025 ( .A(n702), .B(n1325), .Z(n1324) );
  XOR U13026 ( .A(n1326), .B(n1327), .Z(n1325) );
  XOR U13027 ( .A(n1328), .B(n1329), .Z(n1327) );
  XOR U13028 ( .A(n1330), .B(n1331), .Z(n1329) );
  XOR U13029 ( .A(n1332), .B(n1333), .Z(n1331) );
  XOR U13030 ( .A(n1334), .B(n1335), .Z(n1333) );
  XOR U13031 ( .A(n1336), .B(n1337), .Z(n1335) );
  XOR U13032 ( .A(n693), .B(n1338), .Z(n1337) );
  XOR U13033 ( .A(n1339), .B(n694), .Z(n1338) );
  XOR U13034 ( .A(n1340), .B(n1341), .Z(n694) );
  XOR U13035 ( .A(n692), .B(n1342), .Z(n1341) );
  XOR U13036 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U13037 ( .A(n1345), .B(n1346), .Z(n1344) );
  XOR U13038 ( .A(n1347), .B(n1348), .Z(n1346) );
  XOR U13039 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U13040 ( .A(n1351), .B(n1352), .Z(n1350) );
  XOR U13041 ( .A(n1353), .B(n1354), .Z(n1352) );
  XOR U13042 ( .A(n1355), .B(n1356), .Z(n1354) );
  XOR U13043 ( .A(n1357), .B(n1358), .Z(n1356) );
  XOR U13044 ( .A(n1359), .B(n1360), .Z(n1358) );
  AND U13045 ( .A(a[0]), .B(b[125]), .Z(n1359) );
  XNOR U13046 ( .A(n1361), .B(n1360), .Z(n1355) );
  XNOR U13047 ( .A(n1362), .B(n1363), .Z(n1360) );
  ANDN U13048 ( .B(n1364), .A(n1365), .Z(n1362) );
  AND U13049 ( .A(a[1]), .B(b[124]), .Z(n1361) );
  XOR U13050 ( .A(n1366), .B(n1357), .Z(n1351) );
  XOR U13051 ( .A(n1367), .B(n1368), .Z(n1357) );
  ANDN U13052 ( .B(n1369), .A(n1370), .Z(n1367) );
  AND U13053 ( .A(a[2]), .B(b[123]), .Z(n1366) );
  XOR U13054 ( .A(n1371), .B(n1353), .Z(n1347) );
  XOR U13055 ( .A(n1372), .B(n1373), .Z(n1353) );
  ANDN U13056 ( .B(n1374), .A(n1375), .Z(n1372) );
  AND U13057 ( .A(a[3]), .B(b[122]), .Z(n1371) );
  XOR U13058 ( .A(n1376), .B(n1349), .Z(n1343) );
  XOR U13059 ( .A(n1377), .B(n1378), .Z(n1349) );
  ANDN U13060 ( .B(n1379), .A(n1380), .Z(n1377) );
  AND U13061 ( .A(a[4]), .B(b[121]), .Z(n1376) );
  XOR U13062 ( .A(n1381), .B(n1345), .Z(n1340) );
  XOR U13063 ( .A(n1382), .B(n1383), .Z(n1345) );
  ANDN U13064 ( .B(n1384), .A(n1385), .Z(n1382) );
  AND U13065 ( .A(a[5]), .B(b[120]), .Z(n1381) );
  XOR U13066 ( .A(n1386), .B(n692), .Z(n693) );
  XOR U13067 ( .A(n1387), .B(n1388), .Z(n692) );
  ANDN U13068 ( .B(n1389), .A(n1390), .Z(n1387) );
  AND U13069 ( .A(a[6]), .B(b[119]), .Z(n1386) );
  XOR U13070 ( .A(n1391), .B(n1339), .Z(n1334) );
  XOR U13071 ( .A(n1392), .B(n1393), .Z(n1339) );
  ANDN U13072 ( .B(n1394), .A(n1395), .Z(n1392) );
  AND U13073 ( .A(a[7]), .B(b[118]), .Z(n1391) );
  XOR U13074 ( .A(n1396), .B(n1336), .Z(n1330) );
  XOR U13075 ( .A(n1397), .B(n1398), .Z(n1336) );
  ANDN U13076 ( .B(n1399), .A(n1400), .Z(n1397) );
  AND U13077 ( .A(a[8]), .B(b[117]), .Z(n1396) );
  XOR U13078 ( .A(n1401), .B(n1332), .Z(n1326) );
  XOR U13079 ( .A(n1402), .B(n1403), .Z(n1332) );
  ANDN U13080 ( .B(n1404), .A(n1405), .Z(n1402) );
  AND U13081 ( .A(a[9]), .B(b[116]), .Z(n1401) );
  XOR U13082 ( .A(n1406), .B(n1328), .Z(n1323) );
  XOR U13083 ( .A(n1407), .B(n1408), .Z(n1328) );
  ANDN U13084 ( .B(n1409), .A(n1410), .Z(n1407) );
  AND U13085 ( .A(a[10]), .B(b[115]), .Z(n1406) );
  XNOR U13086 ( .A(n1411), .B(n702), .Z(n703) );
  XOR U13087 ( .A(n1412), .B(n1413), .Z(n702) );
  ANDN U13088 ( .B(n1414), .A(n1415), .Z(n1412) );
  AND U13089 ( .A(a[11]), .B(b[114]), .Z(n1411) );
  XOR U13090 ( .A(n1416), .B(n712), .Z(n714) );
  XOR U13091 ( .A(n1417), .B(n1418), .Z(n712) );
  ANDN U13092 ( .B(n1419), .A(n1420), .Z(n1417) );
  AND U13093 ( .A(a[12]), .B(b[113]), .Z(n1416) );
  XOR U13094 ( .A(n1421), .B(n1321), .Z(n1316) );
  XOR U13095 ( .A(n1422), .B(n1423), .Z(n1321) );
  ANDN U13096 ( .B(n1424), .A(n1425), .Z(n1422) );
  AND U13097 ( .A(a[13]), .B(b[112]), .Z(n1421) );
  XOR U13098 ( .A(n1426), .B(n1318), .Z(n1312) );
  XOR U13099 ( .A(n1427), .B(n1428), .Z(n1318) );
  ANDN U13100 ( .B(n1429), .A(n1430), .Z(n1427) );
  AND U13101 ( .A(a[14]), .B(b[111]), .Z(n1426) );
  XOR U13102 ( .A(n1431), .B(n1314), .Z(n1308) );
  XOR U13103 ( .A(n1432), .B(n1433), .Z(n1314) );
  ANDN U13104 ( .B(n1434), .A(n1435), .Z(n1432) );
  AND U13105 ( .A(a[15]), .B(b[110]), .Z(n1431) );
  XOR U13106 ( .A(n1436), .B(n1310), .Z(n1305) );
  XOR U13107 ( .A(n1437), .B(n1438), .Z(n1310) );
  ANDN U13108 ( .B(n1439), .A(n1440), .Z(n1437) );
  AND U13109 ( .A(a[16]), .B(b[109]), .Z(n1436) );
  XNOR U13110 ( .A(n1441), .B(n716), .Z(n717) );
  XOR U13111 ( .A(n1442), .B(n1443), .Z(n716) );
  ANDN U13112 ( .B(n1444), .A(n1445), .Z(n1442) );
  AND U13113 ( .A(a[17]), .B(b[108]), .Z(n1441) );
  XOR U13114 ( .A(n1446), .B(n726), .Z(n728) );
  XOR U13115 ( .A(n1447), .B(n1448), .Z(n726) );
  ANDN U13116 ( .B(n1449), .A(n1450), .Z(n1447) );
  AND U13117 ( .A(a[18]), .B(b[107]), .Z(n1446) );
  XOR U13118 ( .A(n1451), .B(n1303), .Z(n1298) );
  XOR U13119 ( .A(n1452), .B(n1453), .Z(n1303) );
  ANDN U13120 ( .B(n1454), .A(n1455), .Z(n1452) );
  AND U13121 ( .A(a[19]), .B(b[106]), .Z(n1451) );
  XOR U13122 ( .A(n1456), .B(n1300), .Z(n1294) );
  XOR U13123 ( .A(n1457), .B(n1458), .Z(n1300) );
  ANDN U13124 ( .B(n1459), .A(n1460), .Z(n1457) );
  AND U13125 ( .A(a[20]), .B(b[105]), .Z(n1456) );
  XOR U13126 ( .A(n1461), .B(n1296), .Z(n1290) );
  XOR U13127 ( .A(n1462), .B(n1463), .Z(n1296) );
  ANDN U13128 ( .B(n1464), .A(n1465), .Z(n1462) );
  AND U13129 ( .A(a[21]), .B(b[104]), .Z(n1461) );
  XOR U13130 ( .A(n1466), .B(n1292), .Z(n1287) );
  XOR U13131 ( .A(n1467), .B(n1468), .Z(n1292) );
  ANDN U13132 ( .B(n1469), .A(n1470), .Z(n1467) );
  AND U13133 ( .A(a[22]), .B(b[103]), .Z(n1466) );
  XNOR U13134 ( .A(n1471), .B(n730), .Z(n731) );
  XOR U13135 ( .A(n1472), .B(n1473), .Z(n730) );
  ANDN U13136 ( .B(n1474), .A(n1475), .Z(n1472) );
  AND U13137 ( .A(a[23]), .B(b[102]), .Z(n1471) );
  XOR U13138 ( .A(n1476), .B(n740), .Z(n742) );
  XOR U13139 ( .A(n1477), .B(n1478), .Z(n740) );
  ANDN U13140 ( .B(n1479), .A(n1480), .Z(n1477) );
  AND U13141 ( .A(a[24]), .B(b[101]), .Z(n1476) );
  XOR U13142 ( .A(n1481), .B(n1285), .Z(n1280) );
  XOR U13143 ( .A(n1482), .B(n1483), .Z(n1285) );
  ANDN U13144 ( .B(n1484), .A(n1485), .Z(n1482) );
  AND U13145 ( .A(a[25]), .B(b[100]), .Z(n1481) );
  XOR U13146 ( .A(n1486), .B(n1282), .Z(n1276) );
  XOR U13147 ( .A(n1487), .B(n1488), .Z(n1282) );
  ANDN U13148 ( .B(n1489), .A(n1490), .Z(n1487) );
  AND U13149 ( .A(a[26]), .B(b[99]), .Z(n1486) );
  XOR U13150 ( .A(n1491), .B(n1278), .Z(n1272) );
  XOR U13151 ( .A(n1492), .B(n1493), .Z(n1278) );
  ANDN U13152 ( .B(n1494), .A(n1495), .Z(n1492) );
  AND U13153 ( .A(a[27]), .B(b[98]), .Z(n1491) );
  XOR U13154 ( .A(n1496), .B(n1274), .Z(n1269) );
  XOR U13155 ( .A(n1497), .B(n1498), .Z(n1274) );
  ANDN U13156 ( .B(n1499), .A(n1500), .Z(n1497) );
  AND U13157 ( .A(a[28]), .B(b[97]), .Z(n1496) );
  XNOR U13158 ( .A(n1501), .B(n744), .Z(n745) );
  XOR U13159 ( .A(n1502), .B(n1503), .Z(n744) );
  ANDN U13160 ( .B(n1504), .A(n1505), .Z(n1502) );
  AND U13161 ( .A(a[29]), .B(b[96]), .Z(n1501) );
  XOR U13162 ( .A(n1506), .B(n754), .Z(n756) );
  XOR U13163 ( .A(n1507), .B(n1508), .Z(n754) );
  ANDN U13164 ( .B(n1509), .A(n1510), .Z(n1507) );
  AND U13165 ( .A(a[30]), .B(b[95]), .Z(n1506) );
  XOR U13166 ( .A(n1511), .B(n1267), .Z(n1262) );
  XOR U13167 ( .A(n1512), .B(n1513), .Z(n1267) );
  ANDN U13168 ( .B(n1514), .A(n1515), .Z(n1512) );
  AND U13169 ( .A(a[31]), .B(b[94]), .Z(n1511) );
  XOR U13170 ( .A(n1516), .B(n1264), .Z(n1258) );
  XOR U13171 ( .A(n1517), .B(n1518), .Z(n1264) );
  ANDN U13172 ( .B(n1519), .A(n1520), .Z(n1517) );
  AND U13173 ( .A(a[32]), .B(b[93]), .Z(n1516) );
  XOR U13174 ( .A(n1521), .B(n1260), .Z(n1254) );
  XOR U13175 ( .A(n1522), .B(n1523), .Z(n1260) );
  ANDN U13176 ( .B(n1524), .A(n1525), .Z(n1522) );
  AND U13177 ( .A(a[33]), .B(b[92]), .Z(n1521) );
  XOR U13178 ( .A(n1526), .B(n1256), .Z(n1251) );
  XOR U13179 ( .A(n1527), .B(n1528), .Z(n1256) );
  ANDN U13180 ( .B(n1529), .A(n1530), .Z(n1527) );
  AND U13181 ( .A(a[34]), .B(b[91]), .Z(n1526) );
  XNOR U13182 ( .A(n1531), .B(n758), .Z(n759) );
  XOR U13183 ( .A(n1532), .B(n1533), .Z(n758) );
  ANDN U13184 ( .B(n1534), .A(n1535), .Z(n1532) );
  AND U13185 ( .A(a[35]), .B(b[90]), .Z(n1531) );
  XOR U13186 ( .A(n1536), .B(n768), .Z(n770) );
  XOR U13187 ( .A(n1537), .B(n1538), .Z(n768) );
  ANDN U13188 ( .B(n1539), .A(n1540), .Z(n1537) );
  AND U13189 ( .A(a[36]), .B(b[89]), .Z(n1536) );
  XOR U13190 ( .A(n1541), .B(n1249), .Z(n1244) );
  XOR U13191 ( .A(n1542), .B(n1543), .Z(n1249) );
  ANDN U13192 ( .B(n1544), .A(n1545), .Z(n1542) );
  AND U13193 ( .A(a[37]), .B(b[88]), .Z(n1541) );
  XOR U13194 ( .A(n1546), .B(n1246), .Z(n1240) );
  XOR U13195 ( .A(n1547), .B(n1548), .Z(n1246) );
  ANDN U13196 ( .B(n1549), .A(n1550), .Z(n1547) );
  AND U13197 ( .A(a[38]), .B(b[87]), .Z(n1546) );
  XOR U13198 ( .A(n1551), .B(n1242), .Z(n1236) );
  XOR U13199 ( .A(n1552), .B(n1553), .Z(n1242) );
  ANDN U13200 ( .B(n1554), .A(n1555), .Z(n1552) );
  AND U13201 ( .A(a[39]), .B(b[86]), .Z(n1551) );
  XOR U13202 ( .A(n1556), .B(n1238), .Z(n1233) );
  XOR U13203 ( .A(n1557), .B(n1558), .Z(n1238) );
  ANDN U13204 ( .B(n1559), .A(n1560), .Z(n1557) );
  AND U13205 ( .A(a[40]), .B(b[85]), .Z(n1556) );
  XNOR U13206 ( .A(n1561), .B(n772), .Z(n773) );
  XOR U13207 ( .A(n1562), .B(n1563), .Z(n772) );
  ANDN U13208 ( .B(n1564), .A(n1565), .Z(n1562) );
  AND U13209 ( .A(a[41]), .B(b[84]), .Z(n1561) );
  XOR U13210 ( .A(n1566), .B(n782), .Z(n784) );
  XOR U13211 ( .A(n1567), .B(n1568), .Z(n782) );
  ANDN U13212 ( .B(n1569), .A(n1570), .Z(n1567) );
  AND U13213 ( .A(a[42]), .B(b[83]), .Z(n1566) );
  XOR U13214 ( .A(n1571), .B(n1231), .Z(n1226) );
  XOR U13215 ( .A(n1572), .B(n1573), .Z(n1231) );
  ANDN U13216 ( .B(n1574), .A(n1575), .Z(n1572) );
  AND U13217 ( .A(a[43]), .B(b[82]), .Z(n1571) );
  XOR U13218 ( .A(n1576), .B(n1228), .Z(n1222) );
  XOR U13219 ( .A(n1577), .B(n1578), .Z(n1228) );
  ANDN U13220 ( .B(n1579), .A(n1580), .Z(n1577) );
  AND U13221 ( .A(a[44]), .B(b[81]), .Z(n1576) );
  XOR U13222 ( .A(n1581), .B(n1224), .Z(n1218) );
  XOR U13223 ( .A(n1582), .B(n1583), .Z(n1224) );
  ANDN U13224 ( .B(n1584), .A(n1585), .Z(n1582) );
  AND U13225 ( .A(a[45]), .B(b[80]), .Z(n1581) );
  XOR U13226 ( .A(n1586), .B(n1220), .Z(n1215) );
  XOR U13227 ( .A(n1587), .B(n1588), .Z(n1220) );
  ANDN U13228 ( .B(n1589), .A(n1590), .Z(n1587) );
  AND U13229 ( .A(a[46]), .B(b[79]), .Z(n1586) );
  XNOR U13230 ( .A(n1591), .B(n786), .Z(n787) );
  XOR U13231 ( .A(n1592), .B(n1593), .Z(n786) );
  ANDN U13232 ( .B(n1594), .A(n1595), .Z(n1592) );
  AND U13233 ( .A(a[47]), .B(b[78]), .Z(n1591) );
  XOR U13234 ( .A(n1596), .B(n796), .Z(n798) );
  XOR U13235 ( .A(n1597), .B(n1598), .Z(n796) );
  ANDN U13236 ( .B(n1599), .A(n1600), .Z(n1597) );
  AND U13237 ( .A(a[48]), .B(b[77]), .Z(n1596) );
  XOR U13238 ( .A(n1601), .B(n1213), .Z(n1208) );
  XOR U13239 ( .A(n1602), .B(n1603), .Z(n1213) );
  ANDN U13240 ( .B(n1604), .A(n1605), .Z(n1602) );
  AND U13241 ( .A(a[49]), .B(b[76]), .Z(n1601) );
  XOR U13242 ( .A(n1606), .B(n1210), .Z(n1204) );
  XOR U13243 ( .A(n1607), .B(n1608), .Z(n1210) );
  ANDN U13244 ( .B(n1609), .A(n1610), .Z(n1607) );
  AND U13245 ( .A(a[50]), .B(b[75]), .Z(n1606) );
  XOR U13246 ( .A(n1611), .B(n1206), .Z(n1200) );
  XOR U13247 ( .A(n1612), .B(n1613), .Z(n1206) );
  ANDN U13248 ( .B(n1614), .A(n1615), .Z(n1612) );
  AND U13249 ( .A(a[51]), .B(b[74]), .Z(n1611) );
  XOR U13250 ( .A(n1616), .B(n1202), .Z(n1197) );
  XOR U13251 ( .A(n1617), .B(n1618), .Z(n1202) );
  ANDN U13252 ( .B(n1619), .A(n1620), .Z(n1617) );
  AND U13253 ( .A(a[52]), .B(b[73]), .Z(n1616) );
  XNOR U13254 ( .A(n1621), .B(n800), .Z(n801) );
  XOR U13255 ( .A(n1622), .B(n1623), .Z(n800) );
  ANDN U13256 ( .B(n1624), .A(n1625), .Z(n1622) );
  AND U13257 ( .A(a[53]), .B(b[72]), .Z(n1621) );
  XOR U13258 ( .A(n1626), .B(n810), .Z(n812) );
  XOR U13259 ( .A(n1627), .B(n1628), .Z(n810) );
  ANDN U13260 ( .B(n1629), .A(n1630), .Z(n1627) );
  AND U13261 ( .A(a[54]), .B(b[71]), .Z(n1626) );
  XOR U13262 ( .A(n1631), .B(n1195), .Z(n1190) );
  XOR U13263 ( .A(n1632), .B(n1633), .Z(n1195) );
  ANDN U13264 ( .B(n1634), .A(n1635), .Z(n1632) );
  AND U13265 ( .A(a[55]), .B(b[70]), .Z(n1631) );
  XOR U13266 ( .A(n1636), .B(n1192), .Z(n1186) );
  XOR U13267 ( .A(n1637), .B(n1638), .Z(n1192) );
  ANDN U13268 ( .B(n1639), .A(n1640), .Z(n1637) );
  AND U13269 ( .A(a[56]), .B(b[69]), .Z(n1636) );
  XOR U13270 ( .A(n1641), .B(n1188), .Z(n1182) );
  XOR U13271 ( .A(n1642), .B(n1643), .Z(n1188) );
  ANDN U13272 ( .B(n1644), .A(n1645), .Z(n1642) );
  AND U13273 ( .A(a[57]), .B(b[68]), .Z(n1641) );
  XOR U13274 ( .A(n1646), .B(n1184), .Z(n1179) );
  XOR U13275 ( .A(n1647), .B(n1648), .Z(n1184) );
  ANDN U13276 ( .B(n1649), .A(n1650), .Z(n1647) );
  AND U13277 ( .A(a[58]), .B(b[67]), .Z(n1646) );
  XNOR U13278 ( .A(n1651), .B(n814), .Z(n815) );
  XOR U13279 ( .A(n1652), .B(n1653), .Z(n814) );
  ANDN U13280 ( .B(n1654), .A(n1655), .Z(n1652) );
  AND U13281 ( .A(a[59]), .B(b[66]), .Z(n1651) );
  XOR U13282 ( .A(n1656), .B(n824), .Z(n826) );
  XOR U13283 ( .A(n1657), .B(n1658), .Z(n824) );
  ANDN U13284 ( .B(n1659), .A(n1660), .Z(n1657) );
  AND U13285 ( .A(a[60]), .B(b[65]), .Z(n1656) );
  XOR U13286 ( .A(n1661), .B(n1177), .Z(n1172) );
  XOR U13287 ( .A(n1662), .B(n1663), .Z(n1177) );
  ANDN U13288 ( .B(n1664), .A(n1665), .Z(n1662) );
  AND U13289 ( .A(a[61]), .B(b[64]), .Z(n1661) );
  XOR U13290 ( .A(n1666), .B(n1174), .Z(n1168) );
  XOR U13291 ( .A(n1667), .B(n1668), .Z(n1174) );
  ANDN U13292 ( .B(n1669), .A(n1670), .Z(n1667) );
  AND U13293 ( .A(a[62]), .B(b[63]), .Z(n1666) );
  XOR U13294 ( .A(n1671), .B(n1170), .Z(n1164) );
  XOR U13295 ( .A(n1672), .B(n1673), .Z(n1170) );
  ANDN U13296 ( .B(n1674), .A(n1675), .Z(n1672) );
  AND U13297 ( .A(a[63]), .B(b[62]), .Z(n1671) );
  XOR U13298 ( .A(n1676), .B(n1166), .Z(n1161) );
  XOR U13299 ( .A(n1677), .B(n1678), .Z(n1166) );
  ANDN U13300 ( .B(n1679), .A(n1680), .Z(n1677) );
  AND U13301 ( .A(a[64]), .B(b[61]), .Z(n1676) );
  XNOR U13302 ( .A(n1681), .B(n828), .Z(n829) );
  XOR U13303 ( .A(n1682), .B(n1683), .Z(n828) );
  ANDN U13304 ( .B(n1684), .A(n1685), .Z(n1682) );
  AND U13305 ( .A(a[65]), .B(b[60]), .Z(n1681) );
  XOR U13306 ( .A(n1686), .B(n838), .Z(n840) );
  XOR U13307 ( .A(n1687), .B(n1688), .Z(n838) );
  ANDN U13308 ( .B(n1689), .A(n1690), .Z(n1687) );
  AND U13309 ( .A(a[66]), .B(b[59]), .Z(n1686) );
  XOR U13310 ( .A(n1691), .B(n1159), .Z(n1154) );
  XOR U13311 ( .A(n1692), .B(n1693), .Z(n1159) );
  ANDN U13312 ( .B(n1694), .A(n1695), .Z(n1692) );
  AND U13313 ( .A(a[67]), .B(b[58]), .Z(n1691) );
  XOR U13314 ( .A(n1696), .B(n1156), .Z(n1150) );
  XOR U13315 ( .A(n1697), .B(n1698), .Z(n1156) );
  ANDN U13316 ( .B(n1699), .A(n1700), .Z(n1697) );
  AND U13317 ( .A(a[68]), .B(b[57]), .Z(n1696) );
  XOR U13318 ( .A(n1701), .B(n1152), .Z(n1146) );
  XOR U13319 ( .A(n1702), .B(n1703), .Z(n1152) );
  ANDN U13320 ( .B(n1704), .A(n1705), .Z(n1702) );
  AND U13321 ( .A(a[69]), .B(b[56]), .Z(n1701) );
  XOR U13322 ( .A(n1706), .B(n1148), .Z(n1143) );
  XOR U13323 ( .A(n1707), .B(n1708), .Z(n1148) );
  ANDN U13324 ( .B(n1709), .A(n1710), .Z(n1707) );
  AND U13325 ( .A(a[70]), .B(b[55]), .Z(n1706) );
  XNOR U13326 ( .A(n1711), .B(n842), .Z(n843) );
  XOR U13327 ( .A(n1712), .B(n1713), .Z(n842) );
  ANDN U13328 ( .B(n1714), .A(n1715), .Z(n1712) );
  AND U13329 ( .A(a[71]), .B(b[54]), .Z(n1711) );
  XOR U13330 ( .A(n1716), .B(n852), .Z(n854) );
  XOR U13331 ( .A(n1717), .B(n1718), .Z(n852) );
  ANDN U13332 ( .B(n1719), .A(n1720), .Z(n1717) );
  AND U13333 ( .A(a[72]), .B(b[53]), .Z(n1716) );
  XOR U13334 ( .A(n1721), .B(n1141), .Z(n1136) );
  XOR U13335 ( .A(n1722), .B(n1723), .Z(n1141) );
  ANDN U13336 ( .B(n1724), .A(n1725), .Z(n1722) );
  AND U13337 ( .A(a[73]), .B(b[52]), .Z(n1721) );
  XOR U13338 ( .A(n1726), .B(n1138), .Z(n1132) );
  XOR U13339 ( .A(n1727), .B(n1728), .Z(n1138) );
  ANDN U13340 ( .B(n1729), .A(n1730), .Z(n1727) );
  AND U13341 ( .A(a[74]), .B(b[51]), .Z(n1726) );
  XOR U13342 ( .A(n1731), .B(n1134), .Z(n1128) );
  XOR U13343 ( .A(n1732), .B(n1733), .Z(n1134) );
  ANDN U13344 ( .B(n1734), .A(n1735), .Z(n1732) );
  AND U13345 ( .A(a[75]), .B(b[50]), .Z(n1731) );
  XOR U13346 ( .A(n1736), .B(n1130), .Z(n1125) );
  XOR U13347 ( .A(n1737), .B(n1738), .Z(n1130) );
  ANDN U13348 ( .B(n1739), .A(n1740), .Z(n1737) );
  AND U13349 ( .A(a[76]), .B(b[49]), .Z(n1736) );
  XNOR U13350 ( .A(n1741), .B(n856), .Z(n857) );
  XOR U13351 ( .A(n1742), .B(n1743), .Z(n856) );
  ANDN U13352 ( .B(n1744), .A(n1745), .Z(n1742) );
  AND U13353 ( .A(a[77]), .B(b[48]), .Z(n1741) );
  XOR U13354 ( .A(n1746), .B(n866), .Z(n868) );
  XOR U13355 ( .A(n1747), .B(n1748), .Z(n866) );
  ANDN U13356 ( .B(n1749), .A(n1750), .Z(n1747) );
  AND U13357 ( .A(a[78]), .B(b[47]), .Z(n1746) );
  XOR U13358 ( .A(n1751), .B(n1123), .Z(n1118) );
  XOR U13359 ( .A(n1752), .B(n1753), .Z(n1123) );
  ANDN U13360 ( .B(n1754), .A(n1755), .Z(n1752) );
  AND U13361 ( .A(a[79]), .B(b[46]), .Z(n1751) );
  XOR U13362 ( .A(n1756), .B(n1120), .Z(n1114) );
  XOR U13363 ( .A(n1757), .B(n1758), .Z(n1120) );
  ANDN U13364 ( .B(n1759), .A(n1760), .Z(n1757) );
  AND U13365 ( .A(a[80]), .B(b[45]), .Z(n1756) );
  XOR U13366 ( .A(n1761), .B(n1116), .Z(n1110) );
  XOR U13367 ( .A(n1762), .B(n1763), .Z(n1116) );
  ANDN U13368 ( .B(n1764), .A(n1765), .Z(n1762) );
  AND U13369 ( .A(a[81]), .B(b[44]), .Z(n1761) );
  XOR U13370 ( .A(n1766), .B(n1112), .Z(n1107) );
  XOR U13371 ( .A(n1767), .B(n1768), .Z(n1112) );
  ANDN U13372 ( .B(n1769), .A(n1770), .Z(n1767) );
  AND U13373 ( .A(a[82]), .B(b[43]), .Z(n1766) );
  XNOR U13374 ( .A(n1771), .B(n870), .Z(n871) );
  XOR U13375 ( .A(n1772), .B(n1773), .Z(n870) );
  ANDN U13376 ( .B(n1774), .A(n1775), .Z(n1772) );
  AND U13377 ( .A(a[83]), .B(b[42]), .Z(n1771) );
  XOR U13378 ( .A(n1776), .B(n880), .Z(n882) );
  XOR U13379 ( .A(n1777), .B(n1778), .Z(n880) );
  ANDN U13380 ( .B(n1779), .A(n1780), .Z(n1777) );
  AND U13381 ( .A(a[84]), .B(b[41]), .Z(n1776) );
  XOR U13382 ( .A(n1781), .B(n1105), .Z(n1100) );
  XOR U13383 ( .A(n1782), .B(n1783), .Z(n1105) );
  ANDN U13384 ( .B(n1784), .A(n1785), .Z(n1782) );
  AND U13385 ( .A(a[85]), .B(b[40]), .Z(n1781) );
  XOR U13386 ( .A(n1786), .B(n1102), .Z(n1096) );
  XOR U13387 ( .A(n1787), .B(n1788), .Z(n1102) );
  ANDN U13388 ( .B(n1789), .A(n1790), .Z(n1787) );
  AND U13389 ( .A(a[86]), .B(b[39]), .Z(n1786) );
  XOR U13390 ( .A(n1791), .B(n1098), .Z(n1092) );
  XOR U13391 ( .A(n1792), .B(n1793), .Z(n1098) );
  ANDN U13392 ( .B(n1794), .A(n1795), .Z(n1792) );
  AND U13393 ( .A(a[87]), .B(b[38]), .Z(n1791) );
  XOR U13394 ( .A(n1796), .B(n1094), .Z(n1089) );
  XOR U13395 ( .A(n1797), .B(n1798), .Z(n1094) );
  ANDN U13396 ( .B(n1799), .A(n1800), .Z(n1797) );
  AND U13397 ( .A(a[88]), .B(b[37]), .Z(n1796) );
  XNOR U13398 ( .A(n1801), .B(n884), .Z(n885) );
  XOR U13399 ( .A(n1802), .B(n1803), .Z(n884) );
  ANDN U13400 ( .B(n1804), .A(n1805), .Z(n1802) );
  AND U13401 ( .A(a[89]), .B(b[36]), .Z(n1801) );
  XOR U13402 ( .A(n1806), .B(n894), .Z(n896) );
  XOR U13403 ( .A(n1807), .B(n1808), .Z(n894) );
  ANDN U13404 ( .B(n1809), .A(n1810), .Z(n1807) );
  AND U13405 ( .A(a[90]), .B(b[35]), .Z(n1806) );
  XOR U13406 ( .A(n1811), .B(n1087), .Z(n1082) );
  XOR U13407 ( .A(n1812), .B(n1813), .Z(n1087) );
  ANDN U13408 ( .B(n1814), .A(n1815), .Z(n1812) );
  AND U13409 ( .A(a[91]), .B(b[34]), .Z(n1811) );
  XOR U13410 ( .A(n1816), .B(n1084), .Z(n1078) );
  XOR U13411 ( .A(n1817), .B(n1818), .Z(n1084) );
  ANDN U13412 ( .B(n1819), .A(n1820), .Z(n1817) );
  AND U13413 ( .A(a[92]), .B(b[33]), .Z(n1816) );
  XOR U13414 ( .A(n1821), .B(n1080), .Z(n1074) );
  XOR U13415 ( .A(n1822), .B(n1823), .Z(n1080) );
  ANDN U13416 ( .B(n1824), .A(n1825), .Z(n1822) );
  AND U13417 ( .A(a[93]), .B(b[32]), .Z(n1821) );
  XOR U13418 ( .A(n1826), .B(n1076), .Z(n1071) );
  XOR U13419 ( .A(n1827), .B(n1828), .Z(n1076) );
  ANDN U13420 ( .B(n1829), .A(n1830), .Z(n1827) );
  AND U13421 ( .A(a[94]), .B(b[31]), .Z(n1826) );
  XNOR U13422 ( .A(n1831), .B(n898), .Z(n899) );
  XOR U13423 ( .A(n1832), .B(n1833), .Z(n898) );
  ANDN U13424 ( .B(n1834), .A(n1835), .Z(n1832) );
  AND U13425 ( .A(a[95]), .B(b[30]), .Z(n1831) );
  XOR U13426 ( .A(n1836), .B(n908), .Z(n910) );
  XOR U13427 ( .A(n1837), .B(n1838), .Z(n908) );
  ANDN U13428 ( .B(n1839), .A(n1840), .Z(n1837) );
  AND U13429 ( .A(a[96]), .B(b[29]), .Z(n1836) );
  XOR U13430 ( .A(n1841), .B(n1069), .Z(n1064) );
  XOR U13431 ( .A(n1842), .B(n1843), .Z(n1069) );
  ANDN U13432 ( .B(n1844), .A(n1845), .Z(n1842) );
  AND U13433 ( .A(a[97]), .B(b[28]), .Z(n1841) );
  XOR U13434 ( .A(n1846), .B(n1066), .Z(n1060) );
  XOR U13435 ( .A(n1847), .B(n1848), .Z(n1066) );
  ANDN U13436 ( .B(n1849), .A(n1850), .Z(n1847) );
  AND U13437 ( .A(a[98]), .B(b[27]), .Z(n1846) );
  XOR U13438 ( .A(n1851), .B(n1062), .Z(n1056) );
  XOR U13439 ( .A(n1852), .B(n1853), .Z(n1062) );
  ANDN U13440 ( .B(n1854), .A(n1855), .Z(n1852) );
  AND U13441 ( .A(a[99]), .B(b[26]), .Z(n1851) );
  XOR U13442 ( .A(n1856), .B(n1058), .Z(n1053) );
  XOR U13443 ( .A(n1857), .B(n1858), .Z(n1058) );
  ANDN U13444 ( .B(n1859), .A(n1860), .Z(n1857) );
  AND U13445 ( .A(b[25]), .B(a[100]), .Z(n1856) );
  XNOR U13446 ( .A(n1861), .B(n912), .Z(n913) );
  XOR U13447 ( .A(n1862), .B(n1863), .Z(n912) );
  ANDN U13448 ( .B(n1864), .A(n1865), .Z(n1862) );
  AND U13449 ( .A(b[24]), .B(a[101]), .Z(n1861) );
  XOR U13450 ( .A(n1866), .B(n922), .Z(n924) );
  XOR U13451 ( .A(n1867), .B(n1868), .Z(n922) );
  ANDN U13452 ( .B(n1869), .A(n1870), .Z(n1867) );
  AND U13453 ( .A(b[23]), .B(a[102]), .Z(n1866) );
  XOR U13454 ( .A(n1871), .B(n1051), .Z(n1046) );
  XOR U13455 ( .A(n1872), .B(n1873), .Z(n1051) );
  ANDN U13456 ( .B(n1874), .A(n1875), .Z(n1872) );
  AND U13457 ( .A(b[22]), .B(a[103]), .Z(n1871) );
  XOR U13458 ( .A(n1876), .B(n1048), .Z(n1042) );
  XOR U13459 ( .A(n1877), .B(n1878), .Z(n1048) );
  ANDN U13460 ( .B(n1879), .A(n1880), .Z(n1877) );
  AND U13461 ( .A(b[21]), .B(a[104]), .Z(n1876) );
  XOR U13462 ( .A(n1881), .B(n1044), .Z(n1038) );
  XOR U13463 ( .A(n1882), .B(n1883), .Z(n1044) );
  ANDN U13464 ( .B(n1884), .A(n1885), .Z(n1882) );
  AND U13465 ( .A(b[20]), .B(a[105]), .Z(n1881) );
  XOR U13466 ( .A(n1886), .B(n1040), .Z(n1035) );
  XOR U13467 ( .A(n1887), .B(n1888), .Z(n1040) );
  ANDN U13468 ( .B(n1889), .A(n1890), .Z(n1887) );
  AND U13469 ( .A(b[19]), .B(a[106]), .Z(n1886) );
  XNOR U13470 ( .A(n1891), .B(n926), .Z(n927) );
  XOR U13471 ( .A(n1892), .B(n1893), .Z(n926) );
  ANDN U13472 ( .B(n1894), .A(n1895), .Z(n1892) );
  AND U13473 ( .A(b[18]), .B(a[107]), .Z(n1891) );
  XOR U13474 ( .A(n1896), .B(n936), .Z(n938) );
  XOR U13475 ( .A(n1897), .B(n1898), .Z(n936) );
  ANDN U13476 ( .B(n1899), .A(n1900), .Z(n1897) );
  AND U13477 ( .A(b[17]), .B(a[108]), .Z(n1896) );
  XOR U13478 ( .A(n1901), .B(n1033), .Z(n1028) );
  XOR U13479 ( .A(n1902), .B(n1903), .Z(n1033) );
  ANDN U13480 ( .B(n1904), .A(n1905), .Z(n1902) );
  AND U13481 ( .A(b[16]), .B(a[109]), .Z(n1901) );
  XOR U13482 ( .A(n1906), .B(n1030), .Z(n1024) );
  XOR U13483 ( .A(n1907), .B(n1908), .Z(n1030) );
  ANDN U13484 ( .B(n1909), .A(n1910), .Z(n1907) );
  AND U13485 ( .A(b[15]), .B(a[110]), .Z(n1906) );
  XOR U13486 ( .A(n1911), .B(n1026), .Z(n1020) );
  XOR U13487 ( .A(n1912), .B(n1913), .Z(n1026) );
  ANDN U13488 ( .B(n1914), .A(n1915), .Z(n1912) );
  AND U13489 ( .A(b[14]), .B(a[111]), .Z(n1911) );
  XOR U13490 ( .A(n1916), .B(n1022), .Z(n1017) );
  XOR U13491 ( .A(n1917), .B(n1918), .Z(n1022) );
  ANDN U13492 ( .B(n1919), .A(n1920), .Z(n1917) );
  AND U13493 ( .A(b[13]), .B(a[112]), .Z(n1916) );
  XOR U13494 ( .A(n1921), .B(n940), .Z(n941) );
  XOR U13495 ( .A(n1922), .B(n1923), .Z(n940) );
  ANDN U13496 ( .B(n1924), .A(n1925), .Z(n1922) );
  AND U13497 ( .A(b[12]), .B(a[113]), .Z(n1921) );
  XOR U13498 ( .A(n1926), .B(n1016), .Z(n1011) );
  XOR U13499 ( .A(n1927), .B(n1928), .Z(n1016) );
  ANDN U13500 ( .B(n1929), .A(n1930), .Z(n1927) );
  AND U13501 ( .A(b[11]), .B(a[114]), .Z(n1926) );
  XOR U13502 ( .A(n1931), .B(n1013), .Z(n1007) );
  XOR U13503 ( .A(n1932), .B(n1933), .Z(n1013) );
  ANDN U13504 ( .B(n1934), .A(n1935), .Z(n1932) );
  AND U13505 ( .A(b[10]), .B(a[115]), .Z(n1931) );
  XOR U13506 ( .A(n1936), .B(n1009), .Z(n1003) );
  XOR U13507 ( .A(n1937), .B(n1938), .Z(n1009) );
  ANDN U13508 ( .B(n1939), .A(n1940), .Z(n1937) );
  AND U13509 ( .A(b[9]), .B(a[116]), .Z(n1936) );
  XOR U13510 ( .A(n1941), .B(n1005), .Z(n999) );
  XOR U13511 ( .A(n1942), .B(n1943), .Z(n1005) );
  ANDN U13512 ( .B(n1944), .A(n1945), .Z(n1942) );
  AND U13513 ( .A(b[8]), .B(a[117]), .Z(n1941) );
  XOR U13514 ( .A(n1946), .B(n1001), .Z(n996) );
  XOR U13515 ( .A(n1947), .B(n1948), .Z(n1001) );
  ANDN U13516 ( .B(n1949), .A(n1950), .Z(n1947) );
  AND U13517 ( .A(b[7]), .B(a[118]), .Z(n1946) );
  XOR U13518 ( .A(n1951), .B(n951), .Z(n952) );
  XOR U13519 ( .A(n1952), .B(n1953), .Z(n951) );
  ANDN U13520 ( .B(n1954), .A(n1955), .Z(n1952) );
  AND U13521 ( .A(b[6]), .B(a[119]), .Z(n1951) );
  XOR U13522 ( .A(n1956), .B(n995), .Z(n990) );
  XOR U13523 ( .A(n1957), .B(n1958), .Z(n995) );
  ANDN U13524 ( .B(n1959), .A(n1960), .Z(n1957) );
  AND U13525 ( .A(b[5]), .B(a[120]), .Z(n1956) );
  XOR U13526 ( .A(n1961), .B(n992), .Z(n986) );
  XOR U13527 ( .A(n1962), .B(n1963), .Z(n992) );
  ANDN U13528 ( .B(n1964), .A(n1965), .Z(n1962) );
  AND U13529 ( .A(b[4]), .B(a[121]), .Z(n1961) );
  XNOR U13530 ( .A(n1966), .B(n1967), .Z(n980) );
  NANDN U13531 ( .A(n1968), .B(n1969), .Z(n1967) );
  XOR U13532 ( .A(n1970), .B(n988), .Z(n983) );
  XNOR U13533 ( .A(n1971), .B(n1972), .Z(n988) );
  AND U13534 ( .A(n1973), .B(n1974), .Z(n1971) );
  AND U13535 ( .A(b[3]), .B(a[122]), .Z(n1970) );
  NAND U13536 ( .A(a[125]), .B(b[0]), .Z(n973) );
  XNOR U13537 ( .A(n982), .B(n981), .Z(c[124]) );
  XNOR U13538 ( .A(n1968), .B(n1969), .Z(n981) );
  XOR U13539 ( .A(n1966), .B(n1975), .Z(n1969) );
  NAND U13540 ( .A(b[1]), .B(a[123]), .Z(n1975) );
  XOR U13541 ( .A(n1974), .B(n1976), .Z(n1968) );
  XOR U13542 ( .A(n1966), .B(n1973), .Z(n1976) );
  XNOR U13543 ( .A(n1977), .B(n1972), .Z(n1973) );
  AND U13544 ( .A(b[2]), .B(a[122]), .Z(n1977) );
  NANDN U13545 ( .A(n1978), .B(n1979), .Z(n1966) );
  XOR U13546 ( .A(n1972), .B(n1964), .Z(n1980) );
  XNOR U13547 ( .A(n1963), .B(n1959), .Z(n1981) );
  XNOR U13548 ( .A(n1958), .B(n1954), .Z(n1982) );
  XNOR U13549 ( .A(n1953), .B(n1949), .Z(n1983) );
  XNOR U13550 ( .A(n1948), .B(n1944), .Z(n1984) );
  XNOR U13551 ( .A(n1943), .B(n1939), .Z(n1985) );
  XNOR U13552 ( .A(n1938), .B(n1934), .Z(n1986) );
  XNOR U13553 ( .A(n1933), .B(n1929), .Z(n1987) );
  XNOR U13554 ( .A(n1928), .B(n1924), .Z(n1988) );
  XNOR U13555 ( .A(n1923), .B(n1919), .Z(n1989) );
  XNOR U13556 ( .A(n1918), .B(n1914), .Z(n1990) );
  XNOR U13557 ( .A(n1913), .B(n1909), .Z(n1991) );
  XNOR U13558 ( .A(n1908), .B(n1904), .Z(n1992) );
  XNOR U13559 ( .A(n1903), .B(n1899), .Z(n1993) );
  XNOR U13560 ( .A(n1898), .B(n1894), .Z(n1994) );
  XNOR U13561 ( .A(n1893), .B(n1889), .Z(n1995) );
  XNOR U13562 ( .A(n1888), .B(n1884), .Z(n1996) );
  XNOR U13563 ( .A(n1883), .B(n1879), .Z(n1997) );
  XNOR U13564 ( .A(n1878), .B(n1874), .Z(n1998) );
  XNOR U13565 ( .A(n1873), .B(n1869), .Z(n1999) );
  XNOR U13566 ( .A(n1868), .B(n1864), .Z(n2000) );
  XNOR U13567 ( .A(n1863), .B(n1859), .Z(n2001) );
  XNOR U13568 ( .A(n1858), .B(n1854), .Z(n2002) );
  XNOR U13569 ( .A(n1853), .B(n1849), .Z(n2003) );
  XNOR U13570 ( .A(n1848), .B(n1844), .Z(n2004) );
  XNOR U13571 ( .A(n1843), .B(n1839), .Z(n2005) );
  XNOR U13572 ( .A(n1838), .B(n1834), .Z(n2006) );
  XNOR U13573 ( .A(n1833), .B(n1829), .Z(n2007) );
  XNOR U13574 ( .A(n1828), .B(n1824), .Z(n2008) );
  XNOR U13575 ( .A(n1823), .B(n1819), .Z(n2009) );
  XNOR U13576 ( .A(n1818), .B(n1814), .Z(n2010) );
  XNOR U13577 ( .A(n1813), .B(n1809), .Z(n2011) );
  XNOR U13578 ( .A(n1808), .B(n1804), .Z(n2012) );
  XNOR U13579 ( .A(n1803), .B(n1799), .Z(n2013) );
  XNOR U13580 ( .A(n1798), .B(n1794), .Z(n2014) );
  XNOR U13581 ( .A(n1793), .B(n1789), .Z(n2015) );
  XNOR U13582 ( .A(n1788), .B(n1784), .Z(n2016) );
  XNOR U13583 ( .A(n1783), .B(n1779), .Z(n2017) );
  XNOR U13584 ( .A(n1778), .B(n1774), .Z(n2018) );
  XNOR U13585 ( .A(n1773), .B(n1769), .Z(n2019) );
  XNOR U13586 ( .A(n1768), .B(n1764), .Z(n2020) );
  XNOR U13587 ( .A(n1763), .B(n1759), .Z(n2021) );
  XNOR U13588 ( .A(n1758), .B(n1754), .Z(n2022) );
  XNOR U13589 ( .A(n1753), .B(n1749), .Z(n2023) );
  XNOR U13590 ( .A(n1748), .B(n1744), .Z(n2024) );
  XNOR U13591 ( .A(n1743), .B(n1739), .Z(n2025) );
  XNOR U13592 ( .A(n1738), .B(n1734), .Z(n2026) );
  XNOR U13593 ( .A(n1733), .B(n1729), .Z(n2027) );
  XNOR U13594 ( .A(n1728), .B(n1724), .Z(n2028) );
  XNOR U13595 ( .A(n1723), .B(n1719), .Z(n2029) );
  XNOR U13596 ( .A(n1718), .B(n1714), .Z(n2030) );
  XNOR U13597 ( .A(n1713), .B(n1709), .Z(n2031) );
  XNOR U13598 ( .A(n1708), .B(n1704), .Z(n2032) );
  XNOR U13599 ( .A(n1703), .B(n1699), .Z(n2033) );
  XNOR U13600 ( .A(n1698), .B(n1694), .Z(n2034) );
  XNOR U13601 ( .A(n1693), .B(n1689), .Z(n2035) );
  XNOR U13602 ( .A(n1688), .B(n1684), .Z(n2036) );
  XNOR U13603 ( .A(n1683), .B(n1679), .Z(n2037) );
  XNOR U13604 ( .A(n1678), .B(n1674), .Z(n2038) );
  XNOR U13605 ( .A(n1673), .B(n1669), .Z(n2039) );
  XNOR U13606 ( .A(n1668), .B(n1664), .Z(n2040) );
  XNOR U13607 ( .A(n1663), .B(n1659), .Z(n2041) );
  XNOR U13608 ( .A(n1658), .B(n1654), .Z(n2042) );
  XNOR U13609 ( .A(n1653), .B(n1649), .Z(n2043) );
  XNOR U13610 ( .A(n1648), .B(n1644), .Z(n2044) );
  XNOR U13611 ( .A(n1643), .B(n1639), .Z(n2045) );
  XNOR U13612 ( .A(n1638), .B(n1634), .Z(n2046) );
  XNOR U13613 ( .A(n1633), .B(n1629), .Z(n2047) );
  XNOR U13614 ( .A(n1628), .B(n1624), .Z(n2048) );
  XNOR U13615 ( .A(n1623), .B(n1619), .Z(n2049) );
  XNOR U13616 ( .A(n1618), .B(n1614), .Z(n2050) );
  XNOR U13617 ( .A(n1613), .B(n1609), .Z(n2051) );
  XNOR U13618 ( .A(n1608), .B(n1604), .Z(n2052) );
  XNOR U13619 ( .A(n1603), .B(n1599), .Z(n2053) );
  XNOR U13620 ( .A(n1598), .B(n1594), .Z(n2054) );
  XNOR U13621 ( .A(n1593), .B(n1589), .Z(n2055) );
  XNOR U13622 ( .A(n1588), .B(n1584), .Z(n2056) );
  XNOR U13623 ( .A(n1583), .B(n1579), .Z(n2057) );
  XNOR U13624 ( .A(n1578), .B(n1574), .Z(n2058) );
  XNOR U13625 ( .A(n1573), .B(n1569), .Z(n2059) );
  XNOR U13626 ( .A(n1568), .B(n1564), .Z(n2060) );
  XNOR U13627 ( .A(n1563), .B(n1559), .Z(n2061) );
  XNOR U13628 ( .A(n1558), .B(n1554), .Z(n2062) );
  XNOR U13629 ( .A(n1553), .B(n1549), .Z(n2063) );
  XNOR U13630 ( .A(n1548), .B(n1544), .Z(n2064) );
  XNOR U13631 ( .A(n1543), .B(n1539), .Z(n2065) );
  XNOR U13632 ( .A(n1538), .B(n1534), .Z(n2066) );
  XNOR U13633 ( .A(n1533), .B(n1529), .Z(n2067) );
  XNOR U13634 ( .A(n1528), .B(n1524), .Z(n2068) );
  XNOR U13635 ( .A(n1523), .B(n1519), .Z(n2069) );
  XNOR U13636 ( .A(n1518), .B(n1514), .Z(n2070) );
  XNOR U13637 ( .A(n1513), .B(n1509), .Z(n2071) );
  XNOR U13638 ( .A(n1508), .B(n1504), .Z(n2072) );
  XNOR U13639 ( .A(n1503), .B(n1499), .Z(n2073) );
  XNOR U13640 ( .A(n1498), .B(n1494), .Z(n2074) );
  XNOR U13641 ( .A(n1493), .B(n1489), .Z(n2075) );
  XNOR U13642 ( .A(n1488), .B(n1484), .Z(n2076) );
  XNOR U13643 ( .A(n1483), .B(n1479), .Z(n2077) );
  XNOR U13644 ( .A(n1478), .B(n1474), .Z(n2078) );
  XNOR U13645 ( .A(n1473), .B(n1469), .Z(n2079) );
  XNOR U13646 ( .A(n1468), .B(n1464), .Z(n2080) );
  XNOR U13647 ( .A(n1463), .B(n1459), .Z(n2081) );
  XNOR U13648 ( .A(n1458), .B(n1454), .Z(n2082) );
  XNOR U13649 ( .A(n1453), .B(n1449), .Z(n2083) );
  XNOR U13650 ( .A(n1448), .B(n1444), .Z(n2084) );
  XNOR U13651 ( .A(n1443), .B(n1439), .Z(n2085) );
  XNOR U13652 ( .A(n1438), .B(n1434), .Z(n2086) );
  XNOR U13653 ( .A(n1433), .B(n1429), .Z(n2087) );
  XNOR U13654 ( .A(n1428), .B(n1424), .Z(n2088) );
  XNOR U13655 ( .A(n1423), .B(n1419), .Z(n2089) );
  XNOR U13656 ( .A(n1418), .B(n1414), .Z(n2090) );
  XNOR U13657 ( .A(n1413), .B(n1409), .Z(n2091) );
  XNOR U13658 ( .A(n1408), .B(n1404), .Z(n2092) );
  XNOR U13659 ( .A(n1403), .B(n1399), .Z(n2093) );
  XNOR U13660 ( .A(n1398), .B(n1394), .Z(n2094) );
  XNOR U13661 ( .A(n1393), .B(n1389), .Z(n2095) );
  XNOR U13662 ( .A(n1388), .B(n1384), .Z(n2096) );
  XNOR U13663 ( .A(n1383), .B(n1379), .Z(n2097) );
  XNOR U13664 ( .A(n1378), .B(n1374), .Z(n2098) );
  XNOR U13665 ( .A(n1373), .B(n1369), .Z(n2099) );
  XNOR U13666 ( .A(n1368), .B(n1364), .Z(n2100) );
  XOR U13667 ( .A(n2101), .B(n1363), .Z(n1364) );
  AND U13668 ( .A(a[0]), .B(b[124]), .Z(n2101) );
  XNOR U13669 ( .A(n2102), .B(n1363), .Z(n1365) );
  XNOR U13670 ( .A(n2103), .B(n2104), .Z(n1363) );
  ANDN U13671 ( .B(n2105), .A(n2106), .Z(n2103) );
  AND U13672 ( .A(a[1]), .B(b[123]), .Z(n2102) );
  XNOR U13673 ( .A(n2107), .B(n1368), .Z(n1370) );
  XOR U13674 ( .A(n2108), .B(n2109), .Z(n1368) );
  ANDN U13675 ( .B(n2110), .A(n2111), .Z(n2108) );
  AND U13676 ( .A(a[2]), .B(b[122]), .Z(n2107) );
  XNOR U13677 ( .A(n2112), .B(n1373), .Z(n1375) );
  XOR U13678 ( .A(n2113), .B(n2114), .Z(n1373) );
  ANDN U13679 ( .B(n2115), .A(n2116), .Z(n2113) );
  AND U13680 ( .A(a[3]), .B(b[121]), .Z(n2112) );
  XNOR U13681 ( .A(n2117), .B(n1378), .Z(n1380) );
  XOR U13682 ( .A(n2118), .B(n2119), .Z(n1378) );
  ANDN U13683 ( .B(n2120), .A(n2121), .Z(n2118) );
  AND U13684 ( .A(a[4]), .B(b[120]), .Z(n2117) );
  XNOR U13685 ( .A(n2122), .B(n1383), .Z(n1385) );
  XOR U13686 ( .A(n2123), .B(n2124), .Z(n1383) );
  ANDN U13687 ( .B(n2125), .A(n2126), .Z(n2123) );
  AND U13688 ( .A(a[5]), .B(b[119]), .Z(n2122) );
  XNOR U13689 ( .A(n2127), .B(n1388), .Z(n1390) );
  XOR U13690 ( .A(n2128), .B(n2129), .Z(n1388) );
  ANDN U13691 ( .B(n2130), .A(n2131), .Z(n2128) );
  AND U13692 ( .A(a[6]), .B(b[118]), .Z(n2127) );
  XNOR U13693 ( .A(n2132), .B(n1393), .Z(n1395) );
  XOR U13694 ( .A(n2133), .B(n2134), .Z(n1393) );
  ANDN U13695 ( .B(n2135), .A(n2136), .Z(n2133) );
  AND U13696 ( .A(a[7]), .B(b[117]), .Z(n2132) );
  XNOR U13697 ( .A(n2137), .B(n1398), .Z(n1400) );
  XOR U13698 ( .A(n2138), .B(n2139), .Z(n1398) );
  ANDN U13699 ( .B(n2140), .A(n2141), .Z(n2138) );
  AND U13700 ( .A(a[8]), .B(b[116]), .Z(n2137) );
  XNOR U13701 ( .A(n2142), .B(n1403), .Z(n1405) );
  XOR U13702 ( .A(n2143), .B(n2144), .Z(n1403) );
  ANDN U13703 ( .B(n2145), .A(n2146), .Z(n2143) );
  AND U13704 ( .A(a[9]), .B(b[115]), .Z(n2142) );
  XNOR U13705 ( .A(n2147), .B(n1408), .Z(n1410) );
  XOR U13706 ( .A(n2148), .B(n2149), .Z(n1408) );
  ANDN U13707 ( .B(n2150), .A(n2151), .Z(n2148) );
  AND U13708 ( .A(a[10]), .B(b[114]), .Z(n2147) );
  XNOR U13709 ( .A(n2152), .B(n1413), .Z(n1415) );
  XOR U13710 ( .A(n2153), .B(n2154), .Z(n1413) );
  ANDN U13711 ( .B(n2155), .A(n2156), .Z(n2153) );
  AND U13712 ( .A(a[11]), .B(b[113]), .Z(n2152) );
  XNOR U13713 ( .A(n2157), .B(n1418), .Z(n1420) );
  XOR U13714 ( .A(n2158), .B(n2159), .Z(n1418) );
  ANDN U13715 ( .B(n2160), .A(n2161), .Z(n2158) );
  AND U13716 ( .A(a[12]), .B(b[112]), .Z(n2157) );
  XNOR U13717 ( .A(n2162), .B(n1423), .Z(n1425) );
  XOR U13718 ( .A(n2163), .B(n2164), .Z(n1423) );
  ANDN U13719 ( .B(n2165), .A(n2166), .Z(n2163) );
  AND U13720 ( .A(a[13]), .B(b[111]), .Z(n2162) );
  XNOR U13721 ( .A(n2167), .B(n1428), .Z(n1430) );
  XOR U13722 ( .A(n2168), .B(n2169), .Z(n1428) );
  ANDN U13723 ( .B(n2170), .A(n2171), .Z(n2168) );
  AND U13724 ( .A(a[14]), .B(b[110]), .Z(n2167) );
  XNOR U13725 ( .A(n2172), .B(n1433), .Z(n1435) );
  XOR U13726 ( .A(n2173), .B(n2174), .Z(n1433) );
  ANDN U13727 ( .B(n2175), .A(n2176), .Z(n2173) );
  AND U13728 ( .A(a[15]), .B(b[109]), .Z(n2172) );
  XNOR U13729 ( .A(n2177), .B(n1438), .Z(n1440) );
  XOR U13730 ( .A(n2178), .B(n2179), .Z(n1438) );
  ANDN U13731 ( .B(n2180), .A(n2181), .Z(n2178) );
  AND U13732 ( .A(a[16]), .B(b[108]), .Z(n2177) );
  XNOR U13733 ( .A(n2182), .B(n1443), .Z(n1445) );
  XOR U13734 ( .A(n2183), .B(n2184), .Z(n1443) );
  ANDN U13735 ( .B(n2185), .A(n2186), .Z(n2183) );
  AND U13736 ( .A(a[17]), .B(b[107]), .Z(n2182) );
  XNOR U13737 ( .A(n2187), .B(n1448), .Z(n1450) );
  XOR U13738 ( .A(n2188), .B(n2189), .Z(n1448) );
  ANDN U13739 ( .B(n2190), .A(n2191), .Z(n2188) );
  AND U13740 ( .A(a[18]), .B(b[106]), .Z(n2187) );
  XNOR U13741 ( .A(n2192), .B(n1453), .Z(n1455) );
  XOR U13742 ( .A(n2193), .B(n2194), .Z(n1453) );
  ANDN U13743 ( .B(n2195), .A(n2196), .Z(n2193) );
  AND U13744 ( .A(a[19]), .B(b[105]), .Z(n2192) );
  XNOR U13745 ( .A(n2197), .B(n1458), .Z(n1460) );
  XOR U13746 ( .A(n2198), .B(n2199), .Z(n1458) );
  ANDN U13747 ( .B(n2200), .A(n2201), .Z(n2198) );
  AND U13748 ( .A(a[20]), .B(b[104]), .Z(n2197) );
  XNOR U13749 ( .A(n2202), .B(n1463), .Z(n1465) );
  XOR U13750 ( .A(n2203), .B(n2204), .Z(n1463) );
  ANDN U13751 ( .B(n2205), .A(n2206), .Z(n2203) );
  AND U13752 ( .A(a[21]), .B(b[103]), .Z(n2202) );
  XNOR U13753 ( .A(n2207), .B(n1468), .Z(n1470) );
  XOR U13754 ( .A(n2208), .B(n2209), .Z(n1468) );
  ANDN U13755 ( .B(n2210), .A(n2211), .Z(n2208) );
  AND U13756 ( .A(a[22]), .B(b[102]), .Z(n2207) );
  XNOR U13757 ( .A(n2212), .B(n1473), .Z(n1475) );
  XOR U13758 ( .A(n2213), .B(n2214), .Z(n1473) );
  ANDN U13759 ( .B(n2215), .A(n2216), .Z(n2213) );
  AND U13760 ( .A(a[23]), .B(b[101]), .Z(n2212) );
  XNOR U13761 ( .A(n2217), .B(n1478), .Z(n1480) );
  XOR U13762 ( .A(n2218), .B(n2219), .Z(n1478) );
  ANDN U13763 ( .B(n2220), .A(n2221), .Z(n2218) );
  AND U13764 ( .A(a[24]), .B(b[100]), .Z(n2217) );
  XNOR U13765 ( .A(n2222), .B(n1483), .Z(n1485) );
  XOR U13766 ( .A(n2223), .B(n2224), .Z(n1483) );
  ANDN U13767 ( .B(n2225), .A(n2226), .Z(n2223) );
  AND U13768 ( .A(a[25]), .B(b[99]), .Z(n2222) );
  XNOR U13769 ( .A(n2227), .B(n1488), .Z(n1490) );
  XOR U13770 ( .A(n2228), .B(n2229), .Z(n1488) );
  ANDN U13771 ( .B(n2230), .A(n2231), .Z(n2228) );
  AND U13772 ( .A(a[26]), .B(b[98]), .Z(n2227) );
  XNOR U13773 ( .A(n2232), .B(n1493), .Z(n1495) );
  XOR U13774 ( .A(n2233), .B(n2234), .Z(n1493) );
  ANDN U13775 ( .B(n2235), .A(n2236), .Z(n2233) );
  AND U13776 ( .A(a[27]), .B(b[97]), .Z(n2232) );
  XNOR U13777 ( .A(n2237), .B(n1498), .Z(n1500) );
  XOR U13778 ( .A(n2238), .B(n2239), .Z(n1498) );
  ANDN U13779 ( .B(n2240), .A(n2241), .Z(n2238) );
  AND U13780 ( .A(a[28]), .B(b[96]), .Z(n2237) );
  XNOR U13781 ( .A(n2242), .B(n1503), .Z(n1505) );
  XOR U13782 ( .A(n2243), .B(n2244), .Z(n1503) );
  ANDN U13783 ( .B(n2245), .A(n2246), .Z(n2243) );
  AND U13784 ( .A(a[29]), .B(b[95]), .Z(n2242) );
  XNOR U13785 ( .A(n2247), .B(n1508), .Z(n1510) );
  XOR U13786 ( .A(n2248), .B(n2249), .Z(n1508) );
  ANDN U13787 ( .B(n2250), .A(n2251), .Z(n2248) );
  AND U13788 ( .A(a[30]), .B(b[94]), .Z(n2247) );
  XNOR U13789 ( .A(n2252), .B(n1513), .Z(n1515) );
  XOR U13790 ( .A(n2253), .B(n2254), .Z(n1513) );
  ANDN U13791 ( .B(n2255), .A(n2256), .Z(n2253) );
  AND U13792 ( .A(a[31]), .B(b[93]), .Z(n2252) );
  XNOR U13793 ( .A(n2257), .B(n1518), .Z(n1520) );
  XOR U13794 ( .A(n2258), .B(n2259), .Z(n1518) );
  ANDN U13795 ( .B(n2260), .A(n2261), .Z(n2258) );
  AND U13796 ( .A(a[32]), .B(b[92]), .Z(n2257) );
  XNOR U13797 ( .A(n2262), .B(n1523), .Z(n1525) );
  XOR U13798 ( .A(n2263), .B(n2264), .Z(n1523) );
  ANDN U13799 ( .B(n2265), .A(n2266), .Z(n2263) );
  AND U13800 ( .A(a[33]), .B(b[91]), .Z(n2262) );
  XNOR U13801 ( .A(n2267), .B(n1528), .Z(n1530) );
  XOR U13802 ( .A(n2268), .B(n2269), .Z(n1528) );
  ANDN U13803 ( .B(n2270), .A(n2271), .Z(n2268) );
  AND U13804 ( .A(a[34]), .B(b[90]), .Z(n2267) );
  XNOR U13805 ( .A(n2272), .B(n1533), .Z(n1535) );
  XOR U13806 ( .A(n2273), .B(n2274), .Z(n1533) );
  ANDN U13807 ( .B(n2275), .A(n2276), .Z(n2273) );
  AND U13808 ( .A(a[35]), .B(b[89]), .Z(n2272) );
  XNOR U13809 ( .A(n2277), .B(n1538), .Z(n1540) );
  XOR U13810 ( .A(n2278), .B(n2279), .Z(n1538) );
  ANDN U13811 ( .B(n2280), .A(n2281), .Z(n2278) );
  AND U13812 ( .A(a[36]), .B(b[88]), .Z(n2277) );
  XNOR U13813 ( .A(n2282), .B(n1543), .Z(n1545) );
  XOR U13814 ( .A(n2283), .B(n2284), .Z(n1543) );
  ANDN U13815 ( .B(n2285), .A(n2286), .Z(n2283) );
  AND U13816 ( .A(a[37]), .B(b[87]), .Z(n2282) );
  XNOR U13817 ( .A(n2287), .B(n1548), .Z(n1550) );
  XOR U13818 ( .A(n2288), .B(n2289), .Z(n1548) );
  ANDN U13819 ( .B(n2290), .A(n2291), .Z(n2288) );
  AND U13820 ( .A(a[38]), .B(b[86]), .Z(n2287) );
  XNOR U13821 ( .A(n2292), .B(n1553), .Z(n1555) );
  XOR U13822 ( .A(n2293), .B(n2294), .Z(n1553) );
  ANDN U13823 ( .B(n2295), .A(n2296), .Z(n2293) );
  AND U13824 ( .A(a[39]), .B(b[85]), .Z(n2292) );
  XNOR U13825 ( .A(n2297), .B(n1558), .Z(n1560) );
  XOR U13826 ( .A(n2298), .B(n2299), .Z(n1558) );
  ANDN U13827 ( .B(n2300), .A(n2301), .Z(n2298) );
  AND U13828 ( .A(a[40]), .B(b[84]), .Z(n2297) );
  XNOR U13829 ( .A(n2302), .B(n1563), .Z(n1565) );
  XOR U13830 ( .A(n2303), .B(n2304), .Z(n1563) );
  ANDN U13831 ( .B(n2305), .A(n2306), .Z(n2303) );
  AND U13832 ( .A(a[41]), .B(b[83]), .Z(n2302) );
  XNOR U13833 ( .A(n2307), .B(n1568), .Z(n1570) );
  XOR U13834 ( .A(n2308), .B(n2309), .Z(n1568) );
  ANDN U13835 ( .B(n2310), .A(n2311), .Z(n2308) );
  AND U13836 ( .A(a[42]), .B(b[82]), .Z(n2307) );
  XNOR U13837 ( .A(n2312), .B(n1573), .Z(n1575) );
  XOR U13838 ( .A(n2313), .B(n2314), .Z(n1573) );
  ANDN U13839 ( .B(n2315), .A(n2316), .Z(n2313) );
  AND U13840 ( .A(a[43]), .B(b[81]), .Z(n2312) );
  XNOR U13841 ( .A(n2317), .B(n1578), .Z(n1580) );
  XOR U13842 ( .A(n2318), .B(n2319), .Z(n1578) );
  ANDN U13843 ( .B(n2320), .A(n2321), .Z(n2318) );
  AND U13844 ( .A(a[44]), .B(b[80]), .Z(n2317) );
  XNOR U13845 ( .A(n2322), .B(n1583), .Z(n1585) );
  XOR U13846 ( .A(n2323), .B(n2324), .Z(n1583) );
  ANDN U13847 ( .B(n2325), .A(n2326), .Z(n2323) );
  AND U13848 ( .A(a[45]), .B(b[79]), .Z(n2322) );
  XNOR U13849 ( .A(n2327), .B(n1588), .Z(n1590) );
  XOR U13850 ( .A(n2328), .B(n2329), .Z(n1588) );
  ANDN U13851 ( .B(n2330), .A(n2331), .Z(n2328) );
  AND U13852 ( .A(a[46]), .B(b[78]), .Z(n2327) );
  XNOR U13853 ( .A(n2332), .B(n1593), .Z(n1595) );
  XOR U13854 ( .A(n2333), .B(n2334), .Z(n1593) );
  ANDN U13855 ( .B(n2335), .A(n2336), .Z(n2333) );
  AND U13856 ( .A(a[47]), .B(b[77]), .Z(n2332) );
  XNOR U13857 ( .A(n2337), .B(n1598), .Z(n1600) );
  XOR U13858 ( .A(n2338), .B(n2339), .Z(n1598) );
  ANDN U13859 ( .B(n2340), .A(n2341), .Z(n2338) );
  AND U13860 ( .A(a[48]), .B(b[76]), .Z(n2337) );
  XNOR U13861 ( .A(n2342), .B(n1603), .Z(n1605) );
  XOR U13862 ( .A(n2343), .B(n2344), .Z(n1603) );
  ANDN U13863 ( .B(n2345), .A(n2346), .Z(n2343) );
  AND U13864 ( .A(a[49]), .B(b[75]), .Z(n2342) );
  XNOR U13865 ( .A(n2347), .B(n1608), .Z(n1610) );
  XOR U13866 ( .A(n2348), .B(n2349), .Z(n1608) );
  ANDN U13867 ( .B(n2350), .A(n2351), .Z(n2348) );
  AND U13868 ( .A(a[50]), .B(b[74]), .Z(n2347) );
  XNOR U13869 ( .A(n2352), .B(n1613), .Z(n1615) );
  XOR U13870 ( .A(n2353), .B(n2354), .Z(n1613) );
  ANDN U13871 ( .B(n2355), .A(n2356), .Z(n2353) );
  AND U13872 ( .A(a[51]), .B(b[73]), .Z(n2352) );
  XNOR U13873 ( .A(n2357), .B(n1618), .Z(n1620) );
  XOR U13874 ( .A(n2358), .B(n2359), .Z(n1618) );
  ANDN U13875 ( .B(n2360), .A(n2361), .Z(n2358) );
  AND U13876 ( .A(a[52]), .B(b[72]), .Z(n2357) );
  XNOR U13877 ( .A(n2362), .B(n1623), .Z(n1625) );
  XOR U13878 ( .A(n2363), .B(n2364), .Z(n1623) );
  ANDN U13879 ( .B(n2365), .A(n2366), .Z(n2363) );
  AND U13880 ( .A(a[53]), .B(b[71]), .Z(n2362) );
  XNOR U13881 ( .A(n2367), .B(n1628), .Z(n1630) );
  XOR U13882 ( .A(n2368), .B(n2369), .Z(n1628) );
  ANDN U13883 ( .B(n2370), .A(n2371), .Z(n2368) );
  AND U13884 ( .A(a[54]), .B(b[70]), .Z(n2367) );
  XNOR U13885 ( .A(n2372), .B(n1633), .Z(n1635) );
  XOR U13886 ( .A(n2373), .B(n2374), .Z(n1633) );
  ANDN U13887 ( .B(n2375), .A(n2376), .Z(n2373) );
  AND U13888 ( .A(a[55]), .B(b[69]), .Z(n2372) );
  XNOR U13889 ( .A(n2377), .B(n1638), .Z(n1640) );
  XOR U13890 ( .A(n2378), .B(n2379), .Z(n1638) );
  ANDN U13891 ( .B(n2380), .A(n2381), .Z(n2378) );
  AND U13892 ( .A(a[56]), .B(b[68]), .Z(n2377) );
  XNOR U13893 ( .A(n2382), .B(n1643), .Z(n1645) );
  XOR U13894 ( .A(n2383), .B(n2384), .Z(n1643) );
  ANDN U13895 ( .B(n2385), .A(n2386), .Z(n2383) );
  AND U13896 ( .A(a[57]), .B(b[67]), .Z(n2382) );
  XNOR U13897 ( .A(n2387), .B(n1648), .Z(n1650) );
  XOR U13898 ( .A(n2388), .B(n2389), .Z(n1648) );
  ANDN U13899 ( .B(n2390), .A(n2391), .Z(n2388) );
  AND U13900 ( .A(a[58]), .B(b[66]), .Z(n2387) );
  XNOR U13901 ( .A(n2392), .B(n1653), .Z(n1655) );
  XOR U13902 ( .A(n2393), .B(n2394), .Z(n1653) );
  ANDN U13903 ( .B(n2395), .A(n2396), .Z(n2393) );
  AND U13904 ( .A(a[59]), .B(b[65]), .Z(n2392) );
  XNOR U13905 ( .A(n2397), .B(n1658), .Z(n1660) );
  XOR U13906 ( .A(n2398), .B(n2399), .Z(n1658) );
  ANDN U13907 ( .B(n2400), .A(n2401), .Z(n2398) );
  AND U13908 ( .A(a[60]), .B(b[64]), .Z(n2397) );
  XNOR U13909 ( .A(n2402), .B(n1663), .Z(n1665) );
  XOR U13910 ( .A(n2403), .B(n2404), .Z(n1663) );
  ANDN U13911 ( .B(n2405), .A(n2406), .Z(n2403) );
  AND U13912 ( .A(a[61]), .B(b[63]), .Z(n2402) );
  XNOR U13913 ( .A(n2407), .B(n1668), .Z(n1670) );
  XOR U13914 ( .A(n2408), .B(n2409), .Z(n1668) );
  ANDN U13915 ( .B(n2410), .A(n2411), .Z(n2408) );
  AND U13916 ( .A(a[62]), .B(b[62]), .Z(n2407) );
  XNOR U13917 ( .A(n2412), .B(n1673), .Z(n1675) );
  XOR U13918 ( .A(n2413), .B(n2414), .Z(n1673) );
  ANDN U13919 ( .B(n2415), .A(n2416), .Z(n2413) );
  AND U13920 ( .A(a[63]), .B(b[61]), .Z(n2412) );
  XNOR U13921 ( .A(n2417), .B(n1678), .Z(n1680) );
  XOR U13922 ( .A(n2418), .B(n2419), .Z(n1678) );
  ANDN U13923 ( .B(n2420), .A(n2421), .Z(n2418) );
  AND U13924 ( .A(a[64]), .B(b[60]), .Z(n2417) );
  XNOR U13925 ( .A(n2422), .B(n1683), .Z(n1685) );
  XOR U13926 ( .A(n2423), .B(n2424), .Z(n1683) );
  ANDN U13927 ( .B(n2425), .A(n2426), .Z(n2423) );
  AND U13928 ( .A(a[65]), .B(b[59]), .Z(n2422) );
  XNOR U13929 ( .A(n2427), .B(n1688), .Z(n1690) );
  XOR U13930 ( .A(n2428), .B(n2429), .Z(n1688) );
  ANDN U13931 ( .B(n2430), .A(n2431), .Z(n2428) );
  AND U13932 ( .A(a[66]), .B(b[58]), .Z(n2427) );
  XNOR U13933 ( .A(n2432), .B(n1693), .Z(n1695) );
  XOR U13934 ( .A(n2433), .B(n2434), .Z(n1693) );
  ANDN U13935 ( .B(n2435), .A(n2436), .Z(n2433) );
  AND U13936 ( .A(a[67]), .B(b[57]), .Z(n2432) );
  XNOR U13937 ( .A(n2437), .B(n1698), .Z(n1700) );
  XOR U13938 ( .A(n2438), .B(n2439), .Z(n1698) );
  ANDN U13939 ( .B(n2440), .A(n2441), .Z(n2438) );
  AND U13940 ( .A(a[68]), .B(b[56]), .Z(n2437) );
  XNOR U13941 ( .A(n2442), .B(n1703), .Z(n1705) );
  XOR U13942 ( .A(n2443), .B(n2444), .Z(n1703) );
  ANDN U13943 ( .B(n2445), .A(n2446), .Z(n2443) );
  AND U13944 ( .A(a[69]), .B(b[55]), .Z(n2442) );
  XNOR U13945 ( .A(n2447), .B(n1708), .Z(n1710) );
  XOR U13946 ( .A(n2448), .B(n2449), .Z(n1708) );
  ANDN U13947 ( .B(n2450), .A(n2451), .Z(n2448) );
  AND U13948 ( .A(a[70]), .B(b[54]), .Z(n2447) );
  XNOR U13949 ( .A(n2452), .B(n1713), .Z(n1715) );
  XOR U13950 ( .A(n2453), .B(n2454), .Z(n1713) );
  ANDN U13951 ( .B(n2455), .A(n2456), .Z(n2453) );
  AND U13952 ( .A(a[71]), .B(b[53]), .Z(n2452) );
  XNOR U13953 ( .A(n2457), .B(n1718), .Z(n1720) );
  XOR U13954 ( .A(n2458), .B(n2459), .Z(n1718) );
  ANDN U13955 ( .B(n2460), .A(n2461), .Z(n2458) );
  AND U13956 ( .A(a[72]), .B(b[52]), .Z(n2457) );
  XNOR U13957 ( .A(n2462), .B(n1723), .Z(n1725) );
  XOR U13958 ( .A(n2463), .B(n2464), .Z(n1723) );
  ANDN U13959 ( .B(n2465), .A(n2466), .Z(n2463) );
  AND U13960 ( .A(a[73]), .B(b[51]), .Z(n2462) );
  XNOR U13961 ( .A(n2467), .B(n1728), .Z(n1730) );
  XOR U13962 ( .A(n2468), .B(n2469), .Z(n1728) );
  ANDN U13963 ( .B(n2470), .A(n2471), .Z(n2468) );
  AND U13964 ( .A(a[74]), .B(b[50]), .Z(n2467) );
  XNOR U13965 ( .A(n2472), .B(n1733), .Z(n1735) );
  XOR U13966 ( .A(n2473), .B(n2474), .Z(n1733) );
  ANDN U13967 ( .B(n2475), .A(n2476), .Z(n2473) );
  AND U13968 ( .A(a[75]), .B(b[49]), .Z(n2472) );
  XNOR U13969 ( .A(n2477), .B(n1738), .Z(n1740) );
  XOR U13970 ( .A(n2478), .B(n2479), .Z(n1738) );
  ANDN U13971 ( .B(n2480), .A(n2481), .Z(n2478) );
  AND U13972 ( .A(a[76]), .B(b[48]), .Z(n2477) );
  XNOR U13973 ( .A(n2482), .B(n1743), .Z(n1745) );
  XOR U13974 ( .A(n2483), .B(n2484), .Z(n1743) );
  ANDN U13975 ( .B(n2485), .A(n2486), .Z(n2483) );
  AND U13976 ( .A(a[77]), .B(b[47]), .Z(n2482) );
  XNOR U13977 ( .A(n2487), .B(n1748), .Z(n1750) );
  XOR U13978 ( .A(n2488), .B(n2489), .Z(n1748) );
  ANDN U13979 ( .B(n2490), .A(n2491), .Z(n2488) );
  AND U13980 ( .A(a[78]), .B(b[46]), .Z(n2487) );
  XNOR U13981 ( .A(n2492), .B(n1753), .Z(n1755) );
  XOR U13982 ( .A(n2493), .B(n2494), .Z(n1753) );
  ANDN U13983 ( .B(n2495), .A(n2496), .Z(n2493) );
  AND U13984 ( .A(a[79]), .B(b[45]), .Z(n2492) );
  XNOR U13985 ( .A(n2497), .B(n1758), .Z(n1760) );
  XOR U13986 ( .A(n2498), .B(n2499), .Z(n1758) );
  ANDN U13987 ( .B(n2500), .A(n2501), .Z(n2498) );
  AND U13988 ( .A(a[80]), .B(b[44]), .Z(n2497) );
  XNOR U13989 ( .A(n2502), .B(n1763), .Z(n1765) );
  XOR U13990 ( .A(n2503), .B(n2504), .Z(n1763) );
  ANDN U13991 ( .B(n2505), .A(n2506), .Z(n2503) );
  AND U13992 ( .A(a[81]), .B(b[43]), .Z(n2502) );
  XNOR U13993 ( .A(n2507), .B(n1768), .Z(n1770) );
  XOR U13994 ( .A(n2508), .B(n2509), .Z(n1768) );
  ANDN U13995 ( .B(n2510), .A(n2511), .Z(n2508) );
  AND U13996 ( .A(a[82]), .B(b[42]), .Z(n2507) );
  XNOR U13997 ( .A(n2512), .B(n1773), .Z(n1775) );
  XOR U13998 ( .A(n2513), .B(n2514), .Z(n1773) );
  ANDN U13999 ( .B(n2515), .A(n2516), .Z(n2513) );
  AND U14000 ( .A(a[83]), .B(b[41]), .Z(n2512) );
  XNOR U14001 ( .A(n2517), .B(n1778), .Z(n1780) );
  XOR U14002 ( .A(n2518), .B(n2519), .Z(n1778) );
  ANDN U14003 ( .B(n2520), .A(n2521), .Z(n2518) );
  AND U14004 ( .A(a[84]), .B(b[40]), .Z(n2517) );
  XNOR U14005 ( .A(n2522), .B(n1783), .Z(n1785) );
  XOR U14006 ( .A(n2523), .B(n2524), .Z(n1783) );
  ANDN U14007 ( .B(n2525), .A(n2526), .Z(n2523) );
  AND U14008 ( .A(a[85]), .B(b[39]), .Z(n2522) );
  XNOR U14009 ( .A(n2527), .B(n1788), .Z(n1790) );
  XOR U14010 ( .A(n2528), .B(n2529), .Z(n1788) );
  ANDN U14011 ( .B(n2530), .A(n2531), .Z(n2528) );
  AND U14012 ( .A(a[86]), .B(b[38]), .Z(n2527) );
  XNOR U14013 ( .A(n2532), .B(n1793), .Z(n1795) );
  XOR U14014 ( .A(n2533), .B(n2534), .Z(n1793) );
  ANDN U14015 ( .B(n2535), .A(n2536), .Z(n2533) );
  AND U14016 ( .A(a[87]), .B(b[37]), .Z(n2532) );
  XNOR U14017 ( .A(n2537), .B(n1798), .Z(n1800) );
  XOR U14018 ( .A(n2538), .B(n2539), .Z(n1798) );
  ANDN U14019 ( .B(n2540), .A(n2541), .Z(n2538) );
  AND U14020 ( .A(a[88]), .B(b[36]), .Z(n2537) );
  XNOR U14021 ( .A(n2542), .B(n1803), .Z(n1805) );
  XOR U14022 ( .A(n2543), .B(n2544), .Z(n1803) );
  ANDN U14023 ( .B(n2545), .A(n2546), .Z(n2543) );
  AND U14024 ( .A(a[89]), .B(b[35]), .Z(n2542) );
  XNOR U14025 ( .A(n2547), .B(n1808), .Z(n1810) );
  XOR U14026 ( .A(n2548), .B(n2549), .Z(n1808) );
  ANDN U14027 ( .B(n2550), .A(n2551), .Z(n2548) );
  AND U14028 ( .A(a[90]), .B(b[34]), .Z(n2547) );
  XNOR U14029 ( .A(n2552), .B(n1813), .Z(n1815) );
  XOR U14030 ( .A(n2553), .B(n2554), .Z(n1813) );
  ANDN U14031 ( .B(n2555), .A(n2556), .Z(n2553) );
  AND U14032 ( .A(a[91]), .B(b[33]), .Z(n2552) );
  XNOR U14033 ( .A(n2557), .B(n1818), .Z(n1820) );
  XOR U14034 ( .A(n2558), .B(n2559), .Z(n1818) );
  ANDN U14035 ( .B(n2560), .A(n2561), .Z(n2558) );
  AND U14036 ( .A(a[92]), .B(b[32]), .Z(n2557) );
  XNOR U14037 ( .A(n2562), .B(n1823), .Z(n1825) );
  XOR U14038 ( .A(n2563), .B(n2564), .Z(n1823) );
  ANDN U14039 ( .B(n2565), .A(n2566), .Z(n2563) );
  AND U14040 ( .A(a[93]), .B(b[31]), .Z(n2562) );
  XNOR U14041 ( .A(n2567), .B(n1828), .Z(n1830) );
  XOR U14042 ( .A(n2568), .B(n2569), .Z(n1828) );
  ANDN U14043 ( .B(n2570), .A(n2571), .Z(n2568) );
  AND U14044 ( .A(a[94]), .B(b[30]), .Z(n2567) );
  XNOR U14045 ( .A(n2572), .B(n1833), .Z(n1835) );
  XOR U14046 ( .A(n2573), .B(n2574), .Z(n1833) );
  ANDN U14047 ( .B(n2575), .A(n2576), .Z(n2573) );
  AND U14048 ( .A(a[95]), .B(b[29]), .Z(n2572) );
  XNOR U14049 ( .A(n2577), .B(n1838), .Z(n1840) );
  XOR U14050 ( .A(n2578), .B(n2579), .Z(n1838) );
  ANDN U14051 ( .B(n2580), .A(n2581), .Z(n2578) );
  AND U14052 ( .A(a[96]), .B(b[28]), .Z(n2577) );
  XNOR U14053 ( .A(n2582), .B(n1843), .Z(n1845) );
  XOR U14054 ( .A(n2583), .B(n2584), .Z(n1843) );
  ANDN U14055 ( .B(n2585), .A(n2586), .Z(n2583) );
  AND U14056 ( .A(a[97]), .B(b[27]), .Z(n2582) );
  XNOR U14057 ( .A(n2587), .B(n1848), .Z(n1850) );
  XOR U14058 ( .A(n2588), .B(n2589), .Z(n1848) );
  ANDN U14059 ( .B(n2590), .A(n2591), .Z(n2588) );
  AND U14060 ( .A(a[98]), .B(b[26]), .Z(n2587) );
  XNOR U14061 ( .A(n2592), .B(n1853), .Z(n1855) );
  XOR U14062 ( .A(n2593), .B(n2594), .Z(n1853) );
  ANDN U14063 ( .B(n2595), .A(n2596), .Z(n2593) );
  AND U14064 ( .A(a[99]), .B(b[25]), .Z(n2592) );
  XNOR U14065 ( .A(n2597), .B(n1858), .Z(n1860) );
  XOR U14066 ( .A(n2598), .B(n2599), .Z(n1858) );
  ANDN U14067 ( .B(n2600), .A(n2601), .Z(n2598) );
  AND U14068 ( .A(b[24]), .B(a[100]), .Z(n2597) );
  XNOR U14069 ( .A(n2602), .B(n1863), .Z(n1865) );
  XOR U14070 ( .A(n2603), .B(n2604), .Z(n1863) );
  ANDN U14071 ( .B(n2605), .A(n2606), .Z(n2603) );
  AND U14072 ( .A(b[23]), .B(a[101]), .Z(n2602) );
  XNOR U14073 ( .A(n2607), .B(n1868), .Z(n1870) );
  XOR U14074 ( .A(n2608), .B(n2609), .Z(n1868) );
  ANDN U14075 ( .B(n2610), .A(n2611), .Z(n2608) );
  AND U14076 ( .A(b[22]), .B(a[102]), .Z(n2607) );
  XNOR U14077 ( .A(n2612), .B(n1873), .Z(n1875) );
  XOR U14078 ( .A(n2613), .B(n2614), .Z(n1873) );
  ANDN U14079 ( .B(n2615), .A(n2616), .Z(n2613) );
  AND U14080 ( .A(b[21]), .B(a[103]), .Z(n2612) );
  XNOR U14081 ( .A(n2617), .B(n1878), .Z(n1880) );
  XOR U14082 ( .A(n2618), .B(n2619), .Z(n1878) );
  ANDN U14083 ( .B(n2620), .A(n2621), .Z(n2618) );
  AND U14084 ( .A(b[20]), .B(a[104]), .Z(n2617) );
  XNOR U14085 ( .A(n2622), .B(n1883), .Z(n1885) );
  XOR U14086 ( .A(n2623), .B(n2624), .Z(n1883) );
  ANDN U14087 ( .B(n2625), .A(n2626), .Z(n2623) );
  AND U14088 ( .A(b[19]), .B(a[105]), .Z(n2622) );
  XNOR U14089 ( .A(n2627), .B(n1888), .Z(n1890) );
  XOR U14090 ( .A(n2628), .B(n2629), .Z(n1888) );
  ANDN U14091 ( .B(n2630), .A(n2631), .Z(n2628) );
  AND U14092 ( .A(b[18]), .B(a[106]), .Z(n2627) );
  XNOR U14093 ( .A(n2632), .B(n1893), .Z(n1895) );
  XOR U14094 ( .A(n2633), .B(n2634), .Z(n1893) );
  ANDN U14095 ( .B(n2635), .A(n2636), .Z(n2633) );
  AND U14096 ( .A(b[17]), .B(a[107]), .Z(n2632) );
  XNOR U14097 ( .A(n2637), .B(n1898), .Z(n1900) );
  XOR U14098 ( .A(n2638), .B(n2639), .Z(n1898) );
  ANDN U14099 ( .B(n2640), .A(n2641), .Z(n2638) );
  AND U14100 ( .A(b[16]), .B(a[108]), .Z(n2637) );
  XNOR U14101 ( .A(n2642), .B(n1903), .Z(n1905) );
  XOR U14102 ( .A(n2643), .B(n2644), .Z(n1903) );
  ANDN U14103 ( .B(n2645), .A(n2646), .Z(n2643) );
  AND U14104 ( .A(b[15]), .B(a[109]), .Z(n2642) );
  XNOR U14105 ( .A(n2647), .B(n1908), .Z(n1910) );
  XOR U14106 ( .A(n2648), .B(n2649), .Z(n1908) );
  ANDN U14107 ( .B(n2650), .A(n2651), .Z(n2648) );
  AND U14108 ( .A(b[14]), .B(a[110]), .Z(n2647) );
  XNOR U14109 ( .A(n2652), .B(n1913), .Z(n1915) );
  XOR U14110 ( .A(n2653), .B(n2654), .Z(n1913) );
  ANDN U14111 ( .B(n2655), .A(n2656), .Z(n2653) );
  AND U14112 ( .A(b[13]), .B(a[111]), .Z(n2652) );
  XNOR U14113 ( .A(n2657), .B(n1918), .Z(n1920) );
  XOR U14114 ( .A(n2658), .B(n2659), .Z(n1918) );
  ANDN U14115 ( .B(n2660), .A(n2661), .Z(n2658) );
  AND U14116 ( .A(b[12]), .B(a[112]), .Z(n2657) );
  XNOR U14117 ( .A(n2662), .B(n1923), .Z(n1925) );
  XOR U14118 ( .A(n2663), .B(n2664), .Z(n1923) );
  ANDN U14119 ( .B(n2665), .A(n2666), .Z(n2663) );
  AND U14120 ( .A(b[11]), .B(a[113]), .Z(n2662) );
  XNOR U14121 ( .A(n2667), .B(n1928), .Z(n1930) );
  XOR U14122 ( .A(n2668), .B(n2669), .Z(n1928) );
  ANDN U14123 ( .B(n2670), .A(n2671), .Z(n2668) );
  AND U14124 ( .A(b[10]), .B(a[114]), .Z(n2667) );
  XNOR U14125 ( .A(n2672), .B(n1933), .Z(n1935) );
  XOR U14126 ( .A(n2673), .B(n2674), .Z(n1933) );
  ANDN U14127 ( .B(n2675), .A(n2676), .Z(n2673) );
  AND U14128 ( .A(b[9]), .B(a[115]), .Z(n2672) );
  XNOR U14129 ( .A(n2677), .B(n1938), .Z(n1940) );
  XOR U14130 ( .A(n2678), .B(n2679), .Z(n1938) );
  ANDN U14131 ( .B(n2680), .A(n2681), .Z(n2678) );
  AND U14132 ( .A(b[8]), .B(a[116]), .Z(n2677) );
  XNOR U14133 ( .A(n2682), .B(n1943), .Z(n1945) );
  XOR U14134 ( .A(n2683), .B(n2684), .Z(n1943) );
  ANDN U14135 ( .B(n2685), .A(n2686), .Z(n2683) );
  AND U14136 ( .A(b[7]), .B(a[117]), .Z(n2682) );
  XNOR U14137 ( .A(n2687), .B(n1948), .Z(n1950) );
  XOR U14138 ( .A(n2688), .B(n2689), .Z(n1948) );
  ANDN U14139 ( .B(n2690), .A(n2691), .Z(n2688) );
  AND U14140 ( .A(b[6]), .B(a[118]), .Z(n2687) );
  XNOR U14141 ( .A(n2692), .B(n1953), .Z(n1955) );
  XOR U14142 ( .A(n2693), .B(n2694), .Z(n1953) );
  ANDN U14143 ( .B(n2695), .A(n2696), .Z(n2693) );
  AND U14144 ( .A(b[5]), .B(a[119]), .Z(n2692) );
  XNOR U14145 ( .A(n2697), .B(n1958), .Z(n1960) );
  XOR U14146 ( .A(n2698), .B(n2699), .Z(n1958) );
  ANDN U14147 ( .B(n2700), .A(n2701), .Z(n2698) );
  AND U14148 ( .A(b[4]), .B(a[120]), .Z(n2697) );
  XNOR U14149 ( .A(n2702), .B(n2703), .Z(n1972) );
  NANDN U14150 ( .A(n2704), .B(n2705), .Z(n2703) );
  XNOR U14151 ( .A(n2706), .B(n1963), .Z(n1965) );
  XNOR U14152 ( .A(n2707), .B(n2708), .Z(n1963) );
  AND U14153 ( .A(n2709), .B(n2710), .Z(n2707) );
  AND U14154 ( .A(b[3]), .B(a[121]), .Z(n2706) );
  NAND U14155 ( .A(a[124]), .B(b[0]), .Z(n982) );
  XNOR U14156 ( .A(n1978), .B(n1979), .Z(c[123]) );
  XNOR U14157 ( .A(n2704), .B(n2705), .Z(n1979) );
  XOR U14158 ( .A(n2702), .B(n2711), .Z(n2705) );
  NAND U14159 ( .A(b[1]), .B(a[122]), .Z(n2711) );
  XOR U14160 ( .A(n2710), .B(n2712), .Z(n2704) );
  XOR U14161 ( .A(n2702), .B(n2709), .Z(n2712) );
  XNOR U14162 ( .A(n2713), .B(n2708), .Z(n2709) );
  AND U14163 ( .A(b[2]), .B(a[121]), .Z(n2713) );
  NANDN U14164 ( .A(n2714), .B(n2715), .Z(n2702) );
  XOR U14165 ( .A(n2708), .B(n2700), .Z(n2716) );
  XNOR U14166 ( .A(n2699), .B(n2695), .Z(n2717) );
  XNOR U14167 ( .A(n2694), .B(n2690), .Z(n2718) );
  XNOR U14168 ( .A(n2689), .B(n2685), .Z(n2719) );
  XNOR U14169 ( .A(n2684), .B(n2680), .Z(n2720) );
  XNOR U14170 ( .A(n2679), .B(n2675), .Z(n2721) );
  XNOR U14171 ( .A(n2674), .B(n2670), .Z(n2722) );
  XNOR U14172 ( .A(n2669), .B(n2665), .Z(n2723) );
  XNOR U14173 ( .A(n2664), .B(n2660), .Z(n2724) );
  XNOR U14174 ( .A(n2659), .B(n2655), .Z(n2725) );
  XNOR U14175 ( .A(n2654), .B(n2650), .Z(n2726) );
  XNOR U14176 ( .A(n2649), .B(n2645), .Z(n2727) );
  XNOR U14177 ( .A(n2644), .B(n2640), .Z(n2728) );
  XNOR U14178 ( .A(n2639), .B(n2635), .Z(n2729) );
  XNOR U14179 ( .A(n2634), .B(n2630), .Z(n2730) );
  XNOR U14180 ( .A(n2629), .B(n2625), .Z(n2731) );
  XNOR U14181 ( .A(n2624), .B(n2620), .Z(n2732) );
  XNOR U14182 ( .A(n2619), .B(n2615), .Z(n2733) );
  XNOR U14183 ( .A(n2614), .B(n2610), .Z(n2734) );
  XNOR U14184 ( .A(n2609), .B(n2605), .Z(n2735) );
  XNOR U14185 ( .A(n2604), .B(n2600), .Z(n2736) );
  XNOR U14186 ( .A(n2599), .B(n2595), .Z(n2737) );
  XNOR U14187 ( .A(n2594), .B(n2590), .Z(n2738) );
  XNOR U14188 ( .A(n2589), .B(n2585), .Z(n2739) );
  XNOR U14189 ( .A(n2584), .B(n2580), .Z(n2740) );
  XNOR U14190 ( .A(n2579), .B(n2575), .Z(n2741) );
  XNOR U14191 ( .A(n2574), .B(n2570), .Z(n2742) );
  XNOR U14192 ( .A(n2569), .B(n2565), .Z(n2743) );
  XNOR U14193 ( .A(n2564), .B(n2560), .Z(n2744) );
  XNOR U14194 ( .A(n2559), .B(n2555), .Z(n2745) );
  XNOR U14195 ( .A(n2554), .B(n2550), .Z(n2746) );
  XNOR U14196 ( .A(n2549), .B(n2545), .Z(n2747) );
  XNOR U14197 ( .A(n2544), .B(n2540), .Z(n2748) );
  XNOR U14198 ( .A(n2539), .B(n2535), .Z(n2749) );
  XNOR U14199 ( .A(n2534), .B(n2530), .Z(n2750) );
  XNOR U14200 ( .A(n2529), .B(n2525), .Z(n2751) );
  XNOR U14201 ( .A(n2524), .B(n2520), .Z(n2752) );
  XNOR U14202 ( .A(n2519), .B(n2515), .Z(n2753) );
  XNOR U14203 ( .A(n2514), .B(n2510), .Z(n2754) );
  XNOR U14204 ( .A(n2509), .B(n2505), .Z(n2755) );
  XNOR U14205 ( .A(n2504), .B(n2500), .Z(n2756) );
  XNOR U14206 ( .A(n2499), .B(n2495), .Z(n2757) );
  XNOR U14207 ( .A(n2494), .B(n2490), .Z(n2758) );
  XNOR U14208 ( .A(n2489), .B(n2485), .Z(n2759) );
  XNOR U14209 ( .A(n2484), .B(n2480), .Z(n2760) );
  XNOR U14210 ( .A(n2479), .B(n2475), .Z(n2761) );
  XNOR U14211 ( .A(n2474), .B(n2470), .Z(n2762) );
  XNOR U14212 ( .A(n2469), .B(n2465), .Z(n2763) );
  XNOR U14213 ( .A(n2464), .B(n2460), .Z(n2764) );
  XNOR U14214 ( .A(n2459), .B(n2455), .Z(n2765) );
  XNOR U14215 ( .A(n2454), .B(n2450), .Z(n2766) );
  XNOR U14216 ( .A(n2449), .B(n2445), .Z(n2767) );
  XNOR U14217 ( .A(n2444), .B(n2440), .Z(n2768) );
  XNOR U14218 ( .A(n2439), .B(n2435), .Z(n2769) );
  XNOR U14219 ( .A(n2434), .B(n2430), .Z(n2770) );
  XNOR U14220 ( .A(n2429), .B(n2425), .Z(n2771) );
  XNOR U14221 ( .A(n2424), .B(n2420), .Z(n2772) );
  XNOR U14222 ( .A(n2419), .B(n2415), .Z(n2773) );
  XNOR U14223 ( .A(n2414), .B(n2410), .Z(n2774) );
  XNOR U14224 ( .A(n2409), .B(n2405), .Z(n2775) );
  XNOR U14225 ( .A(n2404), .B(n2400), .Z(n2776) );
  XNOR U14226 ( .A(n2399), .B(n2395), .Z(n2777) );
  XNOR U14227 ( .A(n2394), .B(n2390), .Z(n2778) );
  XNOR U14228 ( .A(n2389), .B(n2385), .Z(n2779) );
  XNOR U14229 ( .A(n2384), .B(n2380), .Z(n2780) );
  XNOR U14230 ( .A(n2379), .B(n2375), .Z(n2781) );
  XNOR U14231 ( .A(n2374), .B(n2370), .Z(n2782) );
  XNOR U14232 ( .A(n2369), .B(n2365), .Z(n2783) );
  XNOR U14233 ( .A(n2364), .B(n2360), .Z(n2784) );
  XNOR U14234 ( .A(n2359), .B(n2355), .Z(n2785) );
  XNOR U14235 ( .A(n2354), .B(n2350), .Z(n2786) );
  XNOR U14236 ( .A(n2349), .B(n2345), .Z(n2787) );
  XNOR U14237 ( .A(n2344), .B(n2340), .Z(n2788) );
  XNOR U14238 ( .A(n2339), .B(n2335), .Z(n2789) );
  XNOR U14239 ( .A(n2334), .B(n2330), .Z(n2790) );
  XNOR U14240 ( .A(n2329), .B(n2325), .Z(n2791) );
  XNOR U14241 ( .A(n2324), .B(n2320), .Z(n2792) );
  XNOR U14242 ( .A(n2319), .B(n2315), .Z(n2793) );
  XNOR U14243 ( .A(n2314), .B(n2310), .Z(n2794) );
  XNOR U14244 ( .A(n2309), .B(n2305), .Z(n2795) );
  XNOR U14245 ( .A(n2304), .B(n2300), .Z(n2796) );
  XNOR U14246 ( .A(n2299), .B(n2295), .Z(n2797) );
  XNOR U14247 ( .A(n2294), .B(n2290), .Z(n2798) );
  XNOR U14248 ( .A(n2289), .B(n2285), .Z(n2799) );
  XNOR U14249 ( .A(n2284), .B(n2280), .Z(n2800) );
  XNOR U14250 ( .A(n2279), .B(n2275), .Z(n2801) );
  XNOR U14251 ( .A(n2274), .B(n2270), .Z(n2802) );
  XNOR U14252 ( .A(n2269), .B(n2265), .Z(n2803) );
  XNOR U14253 ( .A(n2264), .B(n2260), .Z(n2804) );
  XNOR U14254 ( .A(n2259), .B(n2255), .Z(n2805) );
  XNOR U14255 ( .A(n2254), .B(n2250), .Z(n2806) );
  XNOR U14256 ( .A(n2249), .B(n2245), .Z(n2807) );
  XNOR U14257 ( .A(n2244), .B(n2240), .Z(n2808) );
  XNOR U14258 ( .A(n2239), .B(n2235), .Z(n2809) );
  XNOR U14259 ( .A(n2234), .B(n2230), .Z(n2810) );
  XNOR U14260 ( .A(n2229), .B(n2225), .Z(n2811) );
  XNOR U14261 ( .A(n2224), .B(n2220), .Z(n2812) );
  XNOR U14262 ( .A(n2219), .B(n2215), .Z(n2813) );
  XNOR U14263 ( .A(n2214), .B(n2210), .Z(n2814) );
  XNOR U14264 ( .A(n2209), .B(n2205), .Z(n2815) );
  XNOR U14265 ( .A(n2204), .B(n2200), .Z(n2816) );
  XNOR U14266 ( .A(n2199), .B(n2195), .Z(n2817) );
  XNOR U14267 ( .A(n2194), .B(n2190), .Z(n2818) );
  XNOR U14268 ( .A(n2189), .B(n2185), .Z(n2819) );
  XNOR U14269 ( .A(n2184), .B(n2180), .Z(n2820) );
  XNOR U14270 ( .A(n2179), .B(n2175), .Z(n2821) );
  XNOR U14271 ( .A(n2174), .B(n2170), .Z(n2822) );
  XNOR U14272 ( .A(n2169), .B(n2165), .Z(n2823) );
  XNOR U14273 ( .A(n2164), .B(n2160), .Z(n2824) );
  XNOR U14274 ( .A(n2159), .B(n2155), .Z(n2825) );
  XNOR U14275 ( .A(n2154), .B(n2150), .Z(n2826) );
  XNOR U14276 ( .A(n2149), .B(n2145), .Z(n2827) );
  XNOR U14277 ( .A(n2144), .B(n2140), .Z(n2828) );
  XNOR U14278 ( .A(n2139), .B(n2135), .Z(n2829) );
  XNOR U14279 ( .A(n2134), .B(n2130), .Z(n2830) );
  XNOR U14280 ( .A(n2129), .B(n2125), .Z(n2831) );
  XNOR U14281 ( .A(n2124), .B(n2120), .Z(n2832) );
  XNOR U14282 ( .A(n2119), .B(n2115), .Z(n2833) );
  XNOR U14283 ( .A(n2114), .B(n2110), .Z(n2834) );
  XNOR U14284 ( .A(n2109), .B(n2105), .Z(n2835) );
  XNOR U14285 ( .A(n2836), .B(n2104), .Z(n2105) );
  AND U14286 ( .A(a[0]), .B(b[123]), .Z(n2836) );
  XOR U14287 ( .A(n2837), .B(n2104), .Z(n2106) );
  XNOR U14288 ( .A(n2838), .B(n2839), .Z(n2104) );
  ANDN U14289 ( .B(n2840), .A(n2841), .Z(n2838) );
  AND U14290 ( .A(a[1]), .B(b[122]), .Z(n2837) );
  XNOR U14291 ( .A(n2842), .B(n2109), .Z(n2111) );
  XOR U14292 ( .A(n2843), .B(n2844), .Z(n2109) );
  ANDN U14293 ( .B(n2845), .A(n2846), .Z(n2843) );
  AND U14294 ( .A(a[2]), .B(b[121]), .Z(n2842) );
  XNOR U14295 ( .A(n2847), .B(n2114), .Z(n2116) );
  XOR U14296 ( .A(n2848), .B(n2849), .Z(n2114) );
  ANDN U14297 ( .B(n2850), .A(n2851), .Z(n2848) );
  AND U14298 ( .A(a[3]), .B(b[120]), .Z(n2847) );
  XNOR U14299 ( .A(n2852), .B(n2119), .Z(n2121) );
  XOR U14300 ( .A(n2853), .B(n2854), .Z(n2119) );
  ANDN U14301 ( .B(n2855), .A(n2856), .Z(n2853) );
  AND U14302 ( .A(a[4]), .B(b[119]), .Z(n2852) );
  XNOR U14303 ( .A(n2857), .B(n2124), .Z(n2126) );
  XOR U14304 ( .A(n2858), .B(n2859), .Z(n2124) );
  ANDN U14305 ( .B(n2860), .A(n2861), .Z(n2858) );
  AND U14306 ( .A(a[5]), .B(b[118]), .Z(n2857) );
  XNOR U14307 ( .A(n2862), .B(n2129), .Z(n2131) );
  XOR U14308 ( .A(n2863), .B(n2864), .Z(n2129) );
  ANDN U14309 ( .B(n2865), .A(n2866), .Z(n2863) );
  AND U14310 ( .A(a[6]), .B(b[117]), .Z(n2862) );
  XNOR U14311 ( .A(n2867), .B(n2134), .Z(n2136) );
  XOR U14312 ( .A(n2868), .B(n2869), .Z(n2134) );
  ANDN U14313 ( .B(n2870), .A(n2871), .Z(n2868) );
  AND U14314 ( .A(a[7]), .B(b[116]), .Z(n2867) );
  XNOR U14315 ( .A(n2872), .B(n2139), .Z(n2141) );
  XOR U14316 ( .A(n2873), .B(n2874), .Z(n2139) );
  ANDN U14317 ( .B(n2875), .A(n2876), .Z(n2873) );
  AND U14318 ( .A(a[8]), .B(b[115]), .Z(n2872) );
  XNOR U14319 ( .A(n2877), .B(n2144), .Z(n2146) );
  XOR U14320 ( .A(n2878), .B(n2879), .Z(n2144) );
  ANDN U14321 ( .B(n2880), .A(n2881), .Z(n2878) );
  AND U14322 ( .A(a[9]), .B(b[114]), .Z(n2877) );
  XNOR U14323 ( .A(n2882), .B(n2149), .Z(n2151) );
  XOR U14324 ( .A(n2883), .B(n2884), .Z(n2149) );
  ANDN U14325 ( .B(n2885), .A(n2886), .Z(n2883) );
  AND U14326 ( .A(a[10]), .B(b[113]), .Z(n2882) );
  XNOR U14327 ( .A(n2887), .B(n2154), .Z(n2156) );
  XOR U14328 ( .A(n2888), .B(n2889), .Z(n2154) );
  ANDN U14329 ( .B(n2890), .A(n2891), .Z(n2888) );
  AND U14330 ( .A(a[11]), .B(b[112]), .Z(n2887) );
  XNOR U14331 ( .A(n2892), .B(n2159), .Z(n2161) );
  XOR U14332 ( .A(n2893), .B(n2894), .Z(n2159) );
  ANDN U14333 ( .B(n2895), .A(n2896), .Z(n2893) );
  AND U14334 ( .A(a[12]), .B(b[111]), .Z(n2892) );
  XNOR U14335 ( .A(n2897), .B(n2164), .Z(n2166) );
  XOR U14336 ( .A(n2898), .B(n2899), .Z(n2164) );
  ANDN U14337 ( .B(n2900), .A(n2901), .Z(n2898) );
  AND U14338 ( .A(a[13]), .B(b[110]), .Z(n2897) );
  XNOR U14339 ( .A(n2902), .B(n2169), .Z(n2171) );
  XOR U14340 ( .A(n2903), .B(n2904), .Z(n2169) );
  ANDN U14341 ( .B(n2905), .A(n2906), .Z(n2903) );
  AND U14342 ( .A(a[14]), .B(b[109]), .Z(n2902) );
  XNOR U14343 ( .A(n2907), .B(n2174), .Z(n2176) );
  XOR U14344 ( .A(n2908), .B(n2909), .Z(n2174) );
  ANDN U14345 ( .B(n2910), .A(n2911), .Z(n2908) );
  AND U14346 ( .A(a[15]), .B(b[108]), .Z(n2907) );
  XNOR U14347 ( .A(n2912), .B(n2179), .Z(n2181) );
  XOR U14348 ( .A(n2913), .B(n2914), .Z(n2179) );
  ANDN U14349 ( .B(n2915), .A(n2916), .Z(n2913) );
  AND U14350 ( .A(a[16]), .B(b[107]), .Z(n2912) );
  XNOR U14351 ( .A(n2917), .B(n2184), .Z(n2186) );
  XOR U14352 ( .A(n2918), .B(n2919), .Z(n2184) );
  ANDN U14353 ( .B(n2920), .A(n2921), .Z(n2918) );
  AND U14354 ( .A(a[17]), .B(b[106]), .Z(n2917) );
  XNOR U14355 ( .A(n2922), .B(n2189), .Z(n2191) );
  XOR U14356 ( .A(n2923), .B(n2924), .Z(n2189) );
  ANDN U14357 ( .B(n2925), .A(n2926), .Z(n2923) );
  AND U14358 ( .A(a[18]), .B(b[105]), .Z(n2922) );
  XNOR U14359 ( .A(n2927), .B(n2194), .Z(n2196) );
  XOR U14360 ( .A(n2928), .B(n2929), .Z(n2194) );
  ANDN U14361 ( .B(n2930), .A(n2931), .Z(n2928) );
  AND U14362 ( .A(a[19]), .B(b[104]), .Z(n2927) );
  XNOR U14363 ( .A(n2932), .B(n2199), .Z(n2201) );
  XOR U14364 ( .A(n2933), .B(n2934), .Z(n2199) );
  ANDN U14365 ( .B(n2935), .A(n2936), .Z(n2933) );
  AND U14366 ( .A(a[20]), .B(b[103]), .Z(n2932) );
  XNOR U14367 ( .A(n2937), .B(n2204), .Z(n2206) );
  XOR U14368 ( .A(n2938), .B(n2939), .Z(n2204) );
  ANDN U14369 ( .B(n2940), .A(n2941), .Z(n2938) );
  AND U14370 ( .A(a[21]), .B(b[102]), .Z(n2937) );
  XNOR U14371 ( .A(n2942), .B(n2209), .Z(n2211) );
  XOR U14372 ( .A(n2943), .B(n2944), .Z(n2209) );
  ANDN U14373 ( .B(n2945), .A(n2946), .Z(n2943) );
  AND U14374 ( .A(a[22]), .B(b[101]), .Z(n2942) );
  XNOR U14375 ( .A(n2947), .B(n2214), .Z(n2216) );
  XOR U14376 ( .A(n2948), .B(n2949), .Z(n2214) );
  ANDN U14377 ( .B(n2950), .A(n2951), .Z(n2948) );
  AND U14378 ( .A(a[23]), .B(b[100]), .Z(n2947) );
  XNOR U14379 ( .A(n2952), .B(n2219), .Z(n2221) );
  XOR U14380 ( .A(n2953), .B(n2954), .Z(n2219) );
  ANDN U14381 ( .B(n2955), .A(n2956), .Z(n2953) );
  AND U14382 ( .A(a[24]), .B(b[99]), .Z(n2952) );
  XNOR U14383 ( .A(n2957), .B(n2224), .Z(n2226) );
  XOR U14384 ( .A(n2958), .B(n2959), .Z(n2224) );
  ANDN U14385 ( .B(n2960), .A(n2961), .Z(n2958) );
  AND U14386 ( .A(a[25]), .B(b[98]), .Z(n2957) );
  XNOR U14387 ( .A(n2962), .B(n2229), .Z(n2231) );
  XOR U14388 ( .A(n2963), .B(n2964), .Z(n2229) );
  ANDN U14389 ( .B(n2965), .A(n2966), .Z(n2963) );
  AND U14390 ( .A(a[26]), .B(b[97]), .Z(n2962) );
  XNOR U14391 ( .A(n2967), .B(n2234), .Z(n2236) );
  XOR U14392 ( .A(n2968), .B(n2969), .Z(n2234) );
  ANDN U14393 ( .B(n2970), .A(n2971), .Z(n2968) );
  AND U14394 ( .A(a[27]), .B(b[96]), .Z(n2967) );
  XNOR U14395 ( .A(n2972), .B(n2239), .Z(n2241) );
  XOR U14396 ( .A(n2973), .B(n2974), .Z(n2239) );
  ANDN U14397 ( .B(n2975), .A(n2976), .Z(n2973) );
  AND U14398 ( .A(a[28]), .B(b[95]), .Z(n2972) );
  XNOR U14399 ( .A(n2977), .B(n2244), .Z(n2246) );
  XOR U14400 ( .A(n2978), .B(n2979), .Z(n2244) );
  ANDN U14401 ( .B(n2980), .A(n2981), .Z(n2978) );
  AND U14402 ( .A(a[29]), .B(b[94]), .Z(n2977) );
  XNOR U14403 ( .A(n2982), .B(n2249), .Z(n2251) );
  XOR U14404 ( .A(n2983), .B(n2984), .Z(n2249) );
  ANDN U14405 ( .B(n2985), .A(n2986), .Z(n2983) );
  AND U14406 ( .A(a[30]), .B(b[93]), .Z(n2982) );
  XNOR U14407 ( .A(n2987), .B(n2254), .Z(n2256) );
  XOR U14408 ( .A(n2988), .B(n2989), .Z(n2254) );
  ANDN U14409 ( .B(n2990), .A(n2991), .Z(n2988) );
  AND U14410 ( .A(a[31]), .B(b[92]), .Z(n2987) );
  XNOR U14411 ( .A(n2992), .B(n2259), .Z(n2261) );
  XOR U14412 ( .A(n2993), .B(n2994), .Z(n2259) );
  ANDN U14413 ( .B(n2995), .A(n2996), .Z(n2993) );
  AND U14414 ( .A(a[32]), .B(b[91]), .Z(n2992) );
  XNOR U14415 ( .A(n2997), .B(n2264), .Z(n2266) );
  XOR U14416 ( .A(n2998), .B(n2999), .Z(n2264) );
  ANDN U14417 ( .B(n3000), .A(n3001), .Z(n2998) );
  AND U14418 ( .A(a[33]), .B(b[90]), .Z(n2997) );
  XNOR U14419 ( .A(n3002), .B(n2269), .Z(n2271) );
  XOR U14420 ( .A(n3003), .B(n3004), .Z(n2269) );
  ANDN U14421 ( .B(n3005), .A(n3006), .Z(n3003) );
  AND U14422 ( .A(a[34]), .B(b[89]), .Z(n3002) );
  XNOR U14423 ( .A(n3007), .B(n2274), .Z(n2276) );
  XOR U14424 ( .A(n3008), .B(n3009), .Z(n2274) );
  ANDN U14425 ( .B(n3010), .A(n3011), .Z(n3008) );
  AND U14426 ( .A(a[35]), .B(b[88]), .Z(n3007) );
  XNOR U14427 ( .A(n3012), .B(n2279), .Z(n2281) );
  XOR U14428 ( .A(n3013), .B(n3014), .Z(n2279) );
  ANDN U14429 ( .B(n3015), .A(n3016), .Z(n3013) );
  AND U14430 ( .A(a[36]), .B(b[87]), .Z(n3012) );
  XNOR U14431 ( .A(n3017), .B(n2284), .Z(n2286) );
  XOR U14432 ( .A(n3018), .B(n3019), .Z(n2284) );
  ANDN U14433 ( .B(n3020), .A(n3021), .Z(n3018) );
  AND U14434 ( .A(a[37]), .B(b[86]), .Z(n3017) );
  XNOR U14435 ( .A(n3022), .B(n2289), .Z(n2291) );
  XOR U14436 ( .A(n3023), .B(n3024), .Z(n2289) );
  ANDN U14437 ( .B(n3025), .A(n3026), .Z(n3023) );
  AND U14438 ( .A(a[38]), .B(b[85]), .Z(n3022) );
  XNOR U14439 ( .A(n3027), .B(n2294), .Z(n2296) );
  XOR U14440 ( .A(n3028), .B(n3029), .Z(n2294) );
  ANDN U14441 ( .B(n3030), .A(n3031), .Z(n3028) );
  AND U14442 ( .A(a[39]), .B(b[84]), .Z(n3027) );
  XNOR U14443 ( .A(n3032), .B(n2299), .Z(n2301) );
  XOR U14444 ( .A(n3033), .B(n3034), .Z(n2299) );
  ANDN U14445 ( .B(n3035), .A(n3036), .Z(n3033) );
  AND U14446 ( .A(a[40]), .B(b[83]), .Z(n3032) );
  XNOR U14447 ( .A(n3037), .B(n2304), .Z(n2306) );
  XOR U14448 ( .A(n3038), .B(n3039), .Z(n2304) );
  ANDN U14449 ( .B(n3040), .A(n3041), .Z(n3038) );
  AND U14450 ( .A(a[41]), .B(b[82]), .Z(n3037) );
  XNOR U14451 ( .A(n3042), .B(n2309), .Z(n2311) );
  XOR U14452 ( .A(n3043), .B(n3044), .Z(n2309) );
  ANDN U14453 ( .B(n3045), .A(n3046), .Z(n3043) );
  AND U14454 ( .A(a[42]), .B(b[81]), .Z(n3042) );
  XNOR U14455 ( .A(n3047), .B(n2314), .Z(n2316) );
  XOR U14456 ( .A(n3048), .B(n3049), .Z(n2314) );
  ANDN U14457 ( .B(n3050), .A(n3051), .Z(n3048) );
  AND U14458 ( .A(a[43]), .B(b[80]), .Z(n3047) );
  XNOR U14459 ( .A(n3052), .B(n2319), .Z(n2321) );
  XOR U14460 ( .A(n3053), .B(n3054), .Z(n2319) );
  ANDN U14461 ( .B(n3055), .A(n3056), .Z(n3053) );
  AND U14462 ( .A(a[44]), .B(b[79]), .Z(n3052) );
  XNOR U14463 ( .A(n3057), .B(n2324), .Z(n2326) );
  XOR U14464 ( .A(n3058), .B(n3059), .Z(n2324) );
  ANDN U14465 ( .B(n3060), .A(n3061), .Z(n3058) );
  AND U14466 ( .A(a[45]), .B(b[78]), .Z(n3057) );
  XNOR U14467 ( .A(n3062), .B(n2329), .Z(n2331) );
  XOR U14468 ( .A(n3063), .B(n3064), .Z(n2329) );
  ANDN U14469 ( .B(n3065), .A(n3066), .Z(n3063) );
  AND U14470 ( .A(a[46]), .B(b[77]), .Z(n3062) );
  XNOR U14471 ( .A(n3067), .B(n2334), .Z(n2336) );
  XOR U14472 ( .A(n3068), .B(n3069), .Z(n2334) );
  ANDN U14473 ( .B(n3070), .A(n3071), .Z(n3068) );
  AND U14474 ( .A(a[47]), .B(b[76]), .Z(n3067) );
  XNOR U14475 ( .A(n3072), .B(n2339), .Z(n2341) );
  XOR U14476 ( .A(n3073), .B(n3074), .Z(n2339) );
  ANDN U14477 ( .B(n3075), .A(n3076), .Z(n3073) );
  AND U14478 ( .A(a[48]), .B(b[75]), .Z(n3072) );
  XNOR U14479 ( .A(n3077), .B(n2344), .Z(n2346) );
  XOR U14480 ( .A(n3078), .B(n3079), .Z(n2344) );
  ANDN U14481 ( .B(n3080), .A(n3081), .Z(n3078) );
  AND U14482 ( .A(a[49]), .B(b[74]), .Z(n3077) );
  XNOR U14483 ( .A(n3082), .B(n2349), .Z(n2351) );
  XOR U14484 ( .A(n3083), .B(n3084), .Z(n2349) );
  ANDN U14485 ( .B(n3085), .A(n3086), .Z(n3083) );
  AND U14486 ( .A(a[50]), .B(b[73]), .Z(n3082) );
  XNOR U14487 ( .A(n3087), .B(n2354), .Z(n2356) );
  XOR U14488 ( .A(n3088), .B(n3089), .Z(n2354) );
  ANDN U14489 ( .B(n3090), .A(n3091), .Z(n3088) );
  AND U14490 ( .A(a[51]), .B(b[72]), .Z(n3087) );
  XNOR U14491 ( .A(n3092), .B(n2359), .Z(n2361) );
  XOR U14492 ( .A(n3093), .B(n3094), .Z(n2359) );
  ANDN U14493 ( .B(n3095), .A(n3096), .Z(n3093) );
  AND U14494 ( .A(a[52]), .B(b[71]), .Z(n3092) );
  XNOR U14495 ( .A(n3097), .B(n2364), .Z(n2366) );
  XOR U14496 ( .A(n3098), .B(n3099), .Z(n2364) );
  ANDN U14497 ( .B(n3100), .A(n3101), .Z(n3098) );
  AND U14498 ( .A(a[53]), .B(b[70]), .Z(n3097) );
  XNOR U14499 ( .A(n3102), .B(n2369), .Z(n2371) );
  XOR U14500 ( .A(n3103), .B(n3104), .Z(n2369) );
  ANDN U14501 ( .B(n3105), .A(n3106), .Z(n3103) );
  AND U14502 ( .A(a[54]), .B(b[69]), .Z(n3102) );
  XNOR U14503 ( .A(n3107), .B(n2374), .Z(n2376) );
  XOR U14504 ( .A(n3108), .B(n3109), .Z(n2374) );
  ANDN U14505 ( .B(n3110), .A(n3111), .Z(n3108) );
  AND U14506 ( .A(a[55]), .B(b[68]), .Z(n3107) );
  XNOR U14507 ( .A(n3112), .B(n2379), .Z(n2381) );
  XOR U14508 ( .A(n3113), .B(n3114), .Z(n2379) );
  ANDN U14509 ( .B(n3115), .A(n3116), .Z(n3113) );
  AND U14510 ( .A(a[56]), .B(b[67]), .Z(n3112) );
  XNOR U14511 ( .A(n3117), .B(n2384), .Z(n2386) );
  XOR U14512 ( .A(n3118), .B(n3119), .Z(n2384) );
  ANDN U14513 ( .B(n3120), .A(n3121), .Z(n3118) );
  AND U14514 ( .A(a[57]), .B(b[66]), .Z(n3117) );
  XNOR U14515 ( .A(n3122), .B(n2389), .Z(n2391) );
  XOR U14516 ( .A(n3123), .B(n3124), .Z(n2389) );
  ANDN U14517 ( .B(n3125), .A(n3126), .Z(n3123) );
  AND U14518 ( .A(a[58]), .B(b[65]), .Z(n3122) );
  XNOR U14519 ( .A(n3127), .B(n2394), .Z(n2396) );
  XOR U14520 ( .A(n3128), .B(n3129), .Z(n2394) );
  ANDN U14521 ( .B(n3130), .A(n3131), .Z(n3128) );
  AND U14522 ( .A(a[59]), .B(b[64]), .Z(n3127) );
  XNOR U14523 ( .A(n3132), .B(n2399), .Z(n2401) );
  XOR U14524 ( .A(n3133), .B(n3134), .Z(n2399) );
  ANDN U14525 ( .B(n3135), .A(n3136), .Z(n3133) );
  AND U14526 ( .A(a[60]), .B(b[63]), .Z(n3132) );
  XNOR U14527 ( .A(n3137), .B(n2404), .Z(n2406) );
  XOR U14528 ( .A(n3138), .B(n3139), .Z(n2404) );
  ANDN U14529 ( .B(n3140), .A(n3141), .Z(n3138) );
  AND U14530 ( .A(a[61]), .B(b[62]), .Z(n3137) );
  XNOR U14531 ( .A(n3142), .B(n2409), .Z(n2411) );
  XOR U14532 ( .A(n3143), .B(n3144), .Z(n2409) );
  ANDN U14533 ( .B(n3145), .A(n3146), .Z(n3143) );
  AND U14534 ( .A(a[62]), .B(b[61]), .Z(n3142) );
  XNOR U14535 ( .A(n3147), .B(n2414), .Z(n2416) );
  XOR U14536 ( .A(n3148), .B(n3149), .Z(n2414) );
  ANDN U14537 ( .B(n3150), .A(n3151), .Z(n3148) );
  AND U14538 ( .A(a[63]), .B(b[60]), .Z(n3147) );
  XNOR U14539 ( .A(n3152), .B(n2419), .Z(n2421) );
  XOR U14540 ( .A(n3153), .B(n3154), .Z(n2419) );
  ANDN U14541 ( .B(n3155), .A(n3156), .Z(n3153) );
  AND U14542 ( .A(a[64]), .B(b[59]), .Z(n3152) );
  XNOR U14543 ( .A(n3157), .B(n2424), .Z(n2426) );
  XOR U14544 ( .A(n3158), .B(n3159), .Z(n2424) );
  ANDN U14545 ( .B(n3160), .A(n3161), .Z(n3158) );
  AND U14546 ( .A(a[65]), .B(b[58]), .Z(n3157) );
  XNOR U14547 ( .A(n3162), .B(n2429), .Z(n2431) );
  XOR U14548 ( .A(n3163), .B(n3164), .Z(n2429) );
  ANDN U14549 ( .B(n3165), .A(n3166), .Z(n3163) );
  AND U14550 ( .A(a[66]), .B(b[57]), .Z(n3162) );
  XNOR U14551 ( .A(n3167), .B(n2434), .Z(n2436) );
  XOR U14552 ( .A(n3168), .B(n3169), .Z(n2434) );
  ANDN U14553 ( .B(n3170), .A(n3171), .Z(n3168) );
  AND U14554 ( .A(a[67]), .B(b[56]), .Z(n3167) );
  XNOR U14555 ( .A(n3172), .B(n2439), .Z(n2441) );
  XOR U14556 ( .A(n3173), .B(n3174), .Z(n2439) );
  ANDN U14557 ( .B(n3175), .A(n3176), .Z(n3173) );
  AND U14558 ( .A(a[68]), .B(b[55]), .Z(n3172) );
  XNOR U14559 ( .A(n3177), .B(n2444), .Z(n2446) );
  XOR U14560 ( .A(n3178), .B(n3179), .Z(n2444) );
  ANDN U14561 ( .B(n3180), .A(n3181), .Z(n3178) );
  AND U14562 ( .A(a[69]), .B(b[54]), .Z(n3177) );
  XNOR U14563 ( .A(n3182), .B(n2449), .Z(n2451) );
  XOR U14564 ( .A(n3183), .B(n3184), .Z(n2449) );
  ANDN U14565 ( .B(n3185), .A(n3186), .Z(n3183) );
  AND U14566 ( .A(a[70]), .B(b[53]), .Z(n3182) );
  XNOR U14567 ( .A(n3187), .B(n2454), .Z(n2456) );
  XOR U14568 ( .A(n3188), .B(n3189), .Z(n2454) );
  ANDN U14569 ( .B(n3190), .A(n3191), .Z(n3188) );
  AND U14570 ( .A(a[71]), .B(b[52]), .Z(n3187) );
  XNOR U14571 ( .A(n3192), .B(n2459), .Z(n2461) );
  XOR U14572 ( .A(n3193), .B(n3194), .Z(n2459) );
  ANDN U14573 ( .B(n3195), .A(n3196), .Z(n3193) );
  AND U14574 ( .A(a[72]), .B(b[51]), .Z(n3192) );
  XNOR U14575 ( .A(n3197), .B(n2464), .Z(n2466) );
  XOR U14576 ( .A(n3198), .B(n3199), .Z(n2464) );
  ANDN U14577 ( .B(n3200), .A(n3201), .Z(n3198) );
  AND U14578 ( .A(a[73]), .B(b[50]), .Z(n3197) );
  XNOR U14579 ( .A(n3202), .B(n2469), .Z(n2471) );
  XOR U14580 ( .A(n3203), .B(n3204), .Z(n2469) );
  ANDN U14581 ( .B(n3205), .A(n3206), .Z(n3203) );
  AND U14582 ( .A(a[74]), .B(b[49]), .Z(n3202) );
  XNOR U14583 ( .A(n3207), .B(n2474), .Z(n2476) );
  XOR U14584 ( .A(n3208), .B(n3209), .Z(n2474) );
  ANDN U14585 ( .B(n3210), .A(n3211), .Z(n3208) );
  AND U14586 ( .A(a[75]), .B(b[48]), .Z(n3207) );
  XNOR U14587 ( .A(n3212), .B(n2479), .Z(n2481) );
  XOR U14588 ( .A(n3213), .B(n3214), .Z(n2479) );
  ANDN U14589 ( .B(n3215), .A(n3216), .Z(n3213) );
  AND U14590 ( .A(a[76]), .B(b[47]), .Z(n3212) );
  XNOR U14591 ( .A(n3217), .B(n2484), .Z(n2486) );
  XOR U14592 ( .A(n3218), .B(n3219), .Z(n2484) );
  ANDN U14593 ( .B(n3220), .A(n3221), .Z(n3218) );
  AND U14594 ( .A(a[77]), .B(b[46]), .Z(n3217) );
  XNOR U14595 ( .A(n3222), .B(n2489), .Z(n2491) );
  XOR U14596 ( .A(n3223), .B(n3224), .Z(n2489) );
  ANDN U14597 ( .B(n3225), .A(n3226), .Z(n3223) );
  AND U14598 ( .A(a[78]), .B(b[45]), .Z(n3222) );
  XNOR U14599 ( .A(n3227), .B(n2494), .Z(n2496) );
  XOR U14600 ( .A(n3228), .B(n3229), .Z(n2494) );
  ANDN U14601 ( .B(n3230), .A(n3231), .Z(n3228) );
  AND U14602 ( .A(a[79]), .B(b[44]), .Z(n3227) );
  XNOR U14603 ( .A(n3232), .B(n2499), .Z(n2501) );
  XOR U14604 ( .A(n3233), .B(n3234), .Z(n2499) );
  ANDN U14605 ( .B(n3235), .A(n3236), .Z(n3233) );
  AND U14606 ( .A(a[80]), .B(b[43]), .Z(n3232) );
  XNOR U14607 ( .A(n3237), .B(n2504), .Z(n2506) );
  XOR U14608 ( .A(n3238), .B(n3239), .Z(n2504) );
  ANDN U14609 ( .B(n3240), .A(n3241), .Z(n3238) );
  AND U14610 ( .A(a[81]), .B(b[42]), .Z(n3237) );
  XNOR U14611 ( .A(n3242), .B(n2509), .Z(n2511) );
  XOR U14612 ( .A(n3243), .B(n3244), .Z(n2509) );
  ANDN U14613 ( .B(n3245), .A(n3246), .Z(n3243) );
  AND U14614 ( .A(a[82]), .B(b[41]), .Z(n3242) );
  XNOR U14615 ( .A(n3247), .B(n2514), .Z(n2516) );
  XOR U14616 ( .A(n3248), .B(n3249), .Z(n2514) );
  ANDN U14617 ( .B(n3250), .A(n3251), .Z(n3248) );
  AND U14618 ( .A(a[83]), .B(b[40]), .Z(n3247) );
  XNOR U14619 ( .A(n3252), .B(n2519), .Z(n2521) );
  XOR U14620 ( .A(n3253), .B(n3254), .Z(n2519) );
  ANDN U14621 ( .B(n3255), .A(n3256), .Z(n3253) );
  AND U14622 ( .A(a[84]), .B(b[39]), .Z(n3252) );
  XNOR U14623 ( .A(n3257), .B(n2524), .Z(n2526) );
  XOR U14624 ( .A(n3258), .B(n3259), .Z(n2524) );
  ANDN U14625 ( .B(n3260), .A(n3261), .Z(n3258) );
  AND U14626 ( .A(a[85]), .B(b[38]), .Z(n3257) );
  XNOR U14627 ( .A(n3262), .B(n2529), .Z(n2531) );
  XOR U14628 ( .A(n3263), .B(n3264), .Z(n2529) );
  ANDN U14629 ( .B(n3265), .A(n3266), .Z(n3263) );
  AND U14630 ( .A(a[86]), .B(b[37]), .Z(n3262) );
  XNOR U14631 ( .A(n3267), .B(n2534), .Z(n2536) );
  XOR U14632 ( .A(n3268), .B(n3269), .Z(n2534) );
  ANDN U14633 ( .B(n3270), .A(n3271), .Z(n3268) );
  AND U14634 ( .A(a[87]), .B(b[36]), .Z(n3267) );
  XNOR U14635 ( .A(n3272), .B(n2539), .Z(n2541) );
  XOR U14636 ( .A(n3273), .B(n3274), .Z(n2539) );
  ANDN U14637 ( .B(n3275), .A(n3276), .Z(n3273) );
  AND U14638 ( .A(a[88]), .B(b[35]), .Z(n3272) );
  XNOR U14639 ( .A(n3277), .B(n2544), .Z(n2546) );
  XOR U14640 ( .A(n3278), .B(n3279), .Z(n2544) );
  ANDN U14641 ( .B(n3280), .A(n3281), .Z(n3278) );
  AND U14642 ( .A(a[89]), .B(b[34]), .Z(n3277) );
  XNOR U14643 ( .A(n3282), .B(n2549), .Z(n2551) );
  XOR U14644 ( .A(n3283), .B(n3284), .Z(n2549) );
  ANDN U14645 ( .B(n3285), .A(n3286), .Z(n3283) );
  AND U14646 ( .A(a[90]), .B(b[33]), .Z(n3282) );
  XNOR U14647 ( .A(n3287), .B(n2554), .Z(n2556) );
  XOR U14648 ( .A(n3288), .B(n3289), .Z(n2554) );
  ANDN U14649 ( .B(n3290), .A(n3291), .Z(n3288) );
  AND U14650 ( .A(a[91]), .B(b[32]), .Z(n3287) );
  XNOR U14651 ( .A(n3292), .B(n2559), .Z(n2561) );
  XOR U14652 ( .A(n3293), .B(n3294), .Z(n2559) );
  ANDN U14653 ( .B(n3295), .A(n3296), .Z(n3293) );
  AND U14654 ( .A(a[92]), .B(b[31]), .Z(n3292) );
  XNOR U14655 ( .A(n3297), .B(n2564), .Z(n2566) );
  XOR U14656 ( .A(n3298), .B(n3299), .Z(n2564) );
  ANDN U14657 ( .B(n3300), .A(n3301), .Z(n3298) );
  AND U14658 ( .A(a[93]), .B(b[30]), .Z(n3297) );
  XNOR U14659 ( .A(n3302), .B(n2569), .Z(n2571) );
  XOR U14660 ( .A(n3303), .B(n3304), .Z(n2569) );
  ANDN U14661 ( .B(n3305), .A(n3306), .Z(n3303) );
  AND U14662 ( .A(a[94]), .B(b[29]), .Z(n3302) );
  XNOR U14663 ( .A(n3307), .B(n2574), .Z(n2576) );
  XOR U14664 ( .A(n3308), .B(n3309), .Z(n2574) );
  ANDN U14665 ( .B(n3310), .A(n3311), .Z(n3308) );
  AND U14666 ( .A(a[95]), .B(b[28]), .Z(n3307) );
  XNOR U14667 ( .A(n3312), .B(n2579), .Z(n2581) );
  XOR U14668 ( .A(n3313), .B(n3314), .Z(n2579) );
  ANDN U14669 ( .B(n3315), .A(n3316), .Z(n3313) );
  AND U14670 ( .A(a[96]), .B(b[27]), .Z(n3312) );
  XNOR U14671 ( .A(n3317), .B(n2584), .Z(n2586) );
  XOR U14672 ( .A(n3318), .B(n3319), .Z(n2584) );
  ANDN U14673 ( .B(n3320), .A(n3321), .Z(n3318) );
  AND U14674 ( .A(a[97]), .B(b[26]), .Z(n3317) );
  XNOR U14675 ( .A(n3322), .B(n2589), .Z(n2591) );
  XOR U14676 ( .A(n3323), .B(n3324), .Z(n2589) );
  ANDN U14677 ( .B(n3325), .A(n3326), .Z(n3323) );
  AND U14678 ( .A(a[98]), .B(b[25]), .Z(n3322) );
  XNOR U14679 ( .A(n3327), .B(n2594), .Z(n2596) );
  XOR U14680 ( .A(n3328), .B(n3329), .Z(n2594) );
  ANDN U14681 ( .B(n3330), .A(n3331), .Z(n3328) );
  AND U14682 ( .A(a[99]), .B(b[24]), .Z(n3327) );
  XNOR U14683 ( .A(n3332), .B(n2599), .Z(n2601) );
  XOR U14684 ( .A(n3333), .B(n3334), .Z(n2599) );
  ANDN U14685 ( .B(n3335), .A(n3336), .Z(n3333) );
  AND U14686 ( .A(b[23]), .B(a[100]), .Z(n3332) );
  XNOR U14687 ( .A(n3337), .B(n2604), .Z(n2606) );
  XOR U14688 ( .A(n3338), .B(n3339), .Z(n2604) );
  ANDN U14689 ( .B(n3340), .A(n3341), .Z(n3338) );
  AND U14690 ( .A(b[22]), .B(a[101]), .Z(n3337) );
  XNOR U14691 ( .A(n3342), .B(n2609), .Z(n2611) );
  XOR U14692 ( .A(n3343), .B(n3344), .Z(n2609) );
  ANDN U14693 ( .B(n3345), .A(n3346), .Z(n3343) );
  AND U14694 ( .A(b[21]), .B(a[102]), .Z(n3342) );
  XNOR U14695 ( .A(n3347), .B(n2614), .Z(n2616) );
  XOR U14696 ( .A(n3348), .B(n3349), .Z(n2614) );
  ANDN U14697 ( .B(n3350), .A(n3351), .Z(n3348) );
  AND U14698 ( .A(b[20]), .B(a[103]), .Z(n3347) );
  XNOR U14699 ( .A(n3352), .B(n2619), .Z(n2621) );
  XOR U14700 ( .A(n3353), .B(n3354), .Z(n2619) );
  ANDN U14701 ( .B(n3355), .A(n3356), .Z(n3353) );
  AND U14702 ( .A(b[19]), .B(a[104]), .Z(n3352) );
  XNOR U14703 ( .A(n3357), .B(n2624), .Z(n2626) );
  XOR U14704 ( .A(n3358), .B(n3359), .Z(n2624) );
  ANDN U14705 ( .B(n3360), .A(n3361), .Z(n3358) );
  AND U14706 ( .A(b[18]), .B(a[105]), .Z(n3357) );
  XNOR U14707 ( .A(n3362), .B(n2629), .Z(n2631) );
  XOR U14708 ( .A(n3363), .B(n3364), .Z(n2629) );
  ANDN U14709 ( .B(n3365), .A(n3366), .Z(n3363) );
  AND U14710 ( .A(b[17]), .B(a[106]), .Z(n3362) );
  XNOR U14711 ( .A(n3367), .B(n2634), .Z(n2636) );
  XOR U14712 ( .A(n3368), .B(n3369), .Z(n2634) );
  ANDN U14713 ( .B(n3370), .A(n3371), .Z(n3368) );
  AND U14714 ( .A(b[16]), .B(a[107]), .Z(n3367) );
  XNOR U14715 ( .A(n3372), .B(n2639), .Z(n2641) );
  XOR U14716 ( .A(n3373), .B(n3374), .Z(n2639) );
  ANDN U14717 ( .B(n3375), .A(n3376), .Z(n3373) );
  AND U14718 ( .A(b[15]), .B(a[108]), .Z(n3372) );
  XNOR U14719 ( .A(n3377), .B(n2644), .Z(n2646) );
  XOR U14720 ( .A(n3378), .B(n3379), .Z(n2644) );
  ANDN U14721 ( .B(n3380), .A(n3381), .Z(n3378) );
  AND U14722 ( .A(b[14]), .B(a[109]), .Z(n3377) );
  XNOR U14723 ( .A(n3382), .B(n2649), .Z(n2651) );
  XOR U14724 ( .A(n3383), .B(n3384), .Z(n2649) );
  ANDN U14725 ( .B(n3385), .A(n3386), .Z(n3383) );
  AND U14726 ( .A(b[13]), .B(a[110]), .Z(n3382) );
  XNOR U14727 ( .A(n3387), .B(n2654), .Z(n2656) );
  XOR U14728 ( .A(n3388), .B(n3389), .Z(n2654) );
  ANDN U14729 ( .B(n3390), .A(n3391), .Z(n3388) );
  AND U14730 ( .A(b[12]), .B(a[111]), .Z(n3387) );
  XNOR U14731 ( .A(n3392), .B(n2659), .Z(n2661) );
  XOR U14732 ( .A(n3393), .B(n3394), .Z(n2659) );
  ANDN U14733 ( .B(n3395), .A(n3396), .Z(n3393) );
  AND U14734 ( .A(b[11]), .B(a[112]), .Z(n3392) );
  XNOR U14735 ( .A(n3397), .B(n2664), .Z(n2666) );
  XOR U14736 ( .A(n3398), .B(n3399), .Z(n2664) );
  ANDN U14737 ( .B(n3400), .A(n3401), .Z(n3398) );
  AND U14738 ( .A(b[10]), .B(a[113]), .Z(n3397) );
  XNOR U14739 ( .A(n3402), .B(n2669), .Z(n2671) );
  XOR U14740 ( .A(n3403), .B(n3404), .Z(n2669) );
  ANDN U14741 ( .B(n3405), .A(n3406), .Z(n3403) );
  AND U14742 ( .A(b[9]), .B(a[114]), .Z(n3402) );
  XNOR U14743 ( .A(n3407), .B(n2674), .Z(n2676) );
  XOR U14744 ( .A(n3408), .B(n3409), .Z(n2674) );
  ANDN U14745 ( .B(n3410), .A(n3411), .Z(n3408) );
  AND U14746 ( .A(b[8]), .B(a[115]), .Z(n3407) );
  XNOR U14747 ( .A(n3412), .B(n2679), .Z(n2681) );
  XOR U14748 ( .A(n3413), .B(n3414), .Z(n2679) );
  ANDN U14749 ( .B(n3415), .A(n3416), .Z(n3413) );
  AND U14750 ( .A(b[7]), .B(a[116]), .Z(n3412) );
  XNOR U14751 ( .A(n3417), .B(n2684), .Z(n2686) );
  XOR U14752 ( .A(n3418), .B(n3419), .Z(n2684) );
  ANDN U14753 ( .B(n3420), .A(n3421), .Z(n3418) );
  AND U14754 ( .A(b[6]), .B(a[117]), .Z(n3417) );
  XNOR U14755 ( .A(n3422), .B(n2689), .Z(n2691) );
  XOR U14756 ( .A(n3423), .B(n3424), .Z(n2689) );
  ANDN U14757 ( .B(n3425), .A(n3426), .Z(n3423) );
  AND U14758 ( .A(b[5]), .B(a[118]), .Z(n3422) );
  XNOR U14759 ( .A(n3427), .B(n2694), .Z(n2696) );
  XOR U14760 ( .A(n3428), .B(n3429), .Z(n2694) );
  ANDN U14761 ( .B(n3430), .A(n3431), .Z(n3428) );
  AND U14762 ( .A(b[4]), .B(a[119]), .Z(n3427) );
  XNOR U14763 ( .A(n3432), .B(n3433), .Z(n2708) );
  NANDN U14764 ( .A(n3434), .B(n3435), .Z(n3433) );
  XNOR U14765 ( .A(n3436), .B(n2699), .Z(n2701) );
  XNOR U14766 ( .A(n3437), .B(n3438), .Z(n2699) );
  AND U14767 ( .A(n3439), .B(n3440), .Z(n3437) );
  AND U14768 ( .A(b[3]), .B(a[120]), .Z(n3436) );
  NAND U14769 ( .A(a[123]), .B(b[0]), .Z(n1978) );
  XNOR U14770 ( .A(n2714), .B(n2715), .Z(c[122]) );
  XNOR U14771 ( .A(n3434), .B(n3435), .Z(n2715) );
  XOR U14772 ( .A(n3432), .B(n3441), .Z(n3435) );
  NAND U14773 ( .A(b[1]), .B(a[121]), .Z(n3441) );
  XOR U14774 ( .A(n3440), .B(n3442), .Z(n3434) );
  XOR U14775 ( .A(n3432), .B(n3439), .Z(n3442) );
  XNOR U14776 ( .A(n3443), .B(n3438), .Z(n3439) );
  AND U14777 ( .A(b[2]), .B(a[120]), .Z(n3443) );
  NANDN U14778 ( .A(n3444), .B(n3445), .Z(n3432) );
  XOR U14779 ( .A(n3438), .B(n3430), .Z(n3446) );
  XNOR U14780 ( .A(n3429), .B(n3425), .Z(n3447) );
  XNOR U14781 ( .A(n3424), .B(n3420), .Z(n3448) );
  XNOR U14782 ( .A(n3419), .B(n3415), .Z(n3449) );
  XNOR U14783 ( .A(n3414), .B(n3410), .Z(n3450) );
  XNOR U14784 ( .A(n3409), .B(n3405), .Z(n3451) );
  XNOR U14785 ( .A(n3404), .B(n3400), .Z(n3452) );
  XNOR U14786 ( .A(n3399), .B(n3395), .Z(n3453) );
  XNOR U14787 ( .A(n3394), .B(n3390), .Z(n3454) );
  XNOR U14788 ( .A(n3389), .B(n3385), .Z(n3455) );
  XNOR U14789 ( .A(n3384), .B(n3380), .Z(n3456) );
  XNOR U14790 ( .A(n3379), .B(n3375), .Z(n3457) );
  XNOR U14791 ( .A(n3374), .B(n3370), .Z(n3458) );
  XNOR U14792 ( .A(n3369), .B(n3365), .Z(n3459) );
  XNOR U14793 ( .A(n3364), .B(n3360), .Z(n3460) );
  XNOR U14794 ( .A(n3359), .B(n3355), .Z(n3461) );
  XNOR U14795 ( .A(n3354), .B(n3350), .Z(n3462) );
  XNOR U14796 ( .A(n3349), .B(n3345), .Z(n3463) );
  XNOR U14797 ( .A(n3344), .B(n3340), .Z(n3464) );
  XNOR U14798 ( .A(n3339), .B(n3335), .Z(n3465) );
  XNOR U14799 ( .A(n3334), .B(n3330), .Z(n3466) );
  XNOR U14800 ( .A(n3329), .B(n3325), .Z(n3467) );
  XNOR U14801 ( .A(n3324), .B(n3320), .Z(n3468) );
  XNOR U14802 ( .A(n3319), .B(n3315), .Z(n3469) );
  XNOR U14803 ( .A(n3314), .B(n3310), .Z(n3470) );
  XNOR U14804 ( .A(n3309), .B(n3305), .Z(n3471) );
  XNOR U14805 ( .A(n3304), .B(n3300), .Z(n3472) );
  XNOR U14806 ( .A(n3299), .B(n3295), .Z(n3473) );
  XNOR U14807 ( .A(n3294), .B(n3290), .Z(n3474) );
  XNOR U14808 ( .A(n3289), .B(n3285), .Z(n3475) );
  XNOR U14809 ( .A(n3284), .B(n3280), .Z(n3476) );
  XNOR U14810 ( .A(n3279), .B(n3275), .Z(n3477) );
  XNOR U14811 ( .A(n3274), .B(n3270), .Z(n3478) );
  XNOR U14812 ( .A(n3269), .B(n3265), .Z(n3479) );
  XNOR U14813 ( .A(n3264), .B(n3260), .Z(n3480) );
  XNOR U14814 ( .A(n3259), .B(n3255), .Z(n3481) );
  XNOR U14815 ( .A(n3254), .B(n3250), .Z(n3482) );
  XNOR U14816 ( .A(n3249), .B(n3245), .Z(n3483) );
  XNOR U14817 ( .A(n3244), .B(n3240), .Z(n3484) );
  XNOR U14818 ( .A(n3239), .B(n3235), .Z(n3485) );
  XNOR U14819 ( .A(n3234), .B(n3230), .Z(n3486) );
  XNOR U14820 ( .A(n3229), .B(n3225), .Z(n3487) );
  XNOR U14821 ( .A(n3224), .B(n3220), .Z(n3488) );
  XNOR U14822 ( .A(n3219), .B(n3215), .Z(n3489) );
  XNOR U14823 ( .A(n3214), .B(n3210), .Z(n3490) );
  XNOR U14824 ( .A(n3209), .B(n3205), .Z(n3491) );
  XNOR U14825 ( .A(n3204), .B(n3200), .Z(n3492) );
  XNOR U14826 ( .A(n3199), .B(n3195), .Z(n3493) );
  XNOR U14827 ( .A(n3194), .B(n3190), .Z(n3494) );
  XNOR U14828 ( .A(n3189), .B(n3185), .Z(n3495) );
  XNOR U14829 ( .A(n3184), .B(n3180), .Z(n3496) );
  XNOR U14830 ( .A(n3179), .B(n3175), .Z(n3497) );
  XNOR U14831 ( .A(n3174), .B(n3170), .Z(n3498) );
  XNOR U14832 ( .A(n3169), .B(n3165), .Z(n3499) );
  XNOR U14833 ( .A(n3164), .B(n3160), .Z(n3500) );
  XNOR U14834 ( .A(n3159), .B(n3155), .Z(n3501) );
  XNOR U14835 ( .A(n3154), .B(n3150), .Z(n3502) );
  XNOR U14836 ( .A(n3149), .B(n3145), .Z(n3503) );
  XNOR U14837 ( .A(n3144), .B(n3140), .Z(n3504) );
  XNOR U14838 ( .A(n3139), .B(n3135), .Z(n3505) );
  XNOR U14839 ( .A(n3134), .B(n3130), .Z(n3506) );
  XNOR U14840 ( .A(n3129), .B(n3125), .Z(n3507) );
  XNOR U14841 ( .A(n3124), .B(n3120), .Z(n3508) );
  XNOR U14842 ( .A(n3119), .B(n3115), .Z(n3509) );
  XNOR U14843 ( .A(n3114), .B(n3110), .Z(n3510) );
  XNOR U14844 ( .A(n3109), .B(n3105), .Z(n3511) );
  XNOR U14845 ( .A(n3104), .B(n3100), .Z(n3512) );
  XNOR U14846 ( .A(n3099), .B(n3095), .Z(n3513) );
  XNOR U14847 ( .A(n3094), .B(n3090), .Z(n3514) );
  XNOR U14848 ( .A(n3089), .B(n3085), .Z(n3515) );
  XNOR U14849 ( .A(n3084), .B(n3080), .Z(n3516) );
  XNOR U14850 ( .A(n3079), .B(n3075), .Z(n3517) );
  XNOR U14851 ( .A(n3074), .B(n3070), .Z(n3518) );
  XNOR U14852 ( .A(n3069), .B(n3065), .Z(n3519) );
  XNOR U14853 ( .A(n3064), .B(n3060), .Z(n3520) );
  XNOR U14854 ( .A(n3059), .B(n3055), .Z(n3521) );
  XNOR U14855 ( .A(n3054), .B(n3050), .Z(n3522) );
  XNOR U14856 ( .A(n3049), .B(n3045), .Z(n3523) );
  XNOR U14857 ( .A(n3044), .B(n3040), .Z(n3524) );
  XNOR U14858 ( .A(n3039), .B(n3035), .Z(n3525) );
  XNOR U14859 ( .A(n3034), .B(n3030), .Z(n3526) );
  XNOR U14860 ( .A(n3029), .B(n3025), .Z(n3527) );
  XNOR U14861 ( .A(n3024), .B(n3020), .Z(n3528) );
  XNOR U14862 ( .A(n3019), .B(n3015), .Z(n3529) );
  XNOR U14863 ( .A(n3014), .B(n3010), .Z(n3530) );
  XNOR U14864 ( .A(n3009), .B(n3005), .Z(n3531) );
  XNOR U14865 ( .A(n3004), .B(n3000), .Z(n3532) );
  XNOR U14866 ( .A(n2999), .B(n2995), .Z(n3533) );
  XNOR U14867 ( .A(n2994), .B(n2990), .Z(n3534) );
  XNOR U14868 ( .A(n2989), .B(n2985), .Z(n3535) );
  XNOR U14869 ( .A(n2984), .B(n2980), .Z(n3536) );
  XNOR U14870 ( .A(n2979), .B(n2975), .Z(n3537) );
  XNOR U14871 ( .A(n2974), .B(n2970), .Z(n3538) );
  XNOR U14872 ( .A(n2969), .B(n2965), .Z(n3539) );
  XNOR U14873 ( .A(n2964), .B(n2960), .Z(n3540) );
  XNOR U14874 ( .A(n2959), .B(n2955), .Z(n3541) );
  XNOR U14875 ( .A(n2954), .B(n2950), .Z(n3542) );
  XNOR U14876 ( .A(n2949), .B(n2945), .Z(n3543) );
  XNOR U14877 ( .A(n2944), .B(n2940), .Z(n3544) );
  XNOR U14878 ( .A(n2939), .B(n2935), .Z(n3545) );
  XNOR U14879 ( .A(n2934), .B(n2930), .Z(n3546) );
  XNOR U14880 ( .A(n2929), .B(n2925), .Z(n3547) );
  XNOR U14881 ( .A(n2924), .B(n2920), .Z(n3548) );
  XNOR U14882 ( .A(n2919), .B(n2915), .Z(n3549) );
  XNOR U14883 ( .A(n2914), .B(n2910), .Z(n3550) );
  XNOR U14884 ( .A(n2909), .B(n2905), .Z(n3551) );
  XNOR U14885 ( .A(n2904), .B(n2900), .Z(n3552) );
  XNOR U14886 ( .A(n2899), .B(n2895), .Z(n3553) );
  XNOR U14887 ( .A(n2894), .B(n2890), .Z(n3554) );
  XNOR U14888 ( .A(n2889), .B(n2885), .Z(n3555) );
  XNOR U14889 ( .A(n2884), .B(n2880), .Z(n3556) );
  XNOR U14890 ( .A(n2879), .B(n2875), .Z(n3557) );
  XNOR U14891 ( .A(n2874), .B(n2870), .Z(n3558) );
  XNOR U14892 ( .A(n2869), .B(n2865), .Z(n3559) );
  XNOR U14893 ( .A(n2864), .B(n2860), .Z(n3560) );
  XNOR U14894 ( .A(n2859), .B(n2855), .Z(n3561) );
  XNOR U14895 ( .A(n2854), .B(n2850), .Z(n3562) );
  XNOR U14896 ( .A(n2849), .B(n2845), .Z(n3563) );
  XNOR U14897 ( .A(n2844), .B(n2840), .Z(n3564) );
  XOR U14898 ( .A(n3565), .B(n2839), .Z(n2840) );
  AND U14899 ( .A(a[0]), .B(b[122]), .Z(n3565) );
  XNOR U14900 ( .A(n3566), .B(n2839), .Z(n2841) );
  XNOR U14901 ( .A(n3567), .B(n3568), .Z(n2839) );
  ANDN U14902 ( .B(n3569), .A(n3570), .Z(n3567) );
  AND U14903 ( .A(a[1]), .B(b[121]), .Z(n3566) );
  XNOR U14904 ( .A(n3571), .B(n2844), .Z(n2846) );
  XOR U14905 ( .A(n3572), .B(n3573), .Z(n2844) );
  ANDN U14906 ( .B(n3574), .A(n3575), .Z(n3572) );
  AND U14907 ( .A(a[2]), .B(b[120]), .Z(n3571) );
  XNOR U14908 ( .A(n3576), .B(n2849), .Z(n2851) );
  XOR U14909 ( .A(n3577), .B(n3578), .Z(n2849) );
  ANDN U14910 ( .B(n3579), .A(n3580), .Z(n3577) );
  AND U14911 ( .A(a[3]), .B(b[119]), .Z(n3576) );
  XNOR U14912 ( .A(n3581), .B(n2854), .Z(n2856) );
  XOR U14913 ( .A(n3582), .B(n3583), .Z(n2854) );
  ANDN U14914 ( .B(n3584), .A(n3585), .Z(n3582) );
  AND U14915 ( .A(a[4]), .B(b[118]), .Z(n3581) );
  XNOR U14916 ( .A(n3586), .B(n2859), .Z(n2861) );
  XOR U14917 ( .A(n3587), .B(n3588), .Z(n2859) );
  ANDN U14918 ( .B(n3589), .A(n3590), .Z(n3587) );
  AND U14919 ( .A(a[5]), .B(b[117]), .Z(n3586) );
  XNOR U14920 ( .A(n3591), .B(n2864), .Z(n2866) );
  XOR U14921 ( .A(n3592), .B(n3593), .Z(n2864) );
  ANDN U14922 ( .B(n3594), .A(n3595), .Z(n3592) );
  AND U14923 ( .A(a[6]), .B(b[116]), .Z(n3591) );
  XNOR U14924 ( .A(n3596), .B(n2869), .Z(n2871) );
  XOR U14925 ( .A(n3597), .B(n3598), .Z(n2869) );
  ANDN U14926 ( .B(n3599), .A(n3600), .Z(n3597) );
  AND U14927 ( .A(a[7]), .B(b[115]), .Z(n3596) );
  XNOR U14928 ( .A(n3601), .B(n2874), .Z(n2876) );
  XOR U14929 ( .A(n3602), .B(n3603), .Z(n2874) );
  ANDN U14930 ( .B(n3604), .A(n3605), .Z(n3602) );
  AND U14931 ( .A(a[8]), .B(b[114]), .Z(n3601) );
  XNOR U14932 ( .A(n3606), .B(n2879), .Z(n2881) );
  XOR U14933 ( .A(n3607), .B(n3608), .Z(n2879) );
  ANDN U14934 ( .B(n3609), .A(n3610), .Z(n3607) );
  AND U14935 ( .A(a[9]), .B(b[113]), .Z(n3606) );
  XNOR U14936 ( .A(n3611), .B(n2884), .Z(n2886) );
  XOR U14937 ( .A(n3612), .B(n3613), .Z(n2884) );
  ANDN U14938 ( .B(n3614), .A(n3615), .Z(n3612) );
  AND U14939 ( .A(a[10]), .B(b[112]), .Z(n3611) );
  XNOR U14940 ( .A(n3616), .B(n2889), .Z(n2891) );
  XOR U14941 ( .A(n3617), .B(n3618), .Z(n2889) );
  ANDN U14942 ( .B(n3619), .A(n3620), .Z(n3617) );
  AND U14943 ( .A(a[11]), .B(b[111]), .Z(n3616) );
  XNOR U14944 ( .A(n3621), .B(n2894), .Z(n2896) );
  XOR U14945 ( .A(n3622), .B(n3623), .Z(n2894) );
  ANDN U14946 ( .B(n3624), .A(n3625), .Z(n3622) );
  AND U14947 ( .A(a[12]), .B(b[110]), .Z(n3621) );
  XNOR U14948 ( .A(n3626), .B(n2899), .Z(n2901) );
  XOR U14949 ( .A(n3627), .B(n3628), .Z(n2899) );
  ANDN U14950 ( .B(n3629), .A(n3630), .Z(n3627) );
  AND U14951 ( .A(a[13]), .B(b[109]), .Z(n3626) );
  XNOR U14952 ( .A(n3631), .B(n2904), .Z(n2906) );
  XOR U14953 ( .A(n3632), .B(n3633), .Z(n2904) );
  ANDN U14954 ( .B(n3634), .A(n3635), .Z(n3632) );
  AND U14955 ( .A(a[14]), .B(b[108]), .Z(n3631) );
  XNOR U14956 ( .A(n3636), .B(n2909), .Z(n2911) );
  XOR U14957 ( .A(n3637), .B(n3638), .Z(n2909) );
  ANDN U14958 ( .B(n3639), .A(n3640), .Z(n3637) );
  AND U14959 ( .A(a[15]), .B(b[107]), .Z(n3636) );
  XNOR U14960 ( .A(n3641), .B(n2914), .Z(n2916) );
  XOR U14961 ( .A(n3642), .B(n3643), .Z(n2914) );
  ANDN U14962 ( .B(n3644), .A(n3645), .Z(n3642) );
  AND U14963 ( .A(a[16]), .B(b[106]), .Z(n3641) );
  XNOR U14964 ( .A(n3646), .B(n2919), .Z(n2921) );
  XOR U14965 ( .A(n3647), .B(n3648), .Z(n2919) );
  ANDN U14966 ( .B(n3649), .A(n3650), .Z(n3647) );
  AND U14967 ( .A(a[17]), .B(b[105]), .Z(n3646) );
  XNOR U14968 ( .A(n3651), .B(n2924), .Z(n2926) );
  XOR U14969 ( .A(n3652), .B(n3653), .Z(n2924) );
  ANDN U14970 ( .B(n3654), .A(n3655), .Z(n3652) );
  AND U14971 ( .A(a[18]), .B(b[104]), .Z(n3651) );
  XNOR U14972 ( .A(n3656), .B(n2929), .Z(n2931) );
  XOR U14973 ( .A(n3657), .B(n3658), .Z(n2929) );
  ANDN U14974 ( .B(n3659), .A(n3660), .Z(n3657) );
  AND U14975 ( .A(a[19]), .B(b[103]), .Z(n3656) );
  XNOR U14976 ( .A(n3661), .B(n2934), .Z(n2936) );
  XOR U14977 ( .A(n3662), .B(n3663), .Z(n2934) );
  ANDN U14978 ( .B(n3664), .A(n3665), .Z(n3662) );
  AND U14979 ( .A(a[20]), .B(b[102]), .Z(n3661) );
  XNOR U14980 ( .A(n3666), .B(n2939), .Z(n2941) );
  XOR U14981 ( .A(n3667), .B(n3668), .Z(n2939) );
  ANDN U14982 ( .B(n3669), .A(n3670), .Z(n3667) );
  AND U14983 ( .A(a[21]), .B(b[101]), .Z(n3666) );
  XNOR U14984 ( .A(n3671), .B(n2944), .Z(n2946) );
  XOR U14985 ( .A(n3672), .B(n3673), .Z(n2944) );
  ANDN U14986 ( .B(n3674), .A(n3675), .Z(n3672) );
  AND U14987 ( .A(a[22]), .B(b[100]), .Z(n3671) );
  XNOR U14988 ( .A(n3676), .B(n2949), .Z(n2951) );
  XOR U14989 ( .A(n3677), .B(n3678), .Z(n2949) );
  ANDN U14990 ( .B(n3679), .A(n3680), .Z(n3677) );
  AND U14991 ( .A(a[23]), .B(b[99]), .Z(n3676) );
  XNOR U14992 ( .A(n3681), .B(n2954), .Z(n2956) );
  XOR U14993 ( .A(n3682), .B(n3683), .Z(n2954) );
  ANDN U14994 ( .B(n3684), .A(n3685), .Z(n3682) );
  AND U14995 ( .A(a[24]), .B(b[98]), .Z(n3681) );
  XNOR U14996 ( .A(n3686), .B(n2959), .Z(n2961) );
  XOR U14997 ( .A(n3687), .B(n3688), .Z(n2959) );
  ANDN U14998 ( .B(n3689), .A(n3690), .Z(n3687) );
  AND U14999 ( .A(a[25]), .B(b[97]), .Z(n3686) );
  XNOR U15000 ( .A(n3691), .B(n2964), .Z(n2966) );
  XOR U15001 ( .A(n3692), .B(n3693), .Z(n2964) );
  ANDN U15002 ( .B(n3694), .A(n3695), .Z(n3692) );
  AND U15003 ( .A(a[26]), .B(b[96]), .Z(n3691) );
  XNOR U15004 ( .A(n3696), .B(n2969), .Z(n2971) );
  XOR U15005 ( .A(n3697), .B(n3698), .Z(n2969) );
  ANDN U15006 ( .B(n3699), .A(n3700), .Z(n3697) );
  AND U15007 ( .A(a[27]), .B(b[95]), .Z(n3696) );
  XNOR U15008 ( .A(n3701), .B(n2974), .Z(n2976) );
  XOR U15009 ( .A(n3702), .B(n3703), .Z(n2974) );
  ANDN U15010 ( .B(n3704), .A(n3705), .Z(n3702) );
  AND U15011 ( .A(a[28]), .B(b[94]), .Z(n3701) );
  XNOR U15012 ( .A(n3706), .B(n2979), .Z(n2981) );
  XOR U15013 ( .A(n3707), .B(n3708), .Z(n2979) );
  ANDN U15014 ( .B(n3709), .A(n3710), .Z(n3707) );
  AND U15015 ( .A(a[29]), .B(b[93]), .Z(n3706) );
  XNOR U15016 ( .A(n3711), .B(n2984), .Z(n2986) );
  XOR U15017 ( .A(n3712), .B(n3713), .Z(n2984) );
  ANDN U15018 ( .B(n3714), .A(n3715), .Z(n3712) );
  AND U15019 ( .A(a[30]), .B(b[92]), .Z(n3711) );
  XNOR U15020 ( .A(n3716), .B(n2989), .Z(n2991) );
  XOR U15021 ( .A(n3717), .B(n3718), .Z(n2989) );
  ANDN U15022 ( .B(n3719), .A(n3720), .Z(n3717) );
  AND U15023 ( .A(a[31]), .B(b[91]), .Z(n3716) );
  XNOR U15024 ( .A(n3721), .B(n2994), .Z(n2996) );
  XOR U15025 ( .A(n3722), .B(n3723), .Z(n2994) );
  ANDN U15026 ( .B(n3724), .A(n3725), .Z(n3722) );
  AND U15027 ( .A(a[32]), .B(b[90]), .Z(n3721) );
  XNOR U15028 ( .A(n3726), .B(n2999), .Z(n3001) );
  XOR U15029 ( .A(n3727), .B(n3728), .Z(n2999) );
  ANDN U15030 ( .B(n3729), .A(n3730), .Z(n3727) );
  AND U15031 ( .A(a[33]), .B(b[89]), .Z(n3726) );
  XNOR U15032 ( .A(n3731), .B(n3004), .Z(n3006) );
  XOR U15033 ( .A(n3732), .B(n3733), .Z(n3004) );
  ANDN U15034 ( .B(n3734), .A(n3735), .Z(n3732) );
  AND U15035 ( .A(a[34]), .B(b[88]), .Z(n3731) );
  XNOR U15036 ( .A(n3736), .B(n3009), .Z(n3011) );
  XOR U15037 ( .A(n3737), .B(n3738), .Z(n3009) );
  ANDN U15038 ( .B(n3739), .A(n3740), .Z(n3737) );
  AND U15039 ( .A(a[35]), .B(b[87]), .Z(n3736) );
  XNOR U15040 ( .A(n3741), .B(n3014), .Z(n3016) );
  XOR U15041 ( .A(n3742), .B(n3743), .Z(n3014) );
  ANDN U15042 ( .B(n3744), .A(n3745), .Z(n3742) );
  AND U15043 ( .A(a[36]), .B(b[86]), .Z(n3741) );
  XNOR U15044 ( .A(n3746), .B(n3019), .Z(n3021) );
  XOR U15045 ( .A(n3747), .B(n3748), .Z(n3019) );
  ANDN U15046 ( .B(n3749), .A(n3750), .Z(n3747) );
  AND U15047 ( .A(a[37]), .B(b[85]), .Z(n3746) );
  XNOR U15048 ( .A(n3751), .B(n3024), .Z(n3026) );
  XOR U15049 ( .A(n3752), .B(n3753), .Z(n3024) );
  ANDN U15050 ( .B(n3754), .A(n3755), .Z(n3752) );
  AND U15051 ( .A(a[38]), .B(b[84]), .Z(n3751) );
  XNOR U15052 ( .A(n3756), .B(n3029), .Z(n3031) );
  XOR U15053 ( .A(n3757), .B(n3758), .Z(n3029) );
  ANDN U15054 ( .B(n3759), .A(n3760), .Z(n3757) );
  AND U15055 ( .A(a[39]), .B(b[83]), .Z(n3756) );
  XNOR U15056 ( .A(n3761), .B(n3034), .Z(n3036) );
  XOR U15057 ( .A(n3762), .B(n3763), .Z(n3034) );
  ANDN U15058 ( .B(n3764), .A(n3765), .Z(n3762) );
  AND U15059 ( .A(a[40]), .B(b[82]), .Z(n3761) );
  XNOR U15060 ( .A(n3766), .B(n3039), .Z(n3041) );
  XOR U15061 ( .A(n3767), .B(n3768), .Z(n3039) );
  ANDN U15062 ( .B(n3769), .A(n3770), .Z(n3767) );
  AND U15063 ( .A(a[41]), .B(b[81]), .Z(n3766) );
  XNOR U15064 ( .A(n3771), .B(n3044), .Z(n3046) );
  XOR U15065 ( .A(n3772), .B(n3773), .Z(n3044) );
  ANDN U15066 ( .B(n3774), .A(n3775), .Z(n3772) );
  AND U15067 ( .A(a[42]), .B(b[80]), .Z(n3771) );
  XNOR U15068 ( .A(n3776), .B(n3049), .Z(n3051) );
  XOR U15069 ( .A(n3777), .B(n3778), .Z(n3049) );
  ANDN U15070 ( .B(n3779), .A(n3780), .Z(n3777) );
  AND U15071 ( .A(a[43]), .B(b[79]), .Z(n3776) );
  XNOR U15072 ( .A(n3781), .B(n3054), .Z(n3056) );
  XOR U15073 ( .A(n3782), .B(n3783), .Z(n3054) );
  ANDN U15074 ( .B(n3784), .A(n3785), .Z(n3782) );
  AND U15075 ( .A(a[44]), .B(b[78]), .Z(n3781) );
  XNOR U15076 ( .A(n3786), .B(n3059), .Z(n3061) );
  XOR U15077 ( .A(n3787), .B(n3788), .Z(n3059) );
  ANDN U15078 ( .B(n3789), .A(n3790), .Z(n3787) );
  AND U15079 ( .A(a[45]), .B(b[77]), .Z(n3786) );
  XNOR U15080 ( .A(n3791), .B(n3064), .Z(n3066) );
  XOR U15081 ( .A(n3792), .B(n3793), .Z(n3064) );
  ANDN U15082 ( .B(n3794), .A(n3795), .Z(n3792) );
  AND U15083 ( .A(a[46]), .B(b[76]), .Z(n3791) );
  XNOR U15084 ( .A(n3796), .B(n3069), .Z(n3071) );
  XOR U15085 ( .A(n3797), .B(n3798), .Z(n3069) );
  ANDN U15086 ( .B(n3799), .A(n3800), .Z(n3797) );
  AND U15087 ( .A(a[47]), .B(b[75]), .Z(n3796) );
  XNOR U15088 ( .A(n3801), .B(n3074), .Z(n3076) );
  XOR U15089 ( .A(n3802), .B(n3803), .Z(n3074) );
  ANDN U15090 ( .B(n3804), .A(n3805), .Z(n3802) );
  AND U15091 ( .A(a[48]), .B(b[74]), .Z(n3801) );
  XNOR U15092 ( .A(n3806), .B(n3079), .Z(n3081) );
  XOR U15093 ( .A(n3807), .B(n3808), .Z(n3079) );
  ANDN U15094 ( .B(n3809), .A(n3810), .Z(n3807) );
  AND U15095 ( .A(a[49]), .B(b[73]), .Z(n3806) );
  XNOR U15096 ( .A(n3811), .B(n3084), .Z(n3086) );
  XOR U15097 ( .A(n3812), .B(n3813), .Z(n3084) );
  ANDN U15098 ( .B(n3814), .A(n3815), .Z(n3812) );
  AND U15099 ( .A(a[50]), .B(b[72]), .Z(n3811) );
  XNOR U15100 ( .A(n3816), .B(n3089), .Z(n3091) );
  XOR U15101 ( .A(n3817), .B(n3818), .Z(n3089) );
  ANDN U15102 ( .B(n3819), .A(n3820), .Z(n3817) );
  AND U15103 ( .A(a[51]), .B(b[71]), .Z(n3816) );
  XNOR U15104 ( .A(n3821), .B(n3094), .Z(n3096) );
  XOR U15105 ( .A(n3822), .B(n3823), .Z(n3094) );
  ANDN U15106 ( .B(n3824), .A(n3825), .Z(n3822) );
  AND U15107 ( .A(a[52]), .B(b[70]), .Z(n3821) );
  XNOR U15108 ( .A(n3826), .B(n3099), .Z(n3101) );
  XOR U15109 ( .A(n3827), .B(n3828), .Z(n3099) );
  ANDN U15110 ( .B(n3829), .A(n3830), .Z(n3827) );
  AND U15111 ( .A(a[53]), .B(b[69]), .Z(n3826) );
  XNOR U15112 ( .A(n3831), .B(n3104), .Z(n3106) );
  XOR U15113 ( .A(n3832), .B(n3833), .Z(n3104) );
  ANDN U15114 ( .B(n3834), .A(n3835), .Z(n3832) );
  AND U15115 ( .A(a[54]), .B(b[68]), .Z(n3831) );
  XNOR U15116 ( .A(n3836), .B(n3109), .Z(n3111) );
  XOR U15117 ( .A(n3837), .B(n3838), .Z(n3109) );
  ANDN U15118 ( .B(n3839), .A(n3840), .Z(n3837) );
  AND U15119 ( .A(a[55]), .B(b[67]), .Z(n3836) );
  XNOR U15120 ( .A(n3841), .B(n3114), .Z(n3116) );
  XOR U15121 ( .A(n3842), .B(n3843), .Z(n3114) );
  ANDN U15122 ( .B(n3844), .A(n3845), .Z(n3842) );
  AND U15123 ( .A(a[56]), .B(b[66]), .Z(n3841) );
  XNOR U15124 ( .A(n3846), .B(n3119), .Z(n3121) );
  XOR U15125 ( .A(n3847), .B(n3848), .Z(n3119) );
  ANDN U15126 ( .B(n3849), .A(n3850), .Z(n3847) );
  AND U15127 ( .A(a[57]), .B(b[65]), .Z(n3846) );
  XNOR U15128 ( .A(n3851), .B(n3124), .Z(n3126) );
  XOR U15129 ( .A(n3852), .B(n3853), .Z(n3124) );
  ANDN U15130 ( .B(n3854), .A(n3855), .Z(n3852) );
  AND U15131 ( .A(a[58]), .B(b[64]), .Z(n3851) );
  XNOR U15132 ( .A(n3856), .B(n3129), .Z(n3131) );
  XOR U15133 ( .A(n3857), .B(n3858), .Z(n3129) );
  ANDN U15134 ( .B(n3859), .A(n3860), .Z(n3857) );
  AND U15135 ( .A(a[59]), .B(b[63]), .Z(n3856) );
  XNOR U15136 ( .A(n3861), .B(n3134), .Z(n3136) );
  XOR U15137 ( .A(n3862), .B(n3863), .Z(n3134) );
  ANDN U15138 ( .B(n3864), .A(n3865), .Z(n3862) );
  AND U15139 ( .A(a[60]), .B(b[62]), .Z(n3861) );
  XNOR U15140 ( .A(n3866), .B(n3139), .Z(n3141) );
  XOR U15141 ( .A(n3867), .B(n3868), .Z(n3139) );
  ANDN U15142 ( .B(n3869), .A(n3870), .Z(n3867) );
  AND U15143 ( .A(a[61]), .B(b[61]), .Z(n3866) );
  XNOR U15144 ( .A(n3871), .B(n3144), .Z(n3146) );
  XOR U15145 ( .A(n3872), .B(n3873), .Z(n3144) );
  ANDN U15146 ( .B(n3874), .A(n3875), .Z(n3872) );
  AND U15147 ( .A(a[62]), .B(b[60]), .Z(n3871) );
  XNOR U15148 ( .A(n3876), .B(n3149), .Z(n3151) );
  XOR U15149 ( .A(n3877), .B(n3878), .Z(n3149) );
  ANDN U15150 ( .B(n3879), .A(n3880), .Z(n3877) );
  AND U15151 ( .A(a[63]), .B(b[59]), .Z(n3876) );
  XNOR U15152 ( .A(n3881), .B(n3154), .Z(n3156) );
  XOR U15153 ( .A(n3882), .B(n3883), .Z(n3154) );
  ANDN U15154 ( .B(n3884), .A(n3885), .Z(n3882) );
  AND U15155 ( .A(a[64]), .B(b[58]), .Z(n3881) );
  XNOR U15156 ( .A(n3886), .B(n3159), .Z(n3161) );
  XOR U15157 ( .A(n3887), .B(n3888), .Z(n3159) );
  ANDN U15158 ( .B(n3889), .A(n3890), .Z(n3887) );
  AND U15159 ( .A(a[65]), .B(b[57]), .Z(n3886) );
  XNOR U15160 ( .A(n3891), .B(n3164), .Z(n3166) );
  XOR U15161 ( .A(n3892), .B(n3893), .Z(n3164) );
  ANDN U15162 ( .B(n3894), .A(n3895), .Z(n3892) );
  AND U15163 ( .A(a[66]), .B(b[56]), .Z(n3891) );
  XNOR U15164 ( .A(n3896), .B(n3169), .Z(n3171) );
  XOR U15165 ( .A(n3897), .B(n3898), .Z(n3169) );
  ANDN U15166 ( .B(n3899), .A(n3900), .Z(n3897) );
  AND U15167 ( .A(a[67]), .B(b[55]), .Z(n3896) );
  XNOR U15168 ( .A(n3901), .B(n3174), .Z(n3176) );
  XOR U15169 ( .A(n3902), .B(n3903), .Z(n3174) );
  ANDN U15170 ( .B(n3904), .A(n3905), .Z(n3902) );
  AND U15171 ( .A(a[68]), .B(b[54]), .Z(n3901) );
  XNOR U15172 ( .A(n3906), .B(n3179), .Z(n3181) );
  XOR U15173 ( .A(n3907), .B(n3908), .Z(n3179) );
  ANDN U15174 ( .B(n3909), .A(n3910), .Z(n3907) );
  AND U15175 ( .A(a[69]), .B(b[53]), .Z(n3906) );
  XNOR U15176 ( .A(n3911), .B(n3184), .Z(n3186) );
  XOR U15177 ( .A(n3912), .B(n3913), .Z(n3184) );
  ANDN U15178 ( .B(n3914), .A(n3915), .Z(n3912) );
  AND U15179 ( .A(a[70]), .B(b[52]), .Z(n3911) );
  XNOR U15180 ( .A(n3916), .B(n3189), .Z(n3191) );
  XOR U15181 ( .A(n3917), .B(n3918), .Z(n3189) );
  ANDN U15182 ( .B(n3919), .A(n3920), .Z(n3917) );
  AND U15183 ( .A(a[71]), .B(b[51]), .Z(n3916) );
  XNOR U15184 ( .A(n3921), .B(n3194), .Z(n3196) );
  XOR U15185 ( .A(n3922), .B(n3923), .Z(n3194) );
  ANDN U15186 ( .B(n3924), .A(n3925), .Z(n3922) );
  AND U15187 ( .A(a[72]), .B(b[50]), .Z(n3921) );
  XNOR U15188 ( .A(n3926), .B(n3199), .Z(n3201) );
  XOR U15189 ( .A(n3927), .B(n3928), .Z(n3199) );
  ANDN U15190 ( .B(n3929), .A(n3930), .Z(n3927) );
  AND U15191 ( .A(a[73]), .B(b[49]), .Z(n3926) );
  XNOR U15192 ( .A(n3931), .B(n3204), .Z(n3206) );
  XOR U15193 ( .A(n3932), .B(n3933), .Z(n3204) );
  ANDN U15194 ( .B(n3934), .A(n3935), .Z(n3932) );
  AND U15195 ( .A(a[74]), .B(b[48]), .Z(n3931) );
  XNOR U15196 ( .A(n3936), .B(n3209), .Z(n3211) );
  XOR U15197 ( .A(n3937), .B(n3938), .Z(n3209) );
  ANDN U15198 ( .B(n3939), .A(n3940), .Z(n3937) );
  AND U15199 ( .A(a[75]), .B(b[47]), .Z(n3936) );
  XNOR U15200 ( .A(n3941), .B(n3214), .Z(n3216) );
  XOR U15201 ( .A(n3942), .B(n3943), .Z(n3214) );
  ANDN U15202 ( .B(n3944), .A(n3945), .Z(n3942) );
  AND U15203 ( .A(a[76]), .B(b[46]), .Z(n3941) );
  XNOR U15204 ( .A(n3946), .B(n3219), .Z(n3221) );
  XOR U15205 ( .A(n3947), .B(n3948), .Z(n3219) );
  ANDN U15206 ( .B(n3949), .A(n3950), .Z(n3947) );
  AND U15207 ( .A(a[77]), .B(b[45]), .Z(n3946) );
  XNOR U15208 ( .A(n3951), .B(n3224), .Z(n3226) );
  XOR U15209 ( .A(n3952), .B(n3953), .Z(n3224) );
  ANDN U15210 ( .B(n3954), .A(n3955), .Z(n3952) );
  AND U15211 ( .A(a[78]), .B(b[44]), .Z(n3951) );
  XNOR U15212 ( .A(n3956), .B(n3229), .Z(n3231) );
  XOR U15213 ( .A(n3957), .B(n3958), .Z(n3229) );
  ANDN U15214 ( .B(n3959), .A(n3960), .Z(n3957) );
  AND U15215 ( .A(a[79]), .B(b[43]), .Z(n3956) );
  XNOR U15216 ( .A(n3961), .B(n3234), .Z(n3236) );
  XOR U15217 ( .A(n3962), .B(n3963), .Z(n3234) );
  ANDN U15218 ( .B(n3964), .A(n3965), .Z(n3962) );
  AND U15219 ( .A(a[80]), .B(b[42]), .Z(n3961) );
  XNOR U15220 ( .A(n3966), .B(n3239), .Z(n3241) );
  XOR U15221 ( .A(n3967), .B(n3968), .Z(n3239) );
  ANDN U15222 ( .B(n3969), .A(n3970), .Z(n3967) );
  AND U15223 ( .A(a[81]), .B(b[41]), .Z(n3966) );
  XNOR U15224 ( .A(n3971), .B(n3244), .Z(n3246) );
  XOR U15225 ( .A(n3972), .B(n3973), .Z(n3244) );
  ANDN U15226 ( .B(n3974), .A(n3975), .Z(n3972) );
  AND U15227 ( .A(a[82]), .B(b[40]), .Z(n3971) );
  XNOR U15228 ( .A(n3976), .B(n3249), .Z(n3251) );
  XOR U15229 ( .A(n3977), .B(n3978), .Z(n3249) );
  ANDN U15230 ( .B(n3979), .A(n3980), .Z(n3977) );
  AND U15231 ( .A(a[83]), .B(b[39]), .Z(n3976) );
  XNOR U15232 ( .A(n3981), .B(n3254), .Z(n3256) );
  XOR U15233 ( .A(n3982), .B(n3983), .Z(n3254) );
  ANDN U15234 ( .B(n3984), .A(n3985), .Z(n3982) );
  AND U15235 ( .A(a[84]), .B(b[38]), .Z(n3981) );
  XNOR U15236 ( .A(n3986), .B(n3259), .Z(n3261) );
  XOR U15237 ( .A(n3987), .B(n3988), .Z(n3259) );
  ANDN U15238 ( .B(n3989), .A(n3990), .Z(n3987) );
  AND U15239 ( .A(a[85]), .B(b[37]), .Z(n3986) );
  XNOR U15240 ( .A(n3991), .B(n3264), .Z(n3266) );
  XOR U15241 ( .A(n3992), .B(n3993), .Z(n3264) );
  ANDN U15242 ( .B(n3994), .A(n3995), .Z(n3992) );
  AND U15243 ( .A(a[86]), .B(b[36]), .Z(n3991) );
  XNOR U15244 ( .A(n3996), .B(n3269), .Z(n3271) );
  XOR U15245 ( .A(n3997), .B(n3998), .Z(n3269) );
  ANDN U15246 ( .B(n3999), .A(n4000), .Z(n3997) );
  AND U15247 ( .A(a[87]), .B(b[35]), .Z(n3996) );
  XNOR U15248 ( .A(n4001), .B(n3274), .Z(n3276) );
  XOR U15249 ( .A(n4002), .B(n4003), .Z(n3274) );
  ANDN U15250 ( .B(n4004), .A(n4005), .Z(n4002) );
  AND U15251 ( .A(a[88]), .B(b[34]), .Z(n4001) );
  XNOR U15252 ( .A(n4006), .B(n3279), .Z(n3281) );
  XOR U15253 ( .A(n4007), .B(n4008), .Z(n3279) );
  ANDN U15254 ( .B(n4009), .A(n4010), .Z(n4007) );
  AND U15255 ( .A(a[89]), .B(b[33]), .Z(n4006) );
  XNOR U15256 ( .A(n4011), .B(n3284), .Z(n3286) );
  XOR U15257 ( .A(n4012), .B(n4013), .Z(n3284) );
  ANDN U15258 ( .B(n4014), .A(n4015), .Z(n4012) );
  AND U15259 ( .A(a[90]), .B(b[32]), .Z(n4011) );
  XNOR U15260 ( .A(n4016), .B(n3289), .Z(n3291) );
  XOR U15261 ( .A(n4017), .B(n4018), .Z(n3289) );
  ANDN U15262 ( .B(n4019), .A(n4020), .Z(n4017) );
  AND U15263 ( .A(a[91]), .B(b[31]), .Z(n4016) );
  XNOR U15264 ( .A(n4021), .B(n3294), .Z(n3296) );
  XOR U15265 ( .A(n4022), .B(n4023), .Z(n3294) );
  ANDN U15266 ( .B(n4024), .A(n4025), .Z(n4022) );
  AND U15267 ( .A(a[92]), .B(b[30]), .Z(n4021) );
  XNOR U15268 ( .A(n4026), .B(n3299), .Z(n3301) );
  XOR U15269 ( .A(n4027), .B(n4028), .Z(n3299) );
  ANDN U15270 ( .B(n4029), .A(n4030), .Z(n4027) );
  AND U15271 ( .A(a[93]), .B(b[29]), .Z(n4026) );
  XNOR U15272 ( .A(n4031), .B(n3304), .Z(n3306) );
  XOR U15273 ( .A(n4032), .B(n4033), .Z(n3304) );
  ANDN U15274 ( .B(n4034), .A(n4035), .Z(n4032) );
  AND U15275 ( .A(a[94]), .B(b[28]), .Z(n4031) );
  XNOR U15276 ( .A(n4036), .B(n3309), .Z(n3311) );
  XOR U15277 ( .A(n4037), .B(n4038), .Z(n3309) );
  ANDN U15278 ( .B(n4039), .A(n4040), .Z(n4037) );
  AND U15279 ( .A(a[95]), .B(b[27]), .Z(n4036) );
  XNOR U15280 ( .A(n4041), .B(n3314), .Z(n3316) );
  XOR U15281 ( .A(n4042), .B(n4043), .Z(n3314) );
  ANDN U15282 ( .B(n4044), .A(n4045), .Z(n4042) );
  AND U15283 ( .A(a[96]), .B(b[26]), .Z(n4041) );
  XNOR U15284 ( .A(n4046), .B(n3319), .Z(n3321) );
  XOR U15285 ( .A(n4047), .B(n4048), .Z(n3319) );
  ANDN U15286 ( .B(n4049), .A(n4050), .Z(n4047) );
  AND U15287 ( .A(a[97]), .B(b[25]), .Z(n4046) );
  XNOR U15288 ( .A(n4051), .B(n3324), .Z(n3326) );
  XOR U15289 ( .A(n4052), .B(n4053), .Z(n3324) );
  ANDN U15290 ( .B(n4054), .A(n4055), .Z(n4052) );
  AND U15291 ( .A(a[98]), .B(b[24]), .Z(n4051) );
  XNOR U15292 ( .A(n4056), .B(n3329), .Z(n3331) );
  XOR U15293 ( .A(n4057), .B(n4058), .Z(n3329) );
  ANDN U15294 ( .B(n4059), .A(n4060), .Z(n4057) );
  AND U15295 ( .A(a[99]), .B(b[23]), .Z(n4056) );
  XNOR U15296 ( .A(n4061), .B(n3334), .Z(n3336) );
  XOR U15297 ( .A(n4062), .B(n4063), .Z(n3334) );
  ANDN U15298 ( .B(n4064), .A(n4065), .Z(n4062) );
  AND U15299 ( .A(b[22]), .B(a[100]), .Z(n4061) );
  XNOR U15300 ( .A(n4066), .B(n3339), .Z(n3341) );
  XOR U15301 ( .A(n4067), .B(n4068), .Z(n3339) );
  ANDN U15302 ( .B(n4069), .A(n4070), .Z(n4067) );
  AND U15303 ( .A(b[21]), .B(a[101]), .Z(n4066) );
  XNOR U15304 ( .A(n4071), .B(n3344), .Z(n3346) );
  XOR U15305 ( .A(n4072), .B(n4073), .Z(n3344) );
  ANDN U15306 ( .B(n4074), .A(n4075), .Z(n4072) );
  AND U15307 ( .A(b[20]), .B(a[102]), .Z(n4071) );
  XNOR U15308 ( .A(n4076), .B(n3349), .Z(n3351) );
  XOR U15309 ( .A(n4077), .B(n4078), .Z(n3349) );
  ANDN U15310 ( .B(n4079), .A(n4080), .Z(n4077) );
  AND U15311 ( .A(b[19]), .B(a[103]), .Z(n4076) );
  XNOR U15312 ( .A(n4081), .B(n3354), .Z(n3356) );
  XOR U15313 ( .A(n4082), .B(n4083), .Z(n3354) );
  ANDN U15314 ( .B(n4084), .A(n4085), .Z(n4082) );
  AND U15315 ( .A(b[18]), .B(a[104]), .Z(n4081) );
  XNOR U15316 ( .A(n4086), .B(n3359), .Z(n3361) );
  XOR U15317 ( .A(n4087), .B(n4088), .Z(n3359) );
  ANDN U15318 ( .B(n4089), .A(n4090), .Z(n4087) );
  AND U15319 ( .A(b[17]), .B(a[105]), .Z(n4086) );
  XNOR U15320 ( .A(n4091), .B(n3364), .Z(n3366) );
  XOR U15321 ( .A(n4092), .B(n4093), .Z(n3364) );
  ANDN U15322 ( .B(n4094), .A(n4095), .Z(n4092) );
  AND U15323 ( .A(b[16]), .B(a[106]), .Z(n4091) );
  XNOR U15324 ( .A(n4096), .B(n3369), .Z(n3371) );
  XOR U15325 ( .A(n4097), .B(n4098), .Z(n3369) );
  ANDN U15326 ( .B(n4099), .A(n4100), .Z(n4097) );
  AND U15327 ( .A(b[15]), .B(a[107]), .Z(n4096) );
  XNOR U15328 ( .A(n4101), .B(n3374), .Z(n3376) );
  XOR U15329 ( .A(n4102), .B(n4103), .Z(n3374) );
  ANDN U15330 ( .B(n4104), .A(n4105), .Z(n4102) );
  AND U15331 ( .A(b[14]), .B(a[108]), .Z(n4101) );
  XNOR U15332 ( .A(n4106), .B(n3379), .Z(n3381) );
  XOR U15333 ( .A(n4107), .B(n4108), .Z(n3379) );
  ANDN U15334 ( .B(n4109), .A(n4110), .Z(n4107) );
  AND U15335 ( .A(b[13]), .B(a[109]), .Z(n4106) );
  XNOR U15336 ( .A(n4111), .B(n3384), .Z(n3386) );
  XOR U15337 ( .A(n4112), .B(n4113), .Z(n3384) );
  ANDN U15338 ( .B(n4114), .A(n4115), .Z(n4112) );
  AND U15339 ( .A(b[12]), .B(a[110]), .Z(n4111) );
  XNOR U15340 ( .A(n4116), .B(n3389), .Z(n3391) );
  XOR U15341 ( .A(n4117), .B(n4118), .Z(n3389) );
  ANDN U15342 ( .B(n4119), .A(n4120), .Z(n4117) );
  AND U15343 ( .A(b[11]), .B(a[111]), .Z(n4116) );
  XNOR U15344 ( .A(n4121), .B(n3394), .Z(n3396) );
  XOR U15345 ( .A(n4122), .B(n4123), .Z(n3394) );
  ANDN U15346 ( .B(n4124), .A(n4125), .Z(n4122) );
  AND U15347 ( .A(b[10]), .B(a[112]), .Z(n4121) );
  XNOR U15348 ( .A(n4126), .B(n3399), .Z(n3401) );
  XOR U15349 ( .A(n4127), .B(n4128), .Z(n3399) );
  ANDN U15350 ( .B(n4129), .A(n4130), .Z(n4127) );
  AND U15351 ( .A(b[9]), .B(a[113]), .Z(n4126) );
  XNOR U15352 ( .A(n4131), .B(n3404), .Z(n3406) );
  XOR U15353 ( .A(n4132), .B(n4133), .Z(n3404) );
  ANDN U15354 ( .B(n4134), .A(n4135), .Z(n4132) );
  AND U15355 ( .A(b[8]), .B(a[114]), .Z(n4131) );
  XNOR U15356 ( .A(n4136), .B(n3409), .Z(n3411) );
  XOR U15357 ( .A(n4137), .B(n4138), .Z(n3409) );
  ANDN U15358 ( .B(n4139), .A(n4140), .Z(n4137) );
  AND U15359 ( .A(b[7]), .B(a[115]), .Z(n4136) );
  XNOR U15360 ( .A(n4141), .B(n3414), .Z(n3416) );
  XOR U15361 ( .A(n4142), .B(n4143), .Z(n3414) );
  ANDN U15362 ( .B(n4144), .A(n4145), .Z(n4142) );
  AND U15363 ( .A(b[6]), .B(a[116]), .Z(n4141) );
  XNOR U15364 ( .A(n4146), .B(n3419), .Z(n3421) );
  XOR U15365 ( .A(n4147), .B(n4148), .Z(n3419) );
  ANDN U15366 ( .B(n4149), .A(n4150), .Z(n4147) );
  AND U15367 ( .A(b[5]), .B(a[117]), .Z(n4146) );
  XNOR U15368 ( .A(n4151), .B(n3424), .Z(n3426) );
  XOR U15369 ( .A(n4152), .B(n4153), .Z(n3424) );
  ANDN U15370 ( .B(n4154), .A(n4155), .Z(n4152) );
  AND U15371 ( .A(b[4]), .B(a[118]), .Z(n4151) );
  XNOR U15372 ( .A(n4156), .B(n4157), .Z(n3438) );
  NANDN U15373 ( .A(n4158), .B(n4159), .Z(n4157) );
  XNOR U15374 ( .A(n4160), .B(n3429), .Z(n3431) );
  XNOR U15375 ( .A(n4161), .B(n4162), .Z(n3429) );
  AND U15376 ( .A(n4163), .B(n4164), .Z(n4161) );
  AND U15377 ( .A(b[3]), .B(a[119]), .Z(n4160) );
  NAND U15378 ( .A(a[122]), .B(b[0]), .Z(n2714) );
  XNOR U15379 ( .A(n3444), .B(n3445), .Z(c[121]) );
  XNOR U15380 ( .A(n4158), .B(n4159), .Z(n3445) );
  XOR U15381 ( .A(n4156), .B(n4165), .Z(n4159) );
  NAND U15382 ( .A(b[1]), .B(a[120]), .Z(n4165) );
  XOR U15383 ( .A(n4164), .B(n4166), .Z(n4158) );
  XOR U15384 ( .A(n4156), .B(n4163), .Z(n4166) );
  XNOR U15385 ( .A(n4167), .B(n4162), .Z(n4163) );
  AND U15386 ( .A(b[2]), .B(a[119]), .Z(n4167) );
  NANDN U15387 ( .A(n4168), .B(n4169), .Z(n4156) );
  XOR U15388 ( .A(n4162), .B(n4154), .Z(n4170) );
  XNOR U15389 ( .A(n4153), .B(n4149), .Z(n4171) );
  XNOR U15390 ( .A(n4148), .B(n4144), .Z(n4172) );
  XNOR U15391 ( .A(n4143), .B(n4139), .Z(n4173) );
  XNOR U15392 ( .A(n4138), .B(n4134), .Z(n4174) );
  XNOR U15393 ( .A(n4133), .B(n4129), .Z(n4175) );
  XNOR U15394 ( .A(n4128), .B(n4124), .Z(n4176) );
  XNOR U15395 ( .A(n4123), .B(n4119), .Z(n4177) );
  XNOR U15396 ( .A(n4118), .B(n4114), .Z(n4178) );
  XNOR U15397 ( .A(n4113), .B(n4109), .Z(n4179) );
  XNOR U15398 ( .A(n4108), .B(n4104), .Z(n4180) );
  XNOR U15399 ( .A(n4103), .B(n4099), .Z(n4181) );
  XNOR U15400 ( .A(n4098), .B(n4094), .Z(n4182) );
  XNOR U15401 ( .A(n4093), .B(n4089), .Z(n4183) );
  XNOR U15402 ( .A(n4088), .B(n4084), .Z(n4184) );
  XNOR U15403 ( .A(n4083), .B(n4079), .Z(n4185) );
  XNOR U15404 ( .A(n4078), .B(n4074), .Z(n4186) );
  XNOR U15405 ( .A(n4073), .B(n4069), .Z(n4187) );
  XNOR U15406 ( .A(n4068), .B(n4064), .Z(n4188) );
  XNOR U15407 ( .A(n4063), .B(n4059), .Z(n4189) );
  XNOR U15408 ( .A(n4058), .B(n4054), .Z(n4190) );
  XNOR U15409 ( .A(n4053), .B(n4049), .Z(n4191) );
  XNOR U15410 ( .A(n4048), .B(n4044), .Z(n4192) );
  XNOR U15411 ( .A(n4043), .B(n4039), .Z(n4193) );
  XNOR U15412 ( .A(n4038), .B(n4034), .Z(n4194) );
  XNOR U15413 ( .A(n4033), .B(n4029), .Z(n4195) );
  XNOR U15414 ( .A(n4028), .B(n4024), .Z(n4196) );
  XNOR U15415 ( .A(n4023), .B(n4019), .Z(n4197) );
  XNOR U15416 ( .A(n4018), .B(n4014), .Z(n4198) );
  XNOR U15417 ( .A(n4013), .B(n4009), .Z(n4199) );
  XNOR U15418 ( .A(n4008), .B(n4004), .Z(n4200) );
  XNOR U15419 ( .A(n4003), .B(n3999), .Z(n4201) );
  XNOR U15420 ( .A(n3998), .B(n3994), .Z(n4202) );
  XNOR U15421 ( .A(n3993), .B(n3989), .Z(n4203) );
  XNOR U15422 ( .A(n3988), .B(n3984), .Z(n4204) );
  XNOR U15423 ( .A(n3983), .B(n3979), .Z(n4205) );
  XNOR U15424 ( .A(n3978), .B(n3974), .Z(n4206) );
  XNOR U15425 ( .A(n3973), .B(n3969), .Z(n4207) );
  XNOR U15426 ( .A(n3968), .B(n3964), .Z(n4208) );
  XNOR U15427 ( .A(n3963), .B(n3959), .Z(n4209) );
  XNOR U15428 ( .A(n3958), .B(n3954), .Z(n4210) );
  XNOR U15429 ( .A(n3953), .B(n3949), .Z(n4211) );
  XNOR U15430 ( .A(n3948), .B(n3944), .Z(n4212) );
  XNOR U15431 ( .A(n3943), .B(n3939), .Z(n4213) );
  XNOR U15432 ( .A(n3938), .B(n3934), .Z(n4214) );
  XNOR U15433 ( .A(n3933), .B(n3929), .Z(n4215) );
  XNOR U15434 ( .A(n3928), .B(n3924), .Z(n4216) );
  XNOR U15435 ( .A(n3923), .B(n3919), .Z(n4217) );
  XNOR U15436 ( .A(n3918), .B(n3914), .Z(n4218) );
  XNOR U15437 ( .A(n3913), .B(n3909), .Z(n4219) );
  XNOR U15438 ( .A(n3908), .B(n3904), .Z(n4220) );
  XNOR U15439 ( .A(n3903), .B(n3899), .Z(n4221) );
  XNOR U15440 ( .A(n3898), .B(n3894), .Z(n4222) );
  XNOR U15441 ( .A(n3893), .B(n3889), .Z(n4223) );
  XNOR U15442 ( .A(n3888), .B(n3884), .Z(n4224) );
  XNOR U15443 ( .A(n3883), .B(n3879), .Z(n4225) );
  XNOR U15444 ( .A(n3878), .B(n3874), .Z(n4226) );
  XNOR U15445 ( .A(n3873), .B(n3869), .Z(n4227) );
  XNOR U15446 ( .A(n3868), .B(n3864), .Z(n4228) );
  XNOR U15447 ( .A(n3863), .B(n3859), .Z(n4229) );
  XNOR U15448 ( .A(n3858), .B(n3854), .Z(n4230) );
  XNOR U15449 ( .A(n3853), .B(n3849), .Z(n4231) );
  XNOR U15450 ( .A(n3848), .B(n3844), .Z(n4232) );
  XNOR U15451 ( .A(n3843), .B(n3839), .Z(n4233) );
  XNOR U15452 ( .A(n3838), .B(n3834), .Z(n4234) );
  XNOR U15453 ( .A(n3833), .B(n3829), .Z(n4235) );
  XNOR U15454 ( .A(n3828), .B(n3824), .Z(n4236) );
  XNOR U15455 ( .A(n3823), .B(n3819), .Z(n4237) );
  XNOR U15456 ( .A(n3818), .B(n3814), .Z(n4238) );
  XNOR U15457 ( .A(n3813), .B(n3809), .Z(n4239) );
  XNOR U15458 ( .A(n3808), .B(n3804), .Z(n4240) );
  XNOR U15459 ( .A(n3803), .B(n3799), .Z(n4241) );
  XNOR U15460 ( .A(n3798), .B(n3794), .Z(n4242) );
  XNOR U15461 ( .A(n3793), .B(n3789), .Z(n4243) );
  XNOR U15462 ( .A(n3788), .B(n3784), .Z(n4244) );
  XNOR U15463 ( .A(n3783), .B(n3779), .Z(n4245) );
  XNOR U15464 ( .A(n3778), .B(n3774), .Z(n4246) );
  XNOR U15465 ( .A(n3773), .B(n3769), .Z(n4247) );
  XNOR U15466 ( .A(n3768), .B(n3764), .Z(n4248) );
  XNOR U15467 ( .A(n3763), .B(n3759), .Z(n4249) );
  XNOR U15468 ( .A(n3758), .B(n3754), .Z(n4250) );
  XNOR U15469 ( .A(n3753), .B(n3749), .Z(n4251) );
  XNOR U15470 ( .A(n3748), .B(n3744), .Z(n4252) );
  XNOR U15471 ( .A(n3743), .B(n3739), .Z(n4253) );
  XNOR U15472 ( .A(n3738), .B(n3734), .Z(n4254) );
  XNOR U15473 ( .A(n3733), .B(n3729), .Z(n4255) );
  XNOR U15474 ( .A(n3728), .B(n3724), .Z(n4256) );
  XNOR U15475 ( .A(n3723), .B(n3719), .Z(n4257) );
  XNOR U15476 ( .A(n3718), .B(n3714), .Z(n4258) );
  XNOR U15477 ( .A(n3713), .B(n3709), .Z(n4259) );
  XNOR U15478 ( .A(n3708), .B(n3704), .Z(n4260) );
  XNOR U15479 ( .A(n3703), .B(n3699), .Z(n4261) );
  XNOR U15480 ( .A(n3698), .B(n3694), .Z(n4262) );
  XNOR U15481 ( .A(n3693), .B(n3689), .Z(n4263) );
  XNOR U15482 ( .A(n3688), .B(n3684), .Z(n4264) );
  XNOR U15483 ( .A(n3683), .B(n3679), .Z(n4265) );
  XNOR U15484 ( .A(n3678), .B(n3674), .Z(n4266) );
  XNOR U15485 ( .A(n3673), .B(n3669), .Z(n4267) );
  XNOR U15486 ( .A(n3668), .B(n3664), .Z(n4268) );
  XNOR U15487 ( .A(n3663), .B(n3659), .Z(n4269) );
  XNOR U15488 ( .A(n3658), .B(n3654), .Z(n4270) );
  XNOR U15489 ( .A(n3653), .B(n3649), .Z(n4271) );
  XNOR U15490 ( .A(n3648), .B(n3644), .Z(n4272) );
  XNOR U15491 ( .A(n3643), .B(n3639), .Z(n4273) );
  XNOR U15492 ( .A(n3638), .B(n3634), .Z(n4274) );
  XNOR U15493 ( .A(n3633), .B(n3629), .Z(n4275) );
  XNOR U15494 ( .A(n3628), .B(n3624), .Z(n4276) );
  XNOR U15495 ( .A(n3623), .B(n3619), .Z(n4277) );
  XNOR U15496 ( .A(n3618), .B(n3614), .Z(n4278) );
  XNOR U15497 ( .A(n3613), .B(n3609), .Z(n4279) );
  XNOR U15498 ( .A(n3608), .B(n3604), .Z(n4280) );
  XNOR U15499 ( .A(n3603), .B(n3599), .Z(n4281) );
  XNOR U15500 ( .A(n3598), .B(n3594), .Z(n4282) );
  XNOR U15501 ( .A(n3593), .B(n3589), .Z(n4283) );
  XNOR U15502 ( .A(n3588), .B(n3584), .Z(n4284) );
  XNOR U15503 ( .A(n3583), .B(n3579), .Z(n4285) );
  XNOR U15504 ( .A(n3578), .B(n3574), .Z(n4286) );
  XNOR U15505 ( .A(n3573), .B(n3569), .Z(n4287) );
  XNOR U15506 ( .A(n4288), .B(n3568), .Z(n3569) );
  AND U15507 ( .A(a[0]), .B(b[121]), .Z(n4288) );
  XOR U15508 ( .A(n4289), .B(n3568), .Z(n3570) );
  XNOR U15509 ( .A(n4290), .B(n4291), .Z(n3568) );
  ANDN U15510 ( .B(n4292), .A(n4293), .Z(n4290) );
  AND U15511 ( .A(a[1]), .B(b[120]), .Z(n4289) );
  XNOR U15512 ( .A(n4294), .B(n3573), .Z(n3575) );
  XOR U15513 ( .A(n4295), .B(n4296), .Z(n3573) );
  ANDN U15514 ( .B(n4297), .A(n4298), .Z(n4295) );
  AND U15515 ( .A(a[2]), .B(b[119]), .Z(n4294) );
  XNOR U15516 ( .A(n4299), .B(n3578), .Z(n3580) );
  XOR U15517 ( .A(n4300), .B(n4301), .Z(n3578) );
  ANDN U15518 ( .B(n4302), .A(n4303), .Z(n4300) );
  AND U15519 ( .A(a[3]), .B(b[118]), .Z(n4299) );
  XNOR U15520 ( .A(n4304), .B(n3583), .Z(n3585) );
  XOR U15521 ( .A(n4305), .B(n4306), .Z(n3583) );
  ANDN U15522 ( .B(n4307), .A(n4308), .Z(n4305) );
  AND U15523 ( .A(a[4]), .B(b[117]), .Z(n4304) );
  XNOR U15524 ( .A(n4309), .B(n3588), .Z(n3590) );
  XOR U15525 ( .A(n4310), .B(n4311), .Z(n3588) );
  ANDN U15526 ( .B(n4312), .A(n4313), .Z(n4310) );
  AND U15527 ( .A(a[5]), .B(b[116]), .Z(n4309) );
  XNOR U15528 ( .A(n4314), .B(n3593), .Z(n3595) );
  XOR U15529 ( .A(n4315), .B(n4316), .Z(n3593) );
  ANDN U15530 ( .B(n4317), .A(n4318), .Z(n4315) );
  AND U15531 ( .A(a[6]), .B(b[115]), .Z(n4314) );
  XNOR U15532 ( .A(n4319), .B(n3598), .Z(n3600) );
  XOR U15533 ( .A(n4320), .B(n4321), .Z(n3598) );
  ANDN U15534 ( .B(n4322), .A(n4323), .Z(n4320) );
  AND U15535 ( .A(a[7]), .B(b[114]), .Z(n4319) );
  XNOR U15536 ( .A(n4324), .B(n3603), .Z(n3605) );
  XOR U15537 ( .A(n4325), .B(n4326), .Z(n3603) );
  ANDN U15538 ( .B(n4327), .A(n4328), .Z(n4325) );
  AND U15539 ( .A(a[8]), .B(b[113]), .Z(n4324) );
  XNOR U15540 ( .A(n4329), .B(n3608), .Z(n3610) );
  XOR U15541 ( .A(n4330), .B(n4331), .Z(n3608) );
  ANDN U15542 ( .B(n4332), .A(n4333), .Z(n4330) );
  AND U15543 ( .A(a[9]), .B(b[112]), .Z(n4329) );
  XNOR U15544 ( .A(n4334), .B(n3613), .Z(n3615) );
  XOR U15545 ( .A(n4335), .B(n4336), .Z(n3613) );
  ANDN U15546 ( .B(n4337), .A(n4338), .Z(n4335) );
  AND U15547 ( .A(a[10]), .B(b[111]), .Z(n4334) );
  XNOR U15548 ( .A(n4339), .B(n3618), .Z(n3620) );
  XOR U15549 ( .A(n4340), .B(n4341), .Z(n3618) );
  ANDN U15550 ( .B(n4342), .A(n4343), .Z(n4340) );
  AND U15551 ( .A(a[11]), .B(b[110]), .Z(n4339) );
  XNOR U15552 ( .A(n4344), .B(n3623), .Z(n3625) );
  XOR U15553 ( .A(n4345), .B(n4346), .Z(n3623) );
  ANDN U15554 ( .B(n4347), .A(n4348), .Z(n4345) );
  AND U15555 ( .A(a[12]), .B(b[109]), .Z(n4344) );
  XNOR U15556 ( .A(n4349), .B(n3628), .Z(n3630) );
  XOR U15557 ( .A(n4350), .B(n4351), .Z(n3628) );
  ANDN U15558 ( .B(n4352), .A(n4353), .Z(n4350) );
  AND U15559 ( .A(a[13]), .B(b[108]), .Z(n4349) );
  XNOR U15560 ( .A(n4354), .B(n3633), .Z(n3635) );
  XOR U15561 ( .A(n4355), .B(n4356), .Z(n3633) );
  ANDN U15562 ( .B(n4357), .A(n4358), .Z(n4355) );
  AND U15563 ( .A(a[14]), .B(b[107]), .Z(n4354) );
  XNOR U15564 ( .A(n4359), .B(n3638), .Z(n3640) );
  XOR U15565 ( .A(n4360), .B(n4361), .Z(n3638) );
  ANDN U15566 ( .B(n4362), .A(n4363), .Z(n4360) );
  AND U15567 ( .A(a[15]), .B(b[106]), .Z(n4359) );
  XNOR U15568 ( .A(n4364), .B(n3643), .Z(n3645) );
  XOR U15569 ( .A(n4365), .B(n4366), .Z(n3643) );
  ANDN U15570 ( .B(n4367), .A(n4368), .Z(n4365) );
  AND U15571 ( .A(a[16]), .B(b[105]), .Z(n4364) );
  XNOR U15572 ( .A(n4369), .B(n3648), .Z(n3650) );
  XOR U15573 ( .A(n4370), .B(n4371), .Z(n3648) );
  ANDN U15574 ( .B(n4372), .A(n4373), .Z(n4370) );
  AND U15575 ( .A(a[17]), .B(b[104]), .Z(n4369) );
  XNOR U15576 ( .A(n4374), .B(n3653), .Z(n3655) );
  XOR U15577 ( .A(n4375), .B(n4376), .Z(n3653) );
  ANDN U15578 ( .B(n4377), .A(n4378), .Z(n4375) );
  AND U15579 ( .A(a[18]), .B(b[103]), .Z(n4374) );
  XNOR U15580 ( .A(n4379), .B(n3658), .Z(n3660) );
  XOR U15581 ( .A(n4380), .B(n4381), .Z(n3658) );
  ANDN U15582 ( .B(n4382), .A(n4383), .Z(n4380) );
  AND U15583 ( .A(a[19]), .B(b[102]), .Z(n4379) );
  XNOR U15584 ( .A(n4384), .B(n3663), .Z(n3665) );
  XOR U15585 ( .A(n4385), .B(n4386), .Z(n3663) );
  ANDN U15586 ( .B(n4387), .A(n4388), .Z(n4385) );
  AND U15587 ( .A(a[20]), .B(b[101]), .Z(n4384) );
  XNOR U15588 ( .A(n4389), .B(n3668), .Z(n3670) );
  XOR U15589 ( .A(n4390), .B(n4391), .Z(n3668) );
  ANDN U15590 ( .B(n4392), .A(n4393), .Z(n4390) );
  AND U15591 ( .A(a[21]), .B(b[100]), .Z(n4389) );
  XNOR U15592 ( .A(n4394), .B(n3673), .Z(n3675) );
  XOR U15593 ( .A(n4395), .B(n4396), .Z(n3673) );
  ANDN U15594 ( .B(n4397), .A(n4398), .Z(n4395) );
  AND U15595 ( .A(a[22]), .B(b[99]), .Z(n4394) );
  XNOR U15596 ( .A(n4399), .B(n3678), .Z(n3680) );
  XOR U15597 ( .A(n4400), .B(n4401), .Z(n3678) );
  ANDN U15598 ( .B(n4402), .A(n4403), .Z(n4400) );
  AND U15599 ( .A(a[23]), .B(b[98]), .Z(n4399) );
  XNOR U15600 ( .A(n4404), .B(n3683), .Z(n3685) );
  XOR U15601 ( .A(n4405), .B(n4406), .Z(n3683) );
  ANDN U15602 ( .B(n4407), .A(n4408), .Z(n4405) );
  AND U15603 ( .A(a[24]), .B(b[97]), .Z(n4404) );
  XNOR U15604 ( .A(n4409), .B(n3688), .Z(n3690) );
  XOR U15605 ( .A(n4410), .B(n4411), .Z(n3688) );
  ANDN U15606 ( .B(n4412), .A(n4413), .Z(n4410) );
  AND U15607 ( .A(a[25]), .B(b[96]), .Z(n4409) );
  XNOR U15608 ( .A(n4414), .B(n3693), .Z(n3695) );
  XOR U15609 ( .A(n4415), .B(n4416), .Z(n3693) );
  ANDN U15610 ( .B(n4417), .A(n4418), .Z(n4415) );
  AND U15611 ( .A(a[26]), .B(b[95]), .Z(n4414) );
  XNOR U15612 ( .A(n4419), .B(n3698), .Z(n3700) );
  XOR U15613 ( .A(n4420), .B(n4421), .Z(n3698) );
  ANDN U15614 ( .B(n4422), .A(n4423), .Z(n4420) );
  AND U15615 ( .A(a[27]), .B(b[94]), .Z(n4419) );
  XNOR U15616 ( .A(n4424), .B(n3703), .Z(n3705) );
  XOR U15617 ( .A(n4425), .B(n4426), .Z(n3703) );
  ANDN U15618 ( .B(n4427), .A(n4428), .Z(n4425) );
  AND U15619 ( .A(a[28]), .B(b[93]), .Z(n4424) );
  XNOR U15620 ( .A(n4429), .B(n3708), .Z(n3710) );
  XOR U15621 ( .A(n4430), .B(n4431), .Z(n3708) );
  ANDN U15622 ( .B(n4432), .A(n4433), .Z(n4430) );
  AND U15623 ( .A(a[29]), .B(b[92]), .Z(n4429) );
  XNOR U15624 ( .A(n4434), .B(n3713), .Z(n3715) );
  XOR U15625 ( .A(n4435), .B(n4436), .Z(n3713) );
  ANDN U15626 ( .B(n4437), .A(n4438), .Z(n4435) );
  AND U15627 ( .A(a[30]), .B(b[91]), .Z(n4434) );
  XNOR U15628 ( .A(n4439), .B(n3718), .Z(n3720) );
  XOR U15629 ( .A(n4440), .B(n4441), .Z(n3718) );
  ANDN U15630 ( .B(n4442), .A(n4443), .Z(n4440) );
  AND U15631 ( .A(a[31]), .B(b[90]), .Z(n4439) );
  XNOR U15632 ( .A(n4444), .B(n3723), .Z(n3725) );
  XOR U15633 ( .A(n4445), .B(n4446), .Z(n3723) );
  ANDN U15634 ( .B(n4447), .A(n4448), .Z(n4445) );
  AND U15635 ( .A(a[32]), .B(b[89]), .Z(n4444) );
  XNOR U15636 ( .A(n4449), .B(n3728), .Z(n3730) );
  XOR U15637 ( .A(n4450), .B(n4451), .Z(n3728) );
  ANDN U15638 ( .B(n4452), .A(n4453), .Z(n4450) );
  AND U15639 ( .A(a[33]), .B(b[88]), .Z(n4449) );
  XNOR U15640 ( .A(n4454), .B(n3733), .Z(n3735) );
  XOR U15641 ( .A(n4455), .B(n4456), .Z(n3733) );
  ANDN U15642 ( .B(n4457), .A(n4458), .Z(n4455) );
  AND U15643 ( .A(a[34]), .B(b[87]), .Z(n4454) );
  XNOR U15644 ( .A(n4459), .B(n3738), .Z(n3740) );
  XOR U15645 ( .A(n4460), .B(n4461), .Z(n3738) );
  ANDN U15646 ( .B(n4462), .A(n4463), .Z(n4460) );
  AND U15647 ( .A(a[35]), .B(b[86]), .Z(n4459) );
  XNOR U15648 ( .A(n4464), .B(n3743), .Z(n3745) );
  XOR U15649 ( .A(n4465), .B(n4466), .Z(n3743) );
  ANDN U15650 ( .B(n4467), .A(n4468), .Z(n4465) );
  AND U15651 ( .A(a[36]), .B(b[85]), .Z(n4464) );
  XNOR U15652 ( .A(n4469), .B(n3748), .Z(n3750) );
  XOR U15653 ( .A(n4470), .B(n4471), .Z(n3748) );
  ANDN U15654 ( .B(n4472), .A(n4473), .Z(n4470) );
  AND U15655 ( .A(a[37]), .B(b[84]), .Z(n4469) );
  XNOR U15656 ( .A(n4474), .B(n3753), .Z(n3755) );
  XOR U15657 ( .A(n4475), .B(n4476), .Z(n3753) );
  ANDN U15658 ( .B(n4477), .A(n4478), .Z(n4475) );
  AND U15659 ( .A(a[38]), .B(b[83]), .Z(n4474) );
  XNOR U15660 ( .A(n4479), .B(n3758), .Z(n3760) );
  XOR U15661 ( .A(n4480), .B(n4481), .Z(n3758) );
  ANDN U15662 ( .B(n4482), .A(n4483), .Z(n4480) );
  AND U15663 ( .A(a[39]), .B(b[82]), .Z(n4479) );
  XNOR U15664 ( .A(n4484), .B(n3763), .Z(n3765) );
  XOR U15665 ( .A(n4485), .B(n4486), .Z(n3763) );
  ANDN U15666 ( .B(n4487), .A(n4488), .Z(n4485) );
  AND U15667 ( .A(a[40]), .B(b[81]), .Z(n4484) );
  XNOR U15668 ( .A(n4489), .B(n3768), .Z(n3770) );
  XOR U15669 ( .A(n4490), .B(n4491), .Z(n3768) );
  ANDN U15670 ( .B(n4492), .A(n4493), .Z(n4490) );
  AND U15671 ( .A(a[41]), .B(b[80]), .Z(n4489) );
  XNOR U15672 ( .A(n4494), .B(n3773), .Z(n3775) );
  XOR U15673 ( .A(n4495), .B(n4496), .Z(n3773) );
  ANDN U15674 ( .B(n4497), .A(n4498), .Z(n4495) );
  AND U15675 ( .A(a[42]), .B(b[79]), .Z(n4494) );
  XNOR U15676 ( .A(n4499), .B(n3778), .Z(n3780) );
  XOR U15677 ( .A(n4500), .B(n4501), .Z(n3778) );
  ANDN U15678 ( .B(n4502), .A(n4503), .Z(n4500) );
  AND U15679 ( .A(a[43]), .B(b[78]), .Z(n4499) );
  XNOR U15680 ( .A(n4504), .B(n3783), .Z(n3785) );
  XOR U15681 ( .A(n4505), .B(n4506), .Z(n3783) );
  ANDN U15682 ( .B(n4507), .A(n4508), .Z(n4505) );
  AND U15683 ( .A(a[44]), .B(b[77]), .Z(n4504) );
  XNOR U15684 ( .A(n4509), .B(n3788), .Z(n3790) );
  XOR U15685 ( .A(n4510), .B(n4511), .Z(n3788) );
  ANDN U15686 ( .B(n4512), .A(n4513), .Z(n4510) );
  AND U15687 ( .A(a[45]), .B(b[76]), .Z(n4509) );
  XNOR U15688 ( .A(n4514), .B(n3793), .Z(n3795) );
  XOR U15689 ( .A(n4515), .B(n4516), .Z(n3793) );
  ANDN U15690 ( .B(n4517), .A(n4518), .Z(n4515) );
  AND U15691 ( .A(a[46]), .B(b[75]), .Z(n4514) );
  XNOR U15692 ( .A(n4519), .B(n3798), .Z(n3800) );
  XOR U15693 ( .A(n4520), .B(n4521), .Z(n3798) );
  ANDN U15694 ( .B(n4522), .A(n4523), .Z(n4520) );
  AND U15695 ( .A(a[47]), .B(b[74]), .Z(n4519) );
  XNOR U15696 ( .A(n4524), .B(n3803), .Z(n3805) );
  XOR U15697 ( .A(n4525), .B(n4526), .Z(n3803) );
  ANDN U15698 ( .B(n4527), .A(n4528), .Z(n4525) );
  AND U15699 ( .A(a[48]), .B(b[73]), .Z(n4524) );
  XNOR U15700 ( .A(n4529), .B(n3808), .Z(n3810) );
  XOR U15701 ( .A(n4530), .B(n4531), .Z(n3808) );
  ANDN U15702 ( .B(n4532), .A(n4533), .Z(n4530) );
  AND U15703 ( .A(a[49]), .B(b[72]), .Z(n4529) );
  XNOR U15704 ( .A(n4534), .B(n3813), .Z(n3815) );
  XOR U15705 ( .A(n4535), .B(n4536), .Z(n3813) );
  ANDN U15706 ( .B(n4537), .A(n4538), .Z(n4535) );
  AND U15707 ( .A(a[50]), .B(b[71]), .Z(n4534) );
  XNOR U15708 ( .A(n4539), .B(n3818), .Z(n3820) );
  XOR U15709 ( .A(n4540), .B(n4541), .Z(n3818) );
  ANDN U15710 ( .B(n4542), .A(n4543), .Z(n4540) );
  AND U15711 ( .A(a[51]), .B(b[70]), .Z(n4539) );
  XNOR U15712 ( .A(n4544), .B(n3823), .Z(n3825) );
  XOR U15713 ( .A(n4545), .B(n4546), .Z(n3823) );
  ANDN U15714 ( .B(n4547), .A(n4548), .Z(n4545) );
  AND U15715 ( .A(a[52]), .B(b[69]), .Z(n4544) );
  XNOR U15716 ( .A(n4549), .B(n3828), .Z(n3830) );
  XOR U15717 ( .A(n4550), .B(n4551), .Z(n3828) );
  ANDN U15718 ( .B(n4552), .A(n4553), .Z(n4550) );
  AND U15719 ( .A(a[53]), .B(b[68]), .Z(n4549) );
  XNOR U15720 ( .A(n4554), .B(n3833), .Z(n3835) );
  XOR U15721 ( .A(n4555), .B(n4556), .Z(n3833) );
  ANDN U15722 ( .B(n4557), .A(n4558), .Z(n4555) );
  AND U15723 ( .A(a[54]), .B(b[67]), .Z(n4554) );
  XNOR U15724 ( .A(n4559), .B(n3838), .Z(n3840) );
  XOR U15725 ( .A(n4560), .B(n4561), .Z(n3838) );
  ANDN U15726 ( .B(n4562), .A(n4563), .Z(n4560) );
  AND U15727 ( .A(a[55]), .B(b[66]), .Z(n4559) );
  XNOR U15728 ( .A(n4564), .B(n3843), .Z(n3845) );
  XOR U15729 ( .A(n4565), .B(n4566), .Z(n3843) );
  ANDN U15730 ( .B(n4567), .A(n4568), .Z(n4565) );
  AND U15731 ( .A(a[56]), .B(b[65]), .Z(n4564) );
  XNOR U15732 ( .A(n4569), .B(n3848), .Z(n3850) );
  XOR U15733 ( .A(n4570), .B(n4571), .Z(n3848) );
  ANDN U15734 ( .B(n4572), .A(n4573), .Z(n4570) );
  AND U15735 ( .A(a[57]), .B(b[64]), .Z(n4569) );
  XNOR U15736 ( .A(n4574), .B(n3853), .Z(n3855) );
  XOR U15737 ( .A(n4575), .B(n4576), .Z(n3853) );
  ANDN U15738 ( .B(n4577), .A(n4578), .Z(n4575) );
  AND U15739 ( .A(a[58]), .B(b[63]), .Z(n4574) );
  XNOR U15740 ( .A(n4579), .B(n3858), .Z(n3860) );
  XOR U15741 ( .A(n4580), .B(n4581), .Z(n3858) );
  ANDN U15742 ( .B(n4582), .A(n4583), .Z(n4580) );
  AND U15743 ( .A(a[59]), .B(b[62]), .Z(n4579) );
  XNOR U15744 ( .A(n4584), .B(n3863), .Z(n3865) );
  XOR U15745 ( .A(n4585), .B(n4586), .Z(n3863) );
  ANDN U15746 ( .B(n4587), .A(n4588), .Z(n4585) );
  AND U15747 ( .A(a[60]), .B(b[61]), .Z(n4584) );
  XNOR U15748 ( .A(n4589), .B(n3868), .Z(n3870) );
  XOR U15749 ( .A(n4590), .B(n4591), .Z(n3868) );
  ANDN U15750 ( .B(n4592), .A(n4593), .Z(n4590) );
  AND U15751 ( .A(a[61]), .B(b[60]), .Z(n4589) );
  XNOR U15752 ( .A(n4594), .B(n3873), .Z(n3875) );
  XOR U15753 ( .A(n4595), .B(n4596), .Z(n3873) );
  ANDN U15754 ( .B(n4597), .A(n4598), .Z(n4595) );
  AND U15755 ( .A(a[62]), .B(b[59]), .Z(n4594) );
  XNOR U15756 ( .A(n4599), .B(n3878), .Z(n3880) );
  XOR U15757 ( .A(n4600), .B(n4601), .Z(n3878) );
  ANDN U15758 ( .B(n4602), .A(n4603), .Z(n4600) );
  AND U15759 ( .A(a[63]), .B(b[58]), .Z(n4599) );
  XNOR U15760 ( .A(n4604), .B(n3883), .Z(n3885) );
  XOR U15761 ( .A(n4605), .B(n4606), .Z(n3883) );
  ANDN U15762 ( .B(n4607), .A(n4608), .Z(n4605) );
  AND U15763 ( .A(a[64]), .B(b[57]), .Z(n4604) );
  XNOR U15764 ( .A(n4609), .B(n3888), .Z(n3890) );
  XOR U15765 ( .A(n4610), .B(n4611), .Z(n3888) );
  ANDN U15766 ( .B(n4612), .A(n4613), .Z(n4610) );
  AND U15767 ( .A(a[65]), .B(b[56]), .Z(n4609) );
  XNOR U15768 ( .A(n4614), .B(n3893), .Z(n3895) );
  XOR U15769 ( .A(n4615), .B(n4616), .Z(n3893) );
  ANDN U15770 ( .B(n4617), .A(n4618), .Z(n4615) );
  AND U15771 ( .A(a[66]), .B(b[55]), .Z(n4614) );
  XNOR U15772 ( .A(n4619), .B(n3898), .Z(n3900) );
  XOR U15773 ( .A(n4620), .B(n4621), .Z(n3898) );
  ANDN U15774 ( .B(n4622), .A(n4623), .Z(n4620) );
  AND U15775 ( .A(a[67]), .B(b[54]), .Z(n4619) );
  XNOR U15776 ( .A(n4624), .B(n3903), .Z(n3905) );
  XOR U15777 ( .A(n4625), .B(n4626), .Z(n3903) );
  ANDN U15778 ( .B(n4627), .A(n4628), .Z(n4625) );
  AND U15779 ( .A(a[68]), .B(b[53]), .Z(n4624) );
  XNOR U15780 ( .A(n4629), .B(n3908), .Z(n3910) );
  XOR U15781 ( .A(n4630), .B(n4631), .Z(n3908) );
  ANDN U15782 ( .B(n4632), .A(n4633), .Z(n4630) );
  AND U15783 ( .A(a[69]), .B(b[52]), .Z(n4629) );
  XNOR U15784 ( .A(n4634), .B(n3913), .Z(n3915) );
  XOR U15785 ( .A(n4635), .B(n4636), .Z(n3913) );
  ANDN U15786 ( .B(n4637), .A(n4638), .Z(n4635) );
  AND U15787 ( .A(a[70]), .B(b[51]), .Z(n4634) );
  XNOR U15788 ( .A(n4639), .B(n3918), .Z(n3920) );
  XOR U15789 ( .A(n4640), .B(n4641), .Z(n3918) );
  ANDN U15790 ( .B(n4642), .A(n4643), .Z(n4640) );
  AND U15791 ( .A(a[71]), .B(b[50]), .Z(n4639) );
  XNOR U15792 ( .A(n4644), .B(n3923), .Z(n3925) );
  XOR U15793 ( .A(n4645), .B(n4646), .Z(n3923) );
  ANDN U15794 ( .B(n4647), .A(n4648), .Z(n4645) );
  AND U15795 ( .A(a[72]), .B(b[49]), .Z(n4644) );
  XNOR U15796 ( .A(n4649), .B(n3928), .Z(n3930) );
  XOR U15797 ( .A(n4650), .B(n4651), .Z(n3928) );
  ANDN U15798 ( .B(n4652), .A(n4653), .Z(n4650) );
  AND U15799 ( .A(a[73]), .B(b[48]), .Z(n4649) );
  XNOR U15800 ( .A(n4654), .B(n3933), .Z(n3935) );
  XOR U15801 ( .A(n4655), .B(n4656), .Z(n3933) );
  ANDN U15802 ( .B(n4657), .A(n4658), .Z(n4655) );
  AND U15803 ( .A(a[74]), .B(b[47]), .Z(n4654) );
  XNOR U15804 ( .A(n4659), .B(n3938), .Z(n3940) );
  XOR U15805 ( .A(n4660), .B(n4661), .Z(n3938) );
  ANDN U15806 ( .B(n4662), .A(n4663), .Z(n4660) );
  AND U15807 ( .A(a[75]), .B(b[46]), .Z(n4659) );
  XNOR U15808 ( .A(n4664), .B(n3943), .Z(n3945) );
  XOR U15809 ( .A(n4665), .B(n4666), .Z(n3943) );
  ANDN U15810 ( .B(n4667), .A(n4668), .Z(n4665) );
  AND U15811 ( .A(a[76]), .B(b[45]), .Z(n4664) );
  XNOR U15812 ( .A(n4669), .B(n3948), .Z(n3950) );
  XOR U15813 ( .A(n4670), .B(n4671), .Z(n3948) );
  ANDN U15814 ( .B(n4672), .A(n4673), .Z(n4670) );
  AND U15815 ( .A(a[77]), .B(b[44]), .Z(n4669) );
  XNOR U15816 ( .A(n4674), .B(n3953), .Z(n3955) );
  XOR U15817 ( .A(n4675), .B(n4676), .Z(n3953) );
  ANDN U15818 ( .B(n4677), .A(n4678), .Z(n4675) );
  AND U15819 ( .A(a[78]), .B(b[43]), .Z(n4674) );
  XNOR U15820 ( .A(n4679), .B(n3958), .Z(n3960) );
  XOR U15821 ( .A(n4680), .B(n4681), .Z(n3958) );
  ANDN U15822 ( .B(n4682), .A(n4683), .Z(n4680) );
  AND U15823 ( .A(a[79]), .B(b[42]), .Z(n4679) );
  XNOR U15824 ( .A(n4684), .B(n3963), .Z(n3965) );
  XOR U15825 ( .A(n4685), .B(n4686), .Z(n3963) );
  ANDN U15826 ( .B(n4687), .A(n4688), .Z(n4685) );
  AND U15827 ( .A(a[80]), .B(b[41]), .Z(n4684) );
  XNOR U15828 ( .A(n4689), .B(n3968), .Z(n3970) );
  XOR U15829 ( .A(n4690), .B(n4691), .Z(n3968) );
  ANDN U15830 ( .B(n4692), .A(n4693), .Z(n4690) );
  AND U15831 ( .A(a[81]), .B(b[40]), .Z(n4689) );
  XNOR U15832 ( .A(n4694), .B(n3973), .Z(n3975) );
  XOR U15833 ( .A(n4695), .B(n4696), .Z(n3973) );
  ANDN U15834 ( .B(n4697), .A(n4698), .Z(n4695) );
  AND U15835 ( .A(a[82]), .B(b[39]), .Z(n4694) );
  XNOR U15836 ( .A(n4699), .B(n3978), .Z(n3980) );
  XOR U15837 ( .A(n4700), .B(n4701), .Z(n3978) );
  ANDN U15838 ( .B(n4702), .A(n4703), .Z(n4700) );
  AND U15839 ( .A(a[83]), .B(b[38]), .Z(n4699) );
  XNOR U15840 ( .A(n4704), .B(n3983), .Z(n3985) );
  XOR U15841 ( .A(n4705), .B(n4706), .Z(n3983) );
  ANDN U15842 ( .B(n4707), .A(n4708), .Z(n4705) );
  AND U15843 ( .A(a[84]), .B(b[37]), .Z(n4704) );
  XNOR U15844 ( .A(n4709), .B(n3988), .Z(n3990) );
  XOR U15845 ( .A(n4710), .B(n4711), .Z(n3988) );
  ANDN U15846 ( .B(n4712), .A(n4713), .Z(n4710) );
  AND U15847 ( .A(a[85]), .B(b[36]), .Z(n4709) );
  XNOR U15848 ( .A(n4714), .B(n3993), .Z(n3995) );
  XOR U15849 ( .A(n4715), .B(n4716), .Z(n3993) );
  ANDN U15850 ( .B(n4717), .A(n4718), .Z(n4715) );
  AND U15851 ( .A(a[86]), .B(b[35]), .Z(n4714) );
  XNOR U15852 ( .A(n4719), .B(n3998), .Z(n4000) );
  XOR U15853 ( .A(n4720), .B(n4721), .Z(n3998) );
  ANDN U15854 ( .B(n4722), .A(n4723), .Z(n4720) );
  AND U15855 ( .A(a[87]), .B(b[34]), .Z(n4719) );
  XNOR U15856 ( .A(n4724), .B(n4003), .Z(n4005) );
  XOR U15857 ( .A(n4725), .B(n4726), .Z(n4003) );
  ANDN U15858 ( .B(n4727), .A(n4728), .Z(n4725) );
  AND U15859 ( .A(a[88]), .B(b[33]), .Z(n4724) );
  XNOR U15860 ( .A(n4729), .B(n4008), .Z(n4010) );
  XOR U15861 ( .A(n4730), .B(n4731), .Z(n4008) );
  ANDN U15862 ( .B(n4732), .A(n4733), .Z(n4730) );
  AND U15863 ( .A(a[89]), .B(b[32]), .Z(n4729) );
  XNOR U15864 ( .A(n4734), .B(n4013), .Z(n4015) );
  XOR U15865 ( .A(n4735), .B(n4736), .Z(n4013) );
  ANDN U15866 ( .B(n4737), .A(n4738), .Z(n4735) );
  AND U15867 ( .A(a[90]), .B(b[31]), .Z(n4734) );
  XNOR U15868 ( .A(n4739), .B(n4018), .Z(n4020) );
  XOR U15869 ( .A(n4740), .B(n4741), .Z(n4018) );
  ANDN U15870 ( .B(n4742), .A(n4743), .Z(n4740) );
  AND U15871 ( .A(a[91]), .B(b[30]), .Z(n4739) );
  XNOR U15872 ( .A(n4744), .B(n4023), .Z(n4025) );
  XOR U15873 ( .A(n4745), .B(n4746), .Z(n4023) );
  ANDN U15874 ( .B(n4747), .A(n4748), .Z(n4745) );
  AND U15875 ( .A(a[92]), .B(b[29]), .Z(n4744) );
  XNOR U15876 ( .A(n4749), .B(n4028), .Z(n4030) );
  XOR U15877 ( .A(n4750), .B(n4751), .Z(n4028) );
  ANDN U15878 ( .B(n4752), .A(n4753), .Z(n4750) );
  AND U15879 ( .A(a[93]), .B(b[28]), .Z(n4749) );
  XNOR U15880 ( .A(n4754), .B(n4033), .Z(n4035) );
  XOR U15881 ( .A(n4755), .B(n4756), .Z(n4033) );
  ANDN U15882 ( .B(n4757), .A(n4758), .Z(n4755) );
  AND U15883 ( .A(a[94]), .B(b[27]), .Z(n4754) );
  XNOR U15884 ( .A(n4759), .B(n4038), .Z(n4040) );
  XOR U15885 ( .A(n4760), .B(n4761), .Z(n4038) );
  ANDN U15886 ( .B(n4762), .A(n4763), .Z(n4760) );
  AND U15887 ( .A(a[95]), .B(b[26]), .Z(n4759) );
  XNOR U15888 ( .A(n4764), .B(n4043), .Z(n4045) );
  XOR U15889 ( .A(n4765), .B(n4766), .Z(n4043) );
  ANDN U15890 ( .B(n4767), .A(n4768), .Z(n4765) );
  AND U15891 ( .A(a[96]), .B(b[25]), .Z(n4764) );
  XNOR U15892 ( .A(n4769), .B(n4048), .Z(n4050) );
  XOR U15893 ( .A(n4770), .B(n4771), .Z(n4048) );
  ANDN U15894 ( .B(n4772), .A(n4773), .Z(n4770) );
  AND U15895 ( .A(a[97]), .B(b[24]), .Z(n4769) );
  XNOR U15896 ( .A(n4774), .B(n4053), .Z(n4055) );
  XOR U15897 ( .A(n4775), .B(n4776), .Z(n4053) );
  ANDN U15898 ( .B(n4777), .A(n4778), .Z(n4775) );
  AND U15899 ( .A(a[98]), .B(b[23]), .Z(n4774) );
  XNOR U15900 ( .A(n4779), .B(n4058), .Z(n4060) );
  XOR U15901 ( .A(n4780), .B(n4781), .Z(n4058) );
  ANDN U15902 ( .B(n4782), .A(n4783), .Z(n4780) );
  AND U15903 ( .A(a[99]), .B(b[22]), .Z(n4779) );
  XNOR U15904 ( .A(n4784), .B(n4063), .Z(n4065) );
  XOR U15905 ( .A(n4785), .B(n4786), .Z(n4063) );
  ANDN U15906 ( .B(n4787), .A(n4788), .Z(n4785) );
  AND U15907 ( .A(b[21]), .B(a[100]), .Z(n4784) );
  XNOR U15908 ( .A(n4789), .B(n4068), .Z(n4070) );
  XOR U15909 ( .A(n4790), .B(n4791), .Z(n4068) );
  ANDN U15910 ( .B(n4792), .A(n4793), .Z(n4790) );
  AND U15911 ( .A(b[20]), .B(a[101]), .Z(n4789) );
  XNOR U15912 ( .A(n4794), .B(n4073), .Z(n4075) );
  XOR U15913 ( .A(n4795), .B(n4796), .Z(n4073) );
  ANDN U15914 ( .B(n4797), .A(n4798), .Z(n4795) );
  AND U15915 ( .A(b[19]), .B(a[102]), .Z(n4794) );
  XNOR U15916 ( .A(n4799), .B(n4078), .Z(n4080) );
  XOR U15917 ( .A(n4800), .B(n4801), .Z(n4078) );
  ANDN U15918 ( .B(n4802), .A(n4803), .Z(n4800) );
  AND U15919 ( .A(b[18]), .B(a[103]), .Z(n4799) );
  XNOR U15920 ( .A(n4804), .B(n4083), .Z(n4085) );
  XOR U15921 ( .A(n4805), .B(n4806), .Z(n4083) );
  ANDN U15922 ( .B(n4807), .A(n4808), .Z(n4805) );
  AND U15923 ( .A(b[17]), .B(a[104]), .Z(n4804) );
  XNOR U15924 ( .A(n4809), .B(n4088), .Z(n4090) );
  XOR U15925 ( .A(n4810), .B(n4811), .Z(n4088) );
  ANDN U15926 ( .B(n4812), .A(n4813), .Z(n4810) );
  AND U15927 ( .A(b[16]), .B(a[105]), .Z(n4809) );
  XNOR U15928 ( .A(n4814), .B(n4093), .Z(n4095) );
  XOR U15929 ( .A(n4815), .B(n4816), .Z(n4093) );
  ANDN U15930 ( .B(n4817), .A(n4818), .Z(n4815) );
  AND U15931 ( .A(b[15]), .B(a[106]), .Z(n4814) );
  XNOR U15932 ( .A(n4819), .B(n4098), .Z(n4100) );
  XOR U15933 ( .A(n4820), .B(n4821), .Z(n4098) );
  ANDN U15934 ( .B(n4822), .A(n4823), .Z(n4820) );
  AND U15935 ( .A(b[14]), .B(a[107]), .Z(n4819) );
  XNOR U15936 ( .A(n4824), .B(n4103), .Z(n4105) );
  XOR U15937 ( .A(n4825), .B(n4826), .Z(n4103) );
  ANDN U15938 ( .B(n4827), .A(n4828), .Z(n4825) );
  AND U15939 ( .A(b[13]), .B(a[108]), .Z(n4824) );
  XNOR U15940 ( .A(n4829), .B(n4108), .Z(n4110) );
  XOR U15941 ( .A(n4830), .B(n4831), .Z(n4108) );
  ANDN U15942 ( .B(n4832), .A(n4833), .Z(n4830) );
  AND U15943 ( .A(b[12]), .B(a[109]), .Z(n4829) );
  XNOR U15944 ( .A(n4834), .B(n4113), .Z(n4115) );
  XOR U15945 ( .A(n4835), .B(n4836), .Z(n4113) );
  ANDN U15946 ( .B(n4837), .A(n4838), .Z(n4835) );
  AND U15947 ( .A(b[11]), .B(a[110]), .Z(n4834) );
  XNOR U15948 ( .A(n4839), .B(n4118), .Z(n4120) );
  XOR U15949 ( .A(n4840), .B(n4841), .Z(n4118) );
  ANDN U15950 ( .B(n4842), .A(n4843), .Z(n4840) );
  AND U15951 ( .A(b[10]), .B(a[111]), .Z(n4839) );
  XNOR U15952 ( .A(n4844), .B(n4123), .Z(n4125) );
  XOR U15953 ( .A(n4845), .B(n4846), .Z(n4123) );
  ANDN U15954 ( .B(n4847), .A(n4848), .Z(n4845) );
  AND U15955 ( .A(b[9]), .B(a[112]), .Z(n4844) );
  XNOR U15956 ( .A(n4849), .B(n4128), .Z(n4130) );
  XOR U15957 ( .A(n4850), .B(n4851), .Z(n4128) );
  ANDN U15958 ( .B(n4852), .A(n4853), .Z(n4850) );
  AND U15959 ( .A(b[8]), .B(a[113]), .Z(n4849) );
  XNOR U15960 ( .A(n4854), .B(n4133), .Z(n4135) );
  XOR U15961 ( .A(n4855), .B(n4856), .Z(n4133) );
  ANDN U15962 ( .B(n4857), .A(n4858), .Z(n4855) );
  AND U15963 ( .A(b[7]), .B(a[114]), .Z(n4854) );
  XNOR U15964 ( .A(n4859), .B(n4138), .Z(n4140) );
  XOR U15965 ( .A(n4860), .B(n4861), .Z(n4138) );
  ANDN U15966 ( .B(n4862), .A(n4863), .Z(n4860) );
  AND U15967 ( .A(b[6]), .B(a[115]), .Z(n4859) );
  XNOR U15968 ( .A(n4864), .B(n4143), .Z(n4145) );
  XOR U15969 ( .A(n4865), .B(n4866), .Z(n4143) );
  ANDN U15970 ( .B(n4867), .A(n4868), .Z(n4865) );
  AND U15971 ( .A(b[5]), .B(a[116]), .Z(n4864) );
  XNOR U15972 ( .A(n4869), .B(n4148), .Z(n4150) );
  XOR U15973 ( .A(n4870), .B(n4871), .Z(n4148) );
  ANDN U15974 ( .B(n4872), .A(n4873), .Z(n4870) );
  AND U15975 ( .A(b[4]), .B(a[117]), .Z(n4869) );
  XNOR U15976 ( .A(n4874), .B(n4875), .Z(n4162) );
  NANDN U15977 ( .A(n4876), .B(n4877), .Z(n4875) );
  XNOR U15978 ( .A(n4878), .B(n4153), .Z(n4155) );
  XNOR U15979 ( .A(n4879), .B(n4880), .Z(n4153) );
  AND U15980 ( .A(n4881), .B(n4882), .Z(n4879) );
  AND U15981 ( .A(b[3]), .B(a[118]), .Z(n4878) );
  NAND U15982 ( .A(a[121]), .B(b[0]), .Z(n3444) );
  XNOR U15983 ( .A(n4168), .B(n4169), .Z(c[120]) );
  XNOR U15984 ( .A(n4876), .B(n4877), .Z(n4169) );
  XOR U15985 ( .A(n4874), .B(n4883), .Z(n4877) );
  NAND U15986 ( .A(b[1]), .B(a[119]), .Z(n4883) );
  XOR U15987 ( .A(n4882), .B(n4884), .Z(n4876) );
  XOR U15988 ( .A(n4874), .B(n4881), .Z(n4884) );
  XNOR U15989 ( .A(n4885), .B(n4880), .Z(n4881) );
  AND U15990 ( .A(b[2]), .B(a[118]), .Z(n4885) );
  NANDN U15991 ( .A(n4886), .B(n4887), .Z(n4874) );
  XOR U15992 ( .A(n4880), .B(n4872), .Z(n4888) );
  XNOR U15993 ( .A(n4871), .B(n4867), .Z(n4889) );
  XNOR U15994 ( .A(n4866), .B(n4862), .Z(n4890) );
  XNOR U15995 ( .A(n4861), .B(n4857), .Z(n4891) );
  XNOR U15996 ( .A(n4856), .B(n4852), .Z(n4892) );
  XNOR U15997 ( .A(n4851), .B(n4847), .Z(n4893) );
  XNOR U15998 ( .A(n4846), .B(n4842), .Z(n4894) );
  XNOR U15999 ( .A(n4841), .B(n4837), .Z(n4895) );
  XNOR U16000 ( .A(n4836), .B(n4832), .Z(n4896) );
  XNOR U16001 ( .A(n4831), .B(n4827), .Z(n4897) );
  XNOR U16002 ( .A(n4826), .B(n4822), .Z(n4898) );
  XNOR U16003 ( .A(n4821), .B(n4817), .Z(n4899) );
  XNOR U16004 ( .A(n4816), .B(n4812), .Z(n4900) );
  XNOR U16005 ( .A(n4811), .B(n4807), .Z(n4901) );
  XNOR U16006 ( .A(n4806), .B(n4802), .Z(n4902) );
  XNOR U16007 ( .A(n4801), .B(n4797), .Z(n4903) );
  XNOR U16008 ( .A(n4796), .B(n4792), .Z(n4904) );
  XNOR U16009 ( .A(n4791), .B(n4787), .Z(n4905) );
  XNOR U16010 ( .A(n4786), .B(n4782), .Z(n4906) );
  XNOR U16011 ( .A(n4781), .B(n4777), .Z(n4907) );
  XNOR U16012 ( .A(n4776), .B(n4772), .Z(n4908) );
  XNOR U16013 ( .A(n4771), .B(n4767), .Z(n4909) );
  XNOR U16014 ( .A(n4766), .B(n4762), .Z(n4910) );
  XNOR U16015 ( .A(n4761), .B(n4757), .Z(n4911) );
  XNOR U16016 ( .A(n4756), .B(n4752), .Z(n4912) );
  XNOR U16017 ( .A(n4751), .B(n4747), .Z(n4913) );
  XNOR U16018 ( .A(n4746), .B(n4742), .Z(n4914) );
  XNOR U16019 ( .A(n4741), .B(n4737), .Z(n4915) );
  XNOR U16020 ( .A(n4736), .B(n4732), .Z(n4916) );
  XNOR U16021 ( .A(n4731), .B(n4727), .Z(n4917) );
  XNOR U16022 ( .A(n4726), .B(n4722), .Z(n4918) );
  XNOR U16023 ( .A(n4721), .B(n4717), .Z(n4919) );
  XNOR U16024 ( .A(n4716), .B(n4712), .Z(n4920) );
  XNOR U16025 ( .A(n4711), .B(n4707), .Z(n4921) );
  XNOR U16026 ( .A(n4706), .B(n4702), .Z(n4922) );
  XNOR U16027 ( .A(n4701), .B(n4697), .Z(n4923) );
  XNOR U16028 ( .A(n4696), .B(n4692), .Z(n4924) );
  XNOR U16029 ( .A(n4691), .B(n4687), .Z(n4925) );
  XNOR U16030 ( .A(n4686), .B(n4682), .Z(n4926) );
  XNOR U16031 ( .A(n4681), .B(n4677), .Z(n4927) );
  XNOR U16032 ( .A(n4676), .B(n4672), .Z(n4928) );
  XNOR U16033 ( .A(n4671), .B(n4667), .Z(n4929) );
  XNOR U16034 ( .A(n4666), .B(n4662), .Z(n4930) );
  XNOR U16035 ( .A(n4661), .B(n4657), .Z(n4931) );
  XNOR U16036 ( .A(n4656), .B(n4652), .Z(n4932) );
  XNOR U16037 ( .A(n4651), .B(n4647), .Z(n4933) );
  XNOR U16038 ( .A(n4646), .B(n4642), .Z(n4934) );
  XNOR U16039 ( .A(n4641), .B(n4637), .Z(n4935) );
  XNOR U16040 ( .A(n4636), .B(n4632), .Z(n4936) );
  XNOR U16041 ( .A(n4631), .B(n4627), .Z(n4937) );
  XNOR U16042 ( .A(n4626), .B(n4622), .Z(n4938) );
  XNOR U16043 ( .A(n4621), .B(n4617), .Z(n4939) );
  XNOR U16044 ( .A(n4616), .B(n4612), .Z(n4940) );
  XNOR U16045 ( .A(n4611), .B(n4607), .Z(n4941) );
  XNOR U16046 ( .A(n4606), .B(n4602), .Z(n4942) );
  XNOR U16047 ( .A(n4601), .B(n4597), .Z(n4943) );
  XNOR U16048 ( .A(n4596), .B(n4592), .Z(n4944) );
  XNOR U16049 ( .A(n4591), .B(n4587), .Z(n4945) );
  XNOR U16050 ( .A(n4586), .B(n4582), .Z(n4946) );
  XNOR U16051 ( .A(n4581), .B(n4577), .Z(n4947) );
  XNOR U16052 ( .A(n4576), .B(n4572), .Z(n4948) );
  XNOR U16053 ( .A(n4571), .B(n4567), .Z(n4949) );
  XNOR U16054 ( .A(n4566), .B(n4562), .Z(n4950) );
  XNOR U16055 ( .A(n4561), .B(n4557), .Z(n4951) );
  XNOR U16056 ( .A(n4556), .B(n4552), .Z(n4952) );
  XNOR U16057 ( .A(n4551), .B(n4547), .Z(n4953) );
  XNOR U16058 ( .A(n4546), .B(n4542), .Z(n4954) );
  XNOR U16059 ( .A(n4541), .B(n4537), .Z(n4955) );
  XNOR U16060 ( .A(n4536), .B(n4532), .Z(n4956) );
  XNOR U16061 ( .A(n4531), .B(n4527), .Z(n4957) );
  XNOR U16062 ( .A(n4526), .B(n4522), .Z(n4958) );
  XNOR U16063 ( .A(n4521), .B(n4517), .Z(n4959) );
  XNOR U16064 ( .A(n4516), .B(n4512), .Z(n4960) );
  XNOR U16065 ( .A(n4511), .B(n4507), .Z(n4961) );
  XNOR U16066 ( .A(n4506), .B(n4502), .Z(n4962) );
  XNOR U16067 ( .A(n4501), .B(n4497), .Z(n4963) );
  XNOR U16068 ( .A(n4496), .B(n4492), .Z(n4964) );
  XNOR U16069 ( .A(n4491), .B(n4487), .Z(n4965) );
  XNOR U16070 ( .A(n4486), .B(n4482), .Z(n4966) );
  XNOR U16071 ( .A(n4481), .B(n4477), .Z(n4967) );
  XNOR U16072 ( .A(n4476), .B(n4472), .Z(n4968) );
  XNOR U16073 ( .A(n4471), .B(n4467), .Z(n4969) );
  XNOR U16074 ( .A(n4466), .B(n4462), .Z(n4970) );
  XNOR U16075 ( .A(n4461), .B(n4457), .Z(n4971) );
  XNOR U16076 ( .A(n4456), .B(n4452), .Z(n4972) );
  XNOR U16077 ( .A(n4451), .B(n4447), .Z(n4973) );
  XNOR U16078 ( .A(n4446), .B(n4442), .Z(n4974) );
  XNOR U16079 ( .A(n4441), .B(n4437), .Z(n4975) );
  XNOR U16080 ( .A(n4436), .B(n4432), .Z(n4976) );
  XNOR U16081 ( .A(n4431), .B(n4427), .Z(n4977) );
  XNOR U16082 ( .A(n4426), .B(n4422), .Z(n4978) );
  XNOR U16083 ( .A(n4421), .B(n4417), .Z(n4979) );
  XNOR U16084 ( .A(n4416), .B(n4412), .Z(n4980) );
  XNOR U16085 ( .A(n4411), .B(n4407), .Z(n4981) );
  XNOR U16086 ( .A(n4406), .B(n4402), .Z(n4982) );
  XNOR U16087 ( .A(n4401), .B(n4397), .Z(n4983) );
  XNOR U16088 ( .A(n4396), .B(n4392), .Z(n4984) );
  XNOR U16089 ( .A(n4391), .B(n4387), .Z(n4985) );
  XNOR U16090 ( .A(n4386), .B(n4382), .Z(n4986) );
  XNOR U16091 ( .A(n4381), .B(n4377), .Z(n4987) );
  XNOR U16092 ( .A(n4376), .B(n4372), .Z(n4988) );
  XNOR U16093 ( .A(n4371), .B(n4367), .Z(n4989) );
  XNOR U16094 ( .A(n4366), .B(n4362), .Z(n4990) );
  XNOR U16095 ( .A(n4361), .B(n4357), .Z(n4991) );
  XNOR U16096 ( .A(n4356), .B(n4352), .Z(n4992) );
  XNOR U16097 ( .A(n4351), .B(n4347), .Z(n4993) );
  XNOR U16098 ( .A(n4346), .B(n4342), .Z(n4994) );
  XNOR U16099 ( .A(n4341), .B(n4337), .Z(n4995) );
  XNOR U16100 ( .A(n4336), .B(n4332), .Z(n4996) );
  XNOR U16101 ( .A(n4331), .B(n4327), .Z(n4997) );
  XNOR U16102 ( .A(n4326), .B(n4322), .Z(n4998) );
  XNOR U16103 ( .A(n4321), .B(n4317), .Z(n4999) );
  XNOR U16104 ( .A(n4316), .B(n4312), .Z(n5000) );
  XNOR U16105 ( .A(n4311), .B(n4307), .Z(n5001) );
  XNOR U16106 ( .A(n4306), .B(n4302), .Z(n5002) );
  XNOR U16107 ( .A(n4301), .B(n4297), .Z(n5003) );
  XNOR U16108 ( .A(n4296), .B(n4292), .Z(n5004) );
  XOR U16109 ( .A(n5005), .B(n4291), .Z(n4292) );
  AND U16110 ( .A(a[0]), .B(b[120]), .Z(n5005) );
  XNOR U16111 ( .A(n5006), .B(n4291), .Z(n4293) );
  XNOR U16112 ( .A(n5007), .B(n5008), .Z(n4291) );
  ANDN U16113 ( .B(n5009), .A(n5010), .Z(n5007) );
  AND U16114 ( .A(a[1]), .B(b[119]), .Z(n5006) );
  XNOR U16115 ( .A(n5011), .B(n4296), .Z(n4298) );
  XOR U16116 ( .A(n5012), .B(n5013), .Z(n4296) );
  ANDN U16117 ( .B(n5014), .A(n5015), .Z(n5012) );
  AND U16118 ( .A(a[2]), .B(b[118]), .Z(n5011) );
  XNOR U16119 ( .A(n5016), .B(n4301), .Z(n4303) );
  XOR U16120 ( .A(n5017), .B(n5018), .Z(n4301) );
  ANDN U16121 ( .B(n5019), .A(n5020), .Z(n5017) );
  AND U16122 ( .A(a[3]), .B(b[117]), .Z(n5016) );
  XNOR U16123 ( .A(n5021), .B(n4306), .Z(n4308) );
  XOR U16124 ( .A(n5022), .B(n5023), .Z(n4306) );
  ANDN U16125 ( .B(n5024), .A(n5025), .Z(n5022) );
  AND U16126 ( .A(a[4]), .B(b[116]), .Z(n5021) );
  XNOR U16127 ( .A(n5026), .B(n4311), .Z(n4313) );
  XOR U16128 ( .A(n5027), .B(n5028), .Z(n4311) );
  ANDN U16129 ( .B(n5029), .A(n5030), .Z(n5027) );
  AND U16130 ( .A(a[5]), .B(b[115]), .Z(n5026) );
  XNOR U16131 ( .A(n5031), .B(n4316), .Z(n4318) );
  XOR U16132 ( .A(n5032), .B(n5033), .Z(n4316) );
  ANDN U16133 ( .B(n5034), .A(n5035), .Z(n5032) );
  AND U16134 ( .A(a[6]), .B(b[114]), .Z(n5031) );
  XNOR U16135 ( .A(n5036), .B(n4321), .Z(n4323) );
  XOR U16136 ( .A(n5037), .B(n5038), .Z(n4321) );
  ANDN U16137 ( .B(n5039), .A(n5040), .Z(n5037) );
  AND U16138 ( .A(a[7]), .B(b[113]), .Z(n5036) );
  XNOR U16139 ( .A(n5041), .B(n4326), .Z(n4328) );
  XOR U16140 ( .A(n5042), .B(n5043), .Z(n4326) );
  ANDN U16141 ( .B(n5044), .A(n5045), .Z(n5042) );
  AND U16142 ( .A(a[8]), .B(b[112]), .Z(n5041) );
  XNOR U16143 ( .A(n5046), .B(n4331), .Z(n4333) );
  XOR U16144 ( .A(n5047), .B(n5048), .Z(n4331) );
  ANDN U16145 ( .B(n5049), .A(n5050), .Z(n5047) );
  AND U16146 ( .A(a[9]), .B(b[111]), .Z(n5046) );
  XNOR U16147 ( .A(n5051), .B(n4336), .Z(n4338) );
  XOR U16148 ( .A(n5052), .B(n5053), .Z(n4336) );
  ANDN U16149 ( .B(n5054), .A(n5055), .Z(n5052) );
  AND U16150 ( .A(a[10]), .B(b[110]), .Z(n5051) );
  XNOR U16151 ( .A(n5056), .B(n4341), .Z(n4343) );
  XOR U16152 ( .A(n5057), .B(n5058), .Z(n4341) );
  ANDN U16153 ( .B(n5059), .A(n5060), .Z(n5057) );
  AND U16154 ( .A(a[11]), .B(b[109]), .Z(n5056) );
  XNOR U16155 ( .A(n5061), .B(n4346), .Z(n4348) );
  XOR U16156 ( .A(n5062), .B(n5063), .Z(n4346) );
  ANDN U16157 ( .B(n5064), .A(n5065), .Z(n5062) );
  AND U16158 ( .A(a[12]), .B(b[108]), .Z(n5061) );
  XNOR U16159 ( .A(n5066), .B(n4351), .Z(n4353) );
  XOR U16160 ( .A(n5067), .B(n5068), .Z(n4351) );
  ANDN U16161 ( .B(n5069), .A(n5070), .Z(n5067) );
  AND U16162 ( .A(a[13]), .B(b[107]), .Z(n5066) );
  XNOR U16163 ( .A(n5071), .B(n4356), .Z(n4358) );
  XOR U16164 ( .A(n5072), .B(n5073), .Z(n4356) );
  ANDN U16165 ( .B(n5074), .A(n5075), .Z(n5072) );
  AND U16166 ( .A(a[14]), .B(b[106]), .Z(n5071) );
  XNOR U16167 ( .A(n5076), .B(n4361), .Z(n4363) );
  XOR U16168 ( .A(n5077), .B(n5078), .Z(n4361) );
  ANDN U16169 ( .B(n5079), .A(n5080), .Z(n5077) );
  AND U16170 ( .A(a[15]), .B(b[105]), .Z(n5076) );
  XNOR U16171 ( .A(n5081), .B(n4366), .Z(n4368) );
  XOR U16172 ( .A(n5082), .B(n5083), .Z(n4366) );
  ANDN U16173 ( .B(n5084), .A(n5085), .Z(n5082) );
  AND U16174 ( .A(a[16]), .B(b[104]), .Z(n5081) );
  XNOR U16175 ( .A(n5086), .B(n4371), .Z(n4373) );
  XOR U16176 ( .A(n5087), .B(n5088), .Z(n4371) );
  ANDN U16177 ( .B(n5089), .A(n5090), .Z(n5087) );
  AND U16178 ( .A(a[17]), .B(b[103]), .Z(n5086) );
  XNOR U16179 ( .A(n5091), .B(n4376), .Z(n4378) );
  XOR U16180 ( .A(n5092), .B(n5093), .Z(n4376) );
  ANDN U16181 ( .B(n5094), .A(n5095), .Z(n5092) );
  AND U16182 ( .A(a[18]), .B(b[102]), .Z(n5091) );
  XNOR U16183 ( .A(n5096), .B(n4381), .Z(n4383) );
  XOR U16184 ( .A(n5097), .B(n5098), .Z(n4381) );
  ANDN U16185 ( .B(n5099), .A(n5100), .Z(n5097) );
  AND U16186 ( .A(a[19]), .B(b[101]), .Z(n5096) );
  XNOR U16187 ( .A(n5101), .B(n4386), .Z(n4388) );
  XOR U16188 ( .A(n5102), .B(n5103), .Z(n4386) );
  ANDN U16189 ( .B(n5104), .A(n5105), .Z(n5102) );
  AND U16190 ( .A(a[20]), .B(b[100]), .Z(n5101) );
  XNOR U16191 ( .A(n5106), .B(n4391), .Z(n4393) );
  XOR U16192 ( .A(n5107), .B(n5108), .Z(n4391) );
  ANDN U16193 ( .B(n5109), .A(n5110), .Z(n5107) );
  AND U16194 ( .A(a[21]), .B(b[99]), .Z(n5106) );
  XNOR U16195 ( .A(n5111), .B(n4396), .Z(n4398) );
  XOR U16196 ( .A(n5112), .B(n5113), .Z(n4396) );
  ANDN U16197 ( .B(n5114), .A(n5115), .Z(n5112) );
  AND U16198 ( .A(a[22]), .B(b[98]), .Z(n5111) );
  XNOR U16199 ( .A(n5116), .B(n4401), .Z(n4403) );
  XOR U16200 ( .A(n5117), .B(n5118), .Z(n4401) );
  ANDN U16201 ( .B(n5119), .A(n5120), .Z(n5117) );
  AND U16202 ( .A(a[23]), .B(b[97]), .Z(n5116) );
  XNOR U16203 ( .A(n5121), .B(n4406), .Z(n4408) );
  XOR U16204 ( .A(n5122), .B(n5123), .Z(n4406) );
  ANDN U16205 ( .B(n5124), .A(n5125), .Z(n5122) );
  AND U16206 ( .A(a[24]), .B(b[96]), .Z(n5121) );
  XNOR U16207 ( .A(n5126), .B(n4411), .Z(n4413) );
  XOR U16208 ( .A(n5127), .B(n5128), .Z(n4411) );
  ANDN U16209 ( .B(n5129), .A(n5130), .Z(n5127) );
  AND U16210 ( .A(a[25]), .B(b[95]), .Z(n5126) );
  XNOR U16211 ( .A(n5131), .B(n4416), .Z(n4418) );
  XOR U16212 ( .A(n5132), .B(n5133), .Z(n4416) );
  ANDN U16213 ( .B(n5134), .A(n5135), .Z(n5132) );
  AND U16214 ( .A(a[26]), .B(b[94]), .Z(n5131) );
  XNOR U16215 ( .A(n5136), .B(n4421), .Z(n4423) );
  XOR U16216 ( .A(n5137), .B(n5138), .Z(n4421) );
  ANDN U16217 ( .B(n5139), .A(n5140), .Z(n5137) );
  AND U16218 ( .A(a[27]), .B(b[93]), .Z(n5136) );
  XNOR U16219 ( .A(n5141), .B(n4426), .Z(n4428) );
  XOR U16220 ( .A(n5142), .B(n5143), .Z(n4426) );
  ANDN U16221 ( .B(n5144), .A(n5145), .Z(n5142) );
  AND U16222 ( .A(a[28]), .B(b[92]), .Z(n5141) );
  XNOR U16223 ( .A(n5146), .B(n4431), .Z(n4433) );
  XOR U16224 ( .A(n5147), .B(n5148), .Z(n4431) );
  ANDN U16225 ( .B(n5149), .A(n5150), .Z(n5147) );
  AND U16226 ( .A(a[29]), .B(b[91]), .Z(n5146) );
  XNOR U16227 ( .A(n5151), .B(n4436), .Z(n4438) );
  XOR U16228 ( .A(n5152), .B(n5153), .Z(n4436) );
  ANDN U16229 ( .B(n5154), .A(n5155), .Z(n5152) );
  AND U16230 ( .A(a[30]), .B(b[90]), .Z(n5151) );
  XNOR U16231 ( .A(n5156), .B(n4441), .Z(n4443) );
  XOR U16232 ( .A(n5157), .B(n5158), .Z(n4441) );
  ANDN U16233 ( .B(n5159), .A(n5160), .Z(n5157) );
  AND U16234 ( .A(a[31]), .B(b[89]), .Z(n5156) );
  XNOR U16235 ( .A(n5161), .B(n4446), .Z(n4448) );
  XOR U16236 ( .A(n5162), .B(n5163), .Z(n4446) );
  ANDN U16237 ( .B(n5164), .A(n5165), .Z(n5162) );
  AND U16238 ( .A(a[32]), .B(b[88]), .Z(n5161) );
  XNOR U16239 ( .A(n5166), .B(n4451), .Z(n4453) );
  XOR U16240 ( .A(n5167), .B(n5168), .Z(n4451) );
  ANDN U16241 ( .B(n5169), .A(n5170), .Z(n5167) );
  AND U16242 ( .A(a[33]), .B(b[87]), .Z(n5166) );
  XNOR U16243 ( .A(n5171), .B(n4456), .Z(n4458) );
  XOR U16244 ( .A(n5172), .B(n5173), .Z(n4456) );
  ANDN U16245 ( .B(n5174), .A(n5175), .Z(n5172) );
  AND U16246 ( .A(a[34]), .B(b[86]), .Z(n5171) );
  XNOR U16247 ( .A(n5176), .B(n4461), .Z(n4463) );
  XOR U16248 ( .A(n5177), .B(n5178), .Z(n4461) );
  ANDN U16249 ( .B(n5179), .A(n5180), .Z(n5177) );
  AND U16250 ( .A(a[35]), .B(b[85]), .Z(n5176) );
  XNOR U16251 ( .A(n5181), .B(n4466), .Z(n4468) );
  XOR U16252 ( .A(n5182), .B(n5183), .Z(n4466) );
  ANDN U16253 ( .B(n5184), .A(n5185), .Z(n5182) );
  AND U16254 ( .A(a[36]), .B(b[84]), .Z(n5181) );
  XNOR U16255 ( .A(n5186), .B(n4471), .Z(n4473) );
  XOR U16256 ( .A(n5187), .B(n5188), .Z(n4471) );
  ANDN U16257 ( .B(n5189), .A(n5190), .Z(n5187) );
  AND U16258 ( .A(a[37]), .B(b[83]), .Z(n5186) );
  XNOR U16259 ( .A(n5191), .B(n4476), .Z(n4478) );
  XOR U16260 ( .A(n5192), .B(n5193), .Z(n4476) );
  ANDN U16261 ( .B(n5194), .A(n5195), .Z(n5192) );
  AND U16262 ( .A(a[38]), .B(b[82]), .Z(n5191) );
  XNOR U16263 ( .A(n5196), .B(n4481), .Z(n4483) );
  XOR U16264 ( .A(n5197), .B(n5198), .Z(n4481) );
  ANDN U16265 ( .B(n5199), .A(n5200), .Z(n5197) );
  AND U16266 ( .A(a[39]), .B(b[81]), .Z(n5196) );
  XNOR U16267 ( .A(n5201), .B(n4486), .Z(n4488) );
  XOR U16268 ( .A(n5202), .B(n5203), .Z(n4486) );
  ANDN U16269 ( .B(n5204), .A(n5205), .Z(n5202) );
  AND U16270 ( .A(a[40]), .B(b[80]), .Z(n5201) );
  XNOR U16271 ( .A(n5206), .B(n4491), .Z(n4493) );
  XOR U16272 ( .A(n5207), .B(n5208), .Z(n4491) );
  ANDN U16273 ( .B(n5209), .A(n5210), .Z(n5207) );
  AND U16274 ( .A(a[41]), .B(b[79]), .Z(n5206) );
  XNOR U16275 ( .A(n5211), .B(n4496), .Z(n4498) );
  XOR U16276 ( .A(n5212), .B(n5213), .Z(n4496) );
  ANDN U16277 ( .B(n5214), .A(n5215), .Z(n5212) );
  AND U16278 ( .A(a[42]), .B(b[78]), .Z(n5211) );
  XNOR U16279 ( .A(n5216), .B(n4501), .Z(n4503) );
  XOR U16280 ( .A(n5217), .B(n5218), .Z(n4501) );
  ANDN U16281 ( .B(n5219), .A(n5220), .Z(n5217) );
  AND U16282 ( .A(a[43]), .B(b[77]), .Z(n5216) );
  XNOR U16283 ( .A(n5221), .B(n4506), .Z(n4508) );
  XOR U16284 ( .A(n5222), .B(n5223), .Z(n4506) );
  ANDN U16285 ( .B(n5224), .A(n5225), .Z(n5222) );
  AND U16286 ( .A(a[44]), .B(b[76]), .Z(n5221) );
  XNOR U16287 ( .A(n5226), .B(n4511), .Z(n4513) );
  XOR U16288 ( .A(n5227), .B(n5228), .Z(n4511) );
  ANDN U16289 ( .B(n5229), .A(n5230), .Z(n5227) );
  AND U16290 ( .A(a[45]), .B(b[75]), .Z(n5226) );
  XNOR U16291 ( .A(n5231), .B(n4516), .Z(n4518) );
  XOR U16292 ( .A(n5232), .B(n5233), .Z(n4516) );
  ANDN U16293 ( .B(n5234), .A(n5235), .Z(n5232) );
  AND U16294 ( .A(a[46]), .B(b[74]), .Z(n5231) );
  XNOR U16295 ( .A(n5236), .B(n4521), .Z(n4523) );
  XOR U16296 ( .A(n5237), .B(n5238), .Z(n4521) );
  ANDN U16297 ( .B(n5239), .A(n5240), .Z(n5237) );
  AND U16298 ( .A(a[47]), .B(b[73]), .Z(n5236) );
  XNOR U16299 ( .A(n5241), .B(n4526), .Z(n4528) );
  XOR U16300 ( .A(n5242), .B(n5243), .Z(n4526) );
  ANDN U16301 ( .B(n5244), .A(n5245), .Z(n5242) );
  AND U16302 ( .A(a[48]), .B(b[72]), .Z(n5241) );
  XNOR U16303 ( .A(n5246), .B(n4531), .Z(n4533) );
  XOR U16304 ( .A(n5247), .B(n5248), .Z(n4531) );
  ANDN U16305 ( .B(n5249), .A(n5250), .Z(n5247) );
  AND U16306 ( .A(a[49]), .B(b[71]), .Z(n5246) );
  XNOR U16307 ( .A(n5251), .B(n4536), .Z(n4538) );
  XOR U16308 ( .A(n5252), .B(n5253), .Z(n4536) );
  ANDN U16309 ( .B(n5254), .A(n5255), .Z(n5252) );
  AND U16310 ( .A(a[50]), .B(b[70]), .Z(n5251) );
  XNOR U16311 ( .A(n5256), .B(n4541), .Z(n4543) );
  XOR U16312 ( .A(n5257), .B(n5258), .Z(n4541) );
  ANDN U16313 ( .B(n5259), .A(n5260), .Z(n5257) );
  AND U16314 ( .A(a[51]), .B(b[69]), .Z(n5256) );
  XNOR U16315 ( .A(n5261), .B(n4546), .Z(n4548) );
  XOR U16316 ( .A(n5262), .B(n5263), .Z(n4546) );
  ANDN U16317 ( .B(n5264), .A(n5265), .Z(n5262) );
  AND U16318 ( .A(a[52]), .B(b[68]), .Z(n5261) );
  XNOR U16319 ( .A(n5266), .B(n4551), .Z(n4553) );
  XOR U16320 ( .A(n5267), .B(n5268), .Z(n4551) );
  ANDN U16321 ( .B(n5269), .A(n5270), .Z(n5267) );
  AND U16322 ( .A(a[53]), .B(b[67]), .Z(n5266) );
  XNOR U16323 ( .A(n5271), .B(n4556), .Z(n4558) );
  XOR U16324 ( .A(n5272), .B(n5273), .Z(n4556) );
  ANDN U16325 ( .B(n5274), .A(n5275), .Z(n5272) );
  AND U16326 ( .A(a[54]), .B(b[66]), .Z(n5271) );
  XNOR U16327 ( .A(n5276), .B(n4561), .Z(n4563) );
  XOR U16328 ( .A(n5277), .B(n5278), .Z(n4561) );
  ANDN U16329 ( .B(n5279), .A(n5280), .Z(n5277) );
  AND U16330 ( .A(a[55]), .B(b[65]), .Z(n5276) );
  XNOR U16331 ( .A(n5281), .B(n4566), .Z(n4568) );
  XOR U16332 ( .A(n5282), .B(n5283), .Z(n4566) );
  ANDN U16333 ( .B(n5284), .A(n5285), .Z(n5282) );
  AND U16334 ( .A(a[56]), .B(b[64]), .Z(n5281) );
  XNOR U16335 ( .A(n5286), .B(n4571), .Z(n4573) );
  XOR U16336 ( .A(n5287), .B(n5288), .Z(n4571) );
  ANDN U16337 ( .B(n5289), .A(n5290), .Z(n5287) );
  AND U16338 ( .A(a[57]), .B(b[63]), .Z(n5286) );
  XNOR U16339 ( .A(n5291), .B(n4576), .Z(n4578) );
  XOR U16340 ( .A(n5292), .B(n5293), .Z(n4576) );
  ANDN U16341 ( .B(n5294), .A(n5295), .Z(n5292) );
  AND U16342 ( .A(a[58]), .B(b[62]), .Z(n5291) );
  XNOR U16343 ( .A(n5296), .B(n4581), .Z(n4583) );
  XOR U16344 ( .A(n5297), .B(n5298), .Z(n4581) );
  ANDN U16345 ( .B(n5299), .A(n5300), .Z(n5297) );
  AND U16346 ( .A(a[59]), .B(b[61]), .Z(n5296) );
  XNOR U16347 ( .A(n5301), .B(n4586), .Z(n4588) );
  XOR U16348 ( .A(n5302), .B(n5303), .Z(n4586) );
  ANDN U16349 ( .B(n5304), .A(n5305), .Z(n5302) );
  AND U16350 ( .A(a[60]), .B(b[60]), .Z(n5301) );
  XNOR U16351 ( .A(n5306), .B(n4591), .Z(n4593) );
  XOR U16352 ( .A(n5307), .B(n5308), .Z(n4591) );
  ANDN U16353 ( .B(n5309), .A(n5310), .Z(n5307) );
  AND U16354 ( .A(a[61]), .B(b[59]), .Z(n5306) );
  XNOR U16355 ( .A(n5311), .B(n4596), .Z(n4598) );
  XOR U16356 ( .A(n5312), .B(n5313), .Z(n4596) );
  ANDN U16357 ( .B(n5314), .A(n5315), .Z(n5312) );
  AND U16358 ( .A(a[62]), .B(b[58]), .Z(n5311) );
  XNOR U16359 ( .A(n5316), .B(n4601), .Z(n4603) );
  XOR U16360 ( .A(n5317), .B(n5318), .Z(n4601) );
  ANDN U16361 ( .B(n5319), .A(n5320), .Z(n5317) );
  AND U16362 ( .A(a[63]), .B(b[57]), .Z(n5316) );
  XNOR U16363 ( .A(n5321), .B(n4606), .Z(n4608) );
  XOR U16364 ( .A(n5322), .B(n5323), .Z(n4606) );
  ANDN U16365 ( .B(n5324), .A(n5325), .Z(n5322) );
  AND U16366 ( .A(a[64]), .B(b[56]), .Z(n5321) );
  XNOR U16367 ( .A(n5326), .B(n4611), .Z(n4613) );
  XOR U16368 ( .A(n5327), .B(n5328), .Z(n4611) );
  ANDN U16369 ( .B(n5329), .A(n5330), .Z(n5327) );
  AND U16370 ( .A(a[65]), .B(b[55]), .Z(n5326) );
  XNOR U16371 ( .A(n5331), .B(n4616), .Z(n4618) );
  XOR U16372 ( .A(n5332), .B(n5333), .Z(n4616) );
  ANDN U16373 ( .B(n5334), .A(n5335), .Z(n5332) );
  AND U16374 ( .A(a[66]), .B(b[54]), .Z(n5331) );
  XNOR U16375 ( .A(n5336), .B(n4621), .Z(n4623) );
  XOR U16376 ( .A(n5337), .B(n5338), .Z(n4621) );
  ANDN U16377 ( .B(n5339), .A(n5340), .Z(n5337) );
  AND U16378 ( .A(a[67]), .B(b[53]), .Z(n5336) );
  XNOR U16379 ( .A(n5341), .B(n4626), .Z(n4628) );
  XOR U16380 ( .A(n5342), .B(n5343), .Z(n4626) );
  ANDN U16381 ( .B(n5344), .A(n5345), .Z(n5342) );
  AND U16382 ( .A(a[68]), .B(b[52]), .Z(n5341) );
  XNOR U16383 ( .A(n5346), .B(n4631), .Z(n4633) );
  XOR U16384 ( .A(n5347), .B(n5348), .Z(n4631) );
  ANDN U16385 ( .B(n5349), .A(n5350), .Z(n5347) );
  AND U16386 ( .A(a[69]), .B(b[51]), .Z(n5346) );
  XNOR U16387 ( .A(n5351), .B(n4636), .Z(n4638) );
  XOR U16388 ( .A(n5352), .B(n5353), .Z(n4636) );
  ANDN U16389 ( .B(n5354), .A(n5355), .Z(n5352) );
  AND U16390 ( .A(a[70]), .B(b[50]), .Z(n5351) );
  XNOR U16391 ( .A(n5356), .B(n4641), .Z(n4643) );
  XOR U16392 ( .A(n5357), .B(n5358), .Z(n4641) );
  ANDN U16393 ( .B(n5359), .A(n5360), .Z(n5357) );
  AND U16394 ( .A(a[71]), .B(b[49]), .Z(n5356) );
  XNOR U16395 ( .A(n5361), .B(n4646), .Z(n4648) );
  XOR U16396 ( .A(n5362), .B(n5363), .Z(n4646) );
  ANDN U16397 ( .B(n5364), .A(n5365), .Z(n5362) );
  AND U16398 ( .A(a[72]), .B(b[48]), .Z(n5361) );
  XNOR U16399 ( .A(n5366), .B(n4651), .Z(n4653) );
  XOR U16400 ( .A(n5367), .B(n5368), .Z(n4651) );
  ANDN U16401 ( .B(n5369), .A(n5370), .Z(n5367) );
  AND U16402 ( .A(a[73]), .B(b[47]), .Z(n5366) );
  XNOR U16403 ( .A(n5371), .B(n4656), .Z(n4658) );
  XOR U16404 ( .A(n5372), .B(n5373), .Z(n4656) );
  ANDN U16405 ( .B(n5374), .A(n5375), .Z(n5372) );
  AND U16406 ( .A(a[74]), .B(b[46]), .Z(n5371) );
  XNOR U16407 ( .A(n5376), .B(n4661), .Z(n4663) );
  XOR U16408 ( .A(n5377), .B(n5378), .Z(n4661) );
  ANDN U16409 ( .B(n5379), .A(n5380), .Z(n5377) );
  AND U16410 ( .A(a[75]), .B(b[45]), .Z(n5376) );
  XNOR U16411 ( .A(n5381), .B(n4666), .Z(n4668) );
  XOR U16412 ( .A(n5382), .B(n5383), .Z(n4666) );
  ANDN U16413 ( .B(n5384), .A(n5385), .Z(n5382) );
  AND U16414 ( .A(a[76]), .B(b[44]), .Z(n5381) );
  XNOR U16415 ( .A(n5386), .B(n4671), .Z(n4673) );
  XOR U16416 ( .A(n5387), .B(n5388), .Z(n4671) );
  ANDN U16417 ( .B(n5389), .A(n5390), .Z(n5387) );
  AND U16418 ( .A(a[77]), .B(b[43]), .Z(n5386) );
  XNOR U16419 ( .A(n5391), .B(n4676), .Z(n4678) );
  XOR U16420 ( .A(n5392), .B(n5393), .Z(n4676) );
  ANDN U16421 ( .B(n5394), .A(n5395), .Z(n5392) );
  AND U16422 ( .A(a[78]), .B(b[42]), .Z(n5391) );
  XNOR U16423 ( .A(n5396), .B(n4681), .Z(n4683) );
  XOR U16424 ( .A(n5397), .B(n5398), .Z(n4681) );
  ANDN U16425 ( .B(n5399), .A(n5400), .Z(n5397) );
  AND U16426 ( .A(a[79]), .B(b[41]), .Z(n5396) );
  XNOR U16427 ( .A(n5401), .B(n4686), .Z(n4688) );
  XOR U16428 ( .A(n5402), .B(n5403), .Z(n4686) );
  ANDN U16429 ( .B(n5404), .A(n5405), .Z(n5402) );
  AND U16430 ( .A(a[80]), .B(b[40]), .Z(n5401) );
  XNOR U16431 ( .A(n5406), .B(n4691), .Z(n4693) );
  XOR U16432 ( .A(n5407), .B(n5408), .Z(n4691) );
  ANDN U16433 ( .B(n5409), .A(n5410), .Z(n5407) );
  AND U16434 ( .A(a[81]), .B(b[39]), .Z(n5406) );
  XNOR U16435 ( .A(n5411), .B(n4696), .Z(n4698) );
  XOR U16436 ( .A(n5412), .B(n5413), .Z(n4696) );
  ANDN U16437 ( .B(n5414), .A(n5415), .Z(n5412) );
  AND U16438 ( .A(a[82]), .B(b[38]), .Z(n5411) );
  XNOR U16439 ( .A(n5416), .B(n4701), .Z(n4703) );
  XOR U16440 ( .A(n5417), .B(n5418), .Z(n4701) );
  ANDN U16441 ( .B(n5419), .A(n5420), .Z(n5417) );
  AND U16442 ( .A(a[83]), .B(b[37]), .Z(n5416) );
  XNOR U16443 ( .A(n5421), .B(n4706), .Z(n4708) );
  XOR U16444 ( .A(n5422), .B(n5423), .Z(n4706) );
  ANDN U16445 ( .B(n5424), .A(n5425), .Z(n5422) );
  AND U16446 ( .A(a[84]), .B(b[36]), .Z(n5421) );
  XNOR U16447 ( .A(n5426), .B(n4711), .Z(n4713) );
  XOR U16448 ( .A(n5427), .B(n5428), .Z(n4711) );
  ANDN U16449 ( .B(n5429), .A(n5430), .Z(n5427) );
  AND U16450 ( .A(a[85]), .B(b[35]), .Z(n5426) );
  XNOR U16451 ( .A(n5431), .B(n4716), .Z(n4718) );
  XOR U16452 ( .A(n5432), .B(n5433), .Z(n4716) );
  ANDN U16453 ( .B(n5434), .A(n5435), .Z(n5432) );
  AND U16454 ( .A(a[86]), .B(b[34]), .Z(n5431) );
  XNOR U16455 ( .A(n5436), .B(n4721), .Z(n4723) );
  XOR U16456 ( .A(n5437), .B(n5438), .Z(n4721) );
  ANDN U16457 ( .B(n5439), .A(n5440), .Z(n5437) );
  AND U16458 ( .A(a[87]), .B(b[33]), .Z(n5436) );
  XNOR U16459 ( .A(n5441), .B(n4726), .Z(n4728) );
  XOR U16460 ( .A(n5442), .B(n5443), .Z(n4726) );
  ANDN U16461 ( .B(n5444), .A(n5445), .Z(n5442) );
  AND U16462 ( .A(a[88]), .B(b[32]), .Z(n5441) );
  XNOR U16463 ( .A(n5446), .B(n4731), .Z(n4733) );
  XOR U16464 ( .A(n5447), .B(n5448), .Z(n4731) );
  ANDN U16465 ( .B(n5449), .A(n5450), .Z(n5447) );
  AND U16466 ( .A(a[89]), .B(b[31]), .Z(n5446) );
  XNOR U16467 ( .A(n5451), .B(n4736), .Z(n4738) );
  XOR U16468 ( .A(n5452), .B(n5453), .Z(n4736) );
  ANDN U16469 ( .B(n5454), .A(n5455), .Z(n5452) );
  AND U16470 ( .A(a[90]), .B(b[30]), .Z(n5451) );
  XNOR U16471 ( .A(n5456), .B(n4741), .Z(n4743) );
  XOR U16472 ( .A(n5457), .B(n5458), .Z(n4741) );
  ANDN U16473 ( .B(n5459), .A(n5460), .Z(n5457) );
  AND U16474 ( .A(a[91]), .B(b[29]), .Z(n5456) );
  XNOR U16475 ( .A(n5461), .B(n4746), .Z(n4748) );
  XOR U16476 ( .A(n5462), .B(n5463), .Z(n4746) );
  ANDN U16477 ( .B(n5464), .A(n5465), .Z(n5462) );
  AND U16478 ( .A(a[92]), .B(b[28]), .Z(n5461) );
  XNOR U16479 ( .A(n5466), .B(n4751), .Z(n4753) );
  XOR U16480 ( .A(n5467), .B(n5468), .Z(n4751) );
  ANDN U16481 ( .B(n5469), .A(n5470), .Z(n5467) );
  AND U16482 ( .A(a[93]), .B(b[27]), .Z(n5466) );
  XNOR U16483 ( .A(n5471), .B(n4756), .Z(n4758) );
  XOR U16484 ( .A(n5472), .B(n5473), .Z(n4756) );
  ANDN U16485 ( .B(n5474), .A(n5475), .Z(n5472) );
  AND U16486 ( .A(a[94]), .B(b[26]), .Z(n5471) );
  XNOR U16487 ( .A(n5476), .B(n4761), .Z(n4763) );
  XOR U16488 ( .A(n5477), .B(n5478), .Z(n4761) );
  ANDN U16489 ( .B(n5479), .A(n5480), .Z(n5477) );
  AND U16490 ( .A(a[95]), .B(b[25]), .Z(n5476) );
  XNOR U16491 ( .A(n5481), .B(n4766), .Z(n4768) );
  XOR U16492 ( .A(n5482), .B(n5483), .Z(n4766) );
  ANDN U16493 ( .B(n5484), .A(n5485), .Z(n5482) );
  AND U16494 ( .A(a[96]), .B(b[24]), .Z(n5481) );
  XNOR U16495 ( .A(n5486), .B(n4771), .Z(n4773) );
  XOR U16496 ( .A(n5487), .B(n5488), .Z(n4771) );
  ANDN U16497 ( .B(n5489), .A(n5490), .Z(n5487) );
  AND U16498 ( .A(a[97]), .B(b[23]), .Z(n5486) );
  XNOR U16499 ( .A(n5491), .B(n4776), .Z(n4778) );
  XOR U16500 ( .A(n5492), .B(n5493), .Z(n4776) );
  ANDN U16501 ( .B(n5494), .A(n5495), .Z(n5492) );
  AND U16502 ( .A(a[98]), .B(b[22]), .Z(n5491) );
  XNOR U16503 ( .A(n5496), .B(n4781), .Z(n4783) );
  XOR U16504 ( .A(n5497), .B(n5498), .Z(n4781) );
  ANDN U16505 ( .B(n5499), .A(n5500), .Z(n5497) );
  AND U16506 ( .A(a[99]), .B(b[21]), .Z(n5496) );
  XNOR U16507 ( .A(n5501), .B(n4786), .Z(n4788) );
  XOR U16508 ( .A(n5502), .B(n5503), .Z(n4786) );
  ANDN U16509 ( .B(n5504), .A(n5505), .Z(n5502) );
  AND U16510 ( .A(b[20]), .B(a[100]), .Z(n5501) );
  XNOR U16511 ( .A(n5506), .B(n4791), .Z(n4793) );
  XOR U16512 ( .A(n5507), .B(n5508), .Z(n4791) );
  ANDN U16513 ( .B(n5509), .A(n5510), .Z(n5507) );
  AND U16514 ( .A(b[19]), .B(a[101]), .Z(n5506) );
  XNOR U16515 ( .A(n5511), .B(n4796), .Z(n4798) );
  XOR U16516 ( .A(n5512), .B(n5513), .Z(n4796) );
  ANDN U16517 ( .B(n5514), .A(n5515), .Z(n5512) );
  AND U16518 ( .A(b[18]), .B(a[102]), .Z(n5511) );
  XNOR U16519 ( .A(n5516), .B(n4801), .Z(n4803) );
  XOR U16520 ( .A(n5517), .B(n5518), .Z(n4801) );
  ANDN U16521 ( .B(n5519), .A(n5520), .Z(n5517) );
  AND U16522 ( .A(b[17]), .B(a[103]), .Z(n5516) );
  XNOR U16523 ( .A(n5521), .B(n4806), .Z(n4808) );
  XOR U16524 ( .A(n5522), .B(n5523), .Z(n4806) );
  ANDN U16525 ( .B(n5524), .A(n5525), .Z(n5522) );
  AND U16526 ( .A(b[16]), .B(a[104]), .Z(n5521) );
  XNOR U16527 ( .A(n5526), .B(n4811), .Z(n4813) );
  XOR U16528 ( .A(n5527), .B(n5528), .Z(n4811) );
  ANDN U16529 ( .B(n5529), .A(n5530), .Z(n5527) );
  AND U16530 ( .A(b[15]), .B(a[105]), .Z(n5526) );
  XNOR U16531 ( .A(n5531), .B(n4816), .Z(n4818) );
  XOR U16532 ( .A(n5532), .B(n5533), .Z(n4816) );
  ANDN U16533 ( .B(n5534), .A(n5535), .Z(n5532) );
  AND U16534 ( .A(b[14]), .B(a[106]), .Z(n5531) );
  XNOR U16535 ( .A(n5536), .B(n4821), .Z(n4823) );
  XOR U16536 ( .A(n5537), .B(n5538), .Z(n4821) );
  ANDN U16537 ( .B(n5539), .A(n5540), .Z(n5537) );
  AND U16538 ( .A(b[13]), .B(a[107]), .Z(n5536) );
  XNOR U16539 ( .A(n5541), .B(n4826), .Z(n4828) );
  XOR U16540 ( .A(n5542), .B(n5543), .Z(n4826) );
  ANDN U16541 ( .B(n5544), .A(n5545), .Z(n5542) );
  AND U16542 ( .A(b[12]), .B(a[108]), .Z(n5541) );
  XNOR U16543 ( .A(n5546), .B(n4831), .Z(n4833) );
  XOR U16544 ( .A(n5547), .B(n5548), .Z(n4831) );
  ANDN U16545 ( .B(n5549), .A(n5550), .Z(n5547) );
  AND U16546 ( .A(b[11]), .B(a[109]), .Z(n5546) );
  XNOR U16547 ( .A(n5551), .B(n4836), .Z(n4838) );
  XOR U16548 ( .A(n5552), .B(n5553), .Z(n4836) );
  ANDN U16549 ( .B(n5554), .A(n5555), .Z(n5552) );
  AND U16550 ( .A(b[10]), .B(a[110]), .Z(n5551) );
  XNOR U16551 ( .A(n5556), .B(n4841), .Z(n4843) );
  XOR U16552 ( .A(n5557), .B(n5558), .Z(n4841) );
  ANDN U16553 ( .B(n5559), .A(n5560), .Z(n5557) );
  AND U16554 ( .A(b[9]), .B(a[111]), .Z(n5556) );
  XNOR U16555 ( .A(n5561), .B(n4846), .Z(n4848) );
  XOR U16556 ( .A(n5562), .B(n5563), .Z(n4846) );
  ANDN U16557 ( .B(n5564), .A(n5565), .Z(n5562) );
  AND U16558 ( .A(b[8]), .B(a[112]), .Z(n5561) );
  XNOR U16559 ( .A(n5566), .B(n4851), .Z(n4853) );
  XOR U16560 ( .A(n5567), .B(n5568), .Z(n4851) );
  ANDN U16561 ( .B(n5569), .A(n5570), .Z(n5567) );
  AND U16562 ( .A(b[7]), .B(a[113]), .Z(n5566) );
  XNOR U16563 ( .A(n5571), .B(n4856), .Z(n4858) );
  XOR U16564 ( .A(n5572), .B(n5573), .Z(n4856) );
  ANDN U16565 ( .B(n5574), .A(n5575), .Z(n5572) );
  AND U16566 ( .A(b[6]), .B(a[114]), .Z(n5571) );
  XNOR U16567 ( .A(n5576), .B(n4861), .Z(n4863) );
  XOR U16568 ( .A(n5577), .B(n5578), .Z(n4861) );
  ANDN U16569 ( .B(n5579), .A(n5580), .Z(n5577) );
  AND U16570 ( .A(b[5]), .B(a[115]), .Z(n5576) );
  XNOR U16571 ( .A(n5581), .B(n4866), .Z(n4868) );
  XOR U16572 ( .A(n5582), .B(n5583), .Z(n4866) );
  ANDN U16573 ( .B(n5584), .A(n5585), .Z(n5582) );
  AND U16574 ( .A(b[4]), .B(a[116]), .Z(n5581) );
  XNOR U16575 ( .A(n5586), .B(n5587), .Z(n4880) );
  NANDN U16576 ( .A(n5588), .B(n5589), .Z(n5587) );
  XNOR U16577 ( .A(n5590), .B(n4871), .Z(n4873) );
  XNOR U16578 ( .A(n5591), .B(n5592), .Z(n4871) );
  AND U16579 ( .A(n5593), .B(n5594), .Z(n5591) );
  AND U16580 ( .A(b[3]), .B(a[117]), .Z(n5590) );
  NAND U16581 ( .A(a[120]), .B(b[0]), .Z(n4168) );
  XNOR U16582 ( .A(n5595), .B(n5596), .Z(c[11]) );
  XNOR U16583 ( .A(n4886), .B(n4887), .Z(c[119]) );
  XNOR U16584 ( .A(n5588), .B(n5589), .Z(n4887) );
  XOR U16585 ( .A(n5586), .B(n5597), .Z(n5589) );
  NAND U16586 ( .A(b[1]), .B(a[118]), .Z(n5597) );
  XOR U16587 ( .A(n5594), .B(n5598), .Z(n5588) );
  XOR U16588 ( .A(n5586), .B(n5593), .Z(n5598) );
  XNOR U16589 ( .A(n5599), .B(n5592), .Z(n5593) );
  AND U16590 ( .A(b[2]), .B(a[117]), .Z(n5599) );
  NANDN U16591 ( .A(n5600), .B(n5601), .Z(n5586) );
  XOR U16592 ( .A(n5592), .B(n5584), .Z(n5602) );
  XNOR U16593 ( .A(n5583), .B(n5579), .Z(n5603) );
  XNOR U16594 ( .A(n5578), .B(n5574), .Z(n5604) );
  XNOR U16595 ( .A(n5573), .B(n5569), .Z(n5605) );
  XNOR U16596 ( .A(n5568), .B(n5564), .Z(n5606) );
  XNOR U16597 ( .A(n5563), .B(n5559), .Z(n5607) );
  XNOR U16598 ( .A(n5558), .B(n5554), .Z(n5608) );
  XNOR U16599 ( .A(n5553), .B(n5549), .Z(n5609) );
  XNOR U16600 ( .A(n5548), .B(n5544), .Z(n5610) );
  XNOR U16601 ( .A(n5543), .B(n5539), .Z(n5611) );
  XNOR U16602 ( .A(n5538), .B(n5534), .Z(n5612) );
  XNOR U16603 ( .A(n5533), .B(n5529), .Z(n5613) );
  XNOR U16604 ( .A(n5528), .B(n5524), .Z(n5614) );
  XNOR U16605 ( .A(n5523), .B(n5519), .Z(n5615) );
  XNOR U16606 ( .A(n5518), .B(n5514), .Z(n5616) );
  XNOR U16607 ( .A(n5513), .B(n5509), .Z(n5617) );
  XNOR U16608 ( .A(n5508), .B(n5504), .Z(n5618) );
  XNOR U16609 ( .A(n5503), .B(n5499), .Z(n5619) );
  XNOR U16610 ( .A(n5498), .B(n5494), .Z(n5620) );
  XNOR U16611 ( .A(n5493), .B(n5489), .Z(n5621) );
  XNOR U16612 ( .A(n5488), .B(n5484), .Z(n5622) );
  XNOR U16613 ( .A(n5483), .B(n5479), .Z(n5623) );
  XNOR U16614 ( .A(n5478), .B(n5474), .Z(n5624) );
  XNOR U16615 ( .A(n5473), .B(n5469), .Z(n5625) );
  XNOR U16616 ( .A(n5468), .B(n5464), .Z(n5626) );
  XNOR U16617 ( .A(n5463), .B(n5459), .Z(n5627) );
  XNOR U16618 ( .A(n5458), .B(n5454), .Z(n5628) );
  XNOR U16619 ( .A(n5453), .B(n5449), .Z(n5629) );
  XNOR U16620 ( .A(n5448), .B(n5444), .Z(n5630) );
  XNOR U16621 ( .A(n5443), .B(n5439), .Z(n5631) );
  XNOR U16622 ( .A(n5438), .B(n5434), .Z(n5632) );
  XNOR U16623 ( .A(n5433), .B(n5429), .Z(n5633) );
  XNOR U16624 ( .A(n5428), .B(n5424), .Z(n5634) );
  XNOR U16625 ( .A(n5423), .B(n5419), .Z(n5635) );
  XNOR U16626 ( .A(n5418), .B(n5414), .Z(n5636) );
  XNOR U16627 ( .A(n5413), .B(n5409), .Z(n5637) );
  XNOR U16628 ( .A(n5408), .B(n5404), .Z(n5638) );
  XNOR U16629 ( .A(n5403), .B(n5399), .Z(n5639) );
  XNOR U16630 ( .A(n5398), .B(n5394), .Z(n5640) );
  XNOR U16631 ( .A(n5393), .B(n5389), .Z(n5641) );
  XNOR U16632 ( .A(n5388), .B(n5384), .Z(n5642) );
  XNOR U16633 ( .A(n5383), .B(n5379), .Z(n5643) );
  XNOR U16634 ( .A(n5378), .B(n5374), .Z(n5644) );
  XNOR U16635 ( .A(n5373), .B(n5369), .Z(n5645) );
  XNOR U16636 ( .A(n5368), .B(n5364), .Z(n5646) );
  XNOR U16637 ( .A(n5363), .B(n5359), .Z(n5647) );
  XNOR U16638 ( .A(n5358), .B(n5354), .Z(n5648) );
  XNOR U16639 ( .A(n5353), .B(n5349), .Z(n5649) );
  XNOR U16640 ( .A(n5348), .B(n5344), .Z(n5650) );
  XNOR U16641 ( .A(n5343), .B(n5339), .Z(n5651) );
  XNOR U16642 ( .A(n5338), .B(n5334), .Z(n5652) );
  XNOR U16643 ( .A(n5333), .B(n5329), .Z(n5653) );
  XNOR U16644 ( .A(n5328), .B(n5324), .Z(n5654) );
  XNOR U16645 ( .A(n5323), .B(n5319), .Z(n5655) );
  XNOR U16646 ( .A(n5318), .B(n5314), .Z(n5656) );
  XNOR U16647 ( .A(n5313), .B(n5309), .Z(n5657) );
  XNOR U16648 ( .A(n5308), .B(n5304), .Z(n5658) );
  XNOR U16649 ( .A(n5303), .B(n5299), .Z(n5659) );
  XNOR U16650 ( .A(n5298), .B(n5294), .Z(n5660) );
  XNOR U16651 ( .A(n5293), .B(n5289), .Z(n5661) );
  XNOR U16652 ( .A(n5288), .B(n5284), .Z(n5662) );
  XNOR U16653 ( .A(n5283), .B(n5279), .Z(n5663) );
  XNOR U16654 ( .A(n5278), .B(n5274), .Z(n5664) );
  XNOR U16655 ( .A(n5273), .B(n5269), .Z(n5665) );
  XNOR U16656 ( .A(n5268), .B(n5264), .Z(n5666) );
  XNOR U16657 ( .A(n5263), .B(n5259), .Z(n5667) );
  XNOR U16658 ( .A(n5258), .B(n5254), .Z(n5668) );
  XNOR U16659 ( .A(n5253), .B(n5249), .Z(n5669) );
  XNOR U16660 ( .A(n5248), .B(n5244), .Z(n5670) );
  XNOR U16661 ( .A(n5243), .B(n5239), .Z(n5671) );
  XNOR U16662 ( .A(n5238), .B(n5234), .Z(n5672) );
  XNOR U16663 ( .A(n5233), .B(n5229), .Z(n5673) );
  XNOR U16664 ( .A(n5228), .B(n5224), .Z(n5674) );
  XNOR U16665 ( .A(n5223), .B(n5219), .Z(n5675) );
  XNOR U16666 ( .A(n5218), .B(n5214), .Z(n5676) );
  XNOR U16667 ( .A(n5213), .B(n5209), .Z(n5677) );
  XNOR U16668 ( .A(n5208), .B(n5204), .Z(n5678) );
  XNOR U16669 ( .A(n5203), .B(n5199), .Z(n5679) );
  XNOR U16670 ( .A(n5198), .B(n5194), .Z(n5680) );
  XNOR U16671 ( .A(n5193), .B(n5189), .Z(n5681) );
  XNOR U16672 ( .A(n5188), .B(n5184), .Z(n5682) );
  XNOR U16673 ( .A(n5183), .B(n5179), .Z(n5683) );
  XNOR U16674 ( .A(n5178), .B(n5174), .Z(n5684) );
  XNOR U16675 ( .A(n5173), .B(n5169), .Z(n5685) );
  XNOR U16676 ( .A(n5168), .B(n5164), .Z(n5686) );
  XNOR U16677 ( .A(n5163), .B(n5159), .Z(n5687) );
  XNOR U16678 ( .A(n5158), .B(n5154), .Z(n5688) );
  XNOR U16679 ( .A(n5153), .B(n5149), .Z(n5689) );
  XNOR U16680 ( .A(n5148), .B(n5144), .Z(n5690) );
  XNOR U16681 ( .A(n5143), .B(n5139), .Z(n5691) );
  XNOR U16682 ( .A(n5138), .B(n5134), .Z(n5692) );
  XNOR U16683 ( .A(n5133), .B(n5129), .Z(n5693) );
  XNOR U16684 ( .A(n5128), .B(n5124), .Z(n5694) );
  XNOR U16685 ( .A(n5123), .B(n5119), .Z(n5695) );
  XNOR U16686 ( .A(n5118), .B(n5114), .Z(n5696) );
  XNOR U16687 ( .A(n5113), .B(n5109), .Z(n5697) );
  XNOR U16688 ( .A(n5108), .B(n5104), .Z(n5698) );
  XNOR U16689 ( .A(n5103), .B(n5099), .Z(n5699) );
  XNOR U16690 ( .A(n5098), .B(n5094), .Z(n5700) );
  XNOR U16691 ( .A(n5093), .B(n5089), .Z(n5701) );
  XNOR U16692 ( .A(n5088), .B(n5084), .Z(n5702) );
  XNOR U16693 ( .A(n5083), .B(n5079), .Z(n5703) );
  XNOR U16694 ( .A(n5078), .B(n5074), .Z(n5704) );
  XNOR U16695 ( .A(n5073), .B(n5069), .Z(n5705) );
  XNOR U16696 ( .A(n5068), .B(n5064), .Z(n5706) );
  XNOR U16697 ( .A(n5063), .B(n5059), .Z(n5707) );
  XNOR U16698 ( .A(n5058), .B(n5054), .Z(n5708) );
  XNOR U16699 ( .A(n5053), .B(n5049), .Z(n5709) );
  XNOR U16700 ( .A(n5048), .B(n5044), .Z(n5710) );
  XNOR U16701 ( .A(n5043), .B(n5039), .Z(n5711) );
  XNOR U16702 ( .A(n5038), .B(n5034), .Z(n5712) );
  XNOR U16703 ( .A(n5033), .B(n5029), .Z(n5713) );
  XNOR U16704 ( .A(n5028), .B(n5024), .Z(n5714) );
  XNOR U16705 ( .A(n5023), .B(n5019), .Z(n5715) );
  XNOR U16706 ( .A(n5018), .B(n5014), .Z(n5716) );
  XNOR U16707 ( .A(n5013), .B(n5009), .Z(n5717) );
  XNOR U16708 ( .A(n5718), .B(n5008), .Z(n5009) );
  AND U16709 ( .A(a[0]), .B(b[119]), .Z(n5718) );
  XOR U16710 ( .A(n5719), .B(n5008), .Z(n5010) );
  XNOR U16711 ( .A(n5720), .B(n5721), .Z(n5008) );
  ANDN U16712 ( .B(n5722), .A(n5723), .Z(n5720) );
  AND U16713 ( .A(a[1]), .B(b[118]), .Z(n5719) );
  XNOR U16714 ( .A(n5724), .B(n5013), .Z(n5015) );
  XOR U16715 ( .A(n5725), .B(n5726), .Z(n5013) );
  ANDN U16716 ( .B(n5727), .A(n5728), .Z(n5725) );
  AND U16717 ( .A(a[2]), .B(b[117]), .Z(n5724) );
  XNOR U16718 ( .A(n5729), .B(n5018), .Z(n5020) );
  XOR U16719 ( .A(n5730), .B(n5731), .Z(n5018) );
  ANDN U16720 ( .B(n5732), .A(n5733), .Z(n5730) );
  AND U16721 ( .A(a[3]), .B(b[116]), .Z(n5729) );
  XNOR U16722 ( .A(n5734), .B(n5023), .Z(n5025) );
  XOR U16723 ( .A(n5735), .B(n5736), .Z(n5023) );
  ANDN U16724 ( .B(n5737), .A(n5738), .Z(n5735) );
  AND U16725 ( .A(a[4]), .B(b[115]), .Z(n5734) );
  XNOR U16726 ( .A(n5739), .B(n5028), .Z(n5030) );
  XOR U16727 ( .A(n5740), .B(n5741), .Z(n5028) );
  ANDN U16728 ( .B(n5742), .A(n5743), .Z(n5740) );
  AND U16729 ( .A(a[5]), .B(b[114]), .Z(n5739) );
  XNOR U16730 ( .A(n5744), .B(n5033), .Z(n5035) );
  XOR U16731 ( .A(n5745), .B(n5746), .Z(n5033) );
  ANDN U16732 ( .B(n5747), .A(n5748), .Z(n5745) );
  AND U16733 ( .A(a[6]), .B(b[113]), .Z(n5744) );
  XNOR U16734 ( .A(n5749), .B(n5038), .Z(n5040) );
  XOR U16735 ( .A(n5750), .B(n5751), .Z(n5038) );
  ANDN U16736 ( .B(n5752), .A(n5753), .Z(n5750) );
  AND U16737 ( .A(a[7]), .B(b[112]), .Z(n5749) );
  XNOR U16738 ( .A(n5754), .B(n5043), .Z(n5045) );
  XOR U16739 ( .A(n5755), .B(n5756), .Z(n5043) );
  ANDN U16740 ( .B(n5757), .A(n5758), .Z(n5755) );
  AND U16741 ( .A(a[8]), .B(b[111]), .Z(n5754) );
  XNOR U16742 ( .A(n5759), .B(n5048), .Z(n5050) );
  XOR U16743 ( .A(n5760), .B(n5761), .Z(n5048) );
  ANDN U16744 ( .B(n5762), .A(n5763), .Z(n5760) );
  AND U16745 ( .A(a[9]), .B(b[110]), .Z(n5759) );
  XNOR U16746 ( .A(n5764), .B(n5053), .Z(n5055) );
  XOR U16747 ( .A(n5765), .B(n5766), .Z(n5053) );
  ANDN U16748 ( .B(n5767), .A(n5768), .Z(n5765) );
  AND U16749 ( .A(a[10]), .B(b[109]), .Z(n5764) );
  XNOR U16750 ( .A(n5769), .B(n5058), .Z(n5060) );
  XOR U16751 ( .A(n5770), .B(n5771), .Z(n5058) );
  ANDN U16752 ( .B(n5772), .A(n5773), .Z(n5770) );
  AND U16753 ( .A(a[11]), .B(b[108]), .Z(n5769) );
  XNOR U16754 ( .A(n5774), .B(n5063), .Z(n5065) );
  XOR U16755 ( .A(n5775), .B(n5776), .Z(n5063) );
  ANDN U16756 ( .B(n5777), .A(n5778), .Z(n5775) );
  AND U16757 ( .A(a[12]), .B(b[107]), .Z(n5774) );
  XNOR U16758 ( .A(n5779), .B(n5068), .Z(n5070) );
  XOR U16759 ( .A(n5780), .B(n5781), .Z(n5068) );
  ANDN U16760 ( .B(n5782), .A(n5783), .Z(n5780) );
  AND U16761 ( .A(a[13]), .B(b[106]), .Z(n5779) );
  XNOR U16762 ( .A(n5784), .B(n5073), .Z(n5075) );
  XOR U16763 ( .A(n5785), .B(n5786), .Z(n5073) );
  ANDN U16764 ( .B(n5787), .A(n5788), .Z(n5785) );
  AND U16765 ( .A(a[14]), .B(b[105]), .Z(n5784) );
  XNOR U16766 ( .A(n5789), .B(n5078), .Z(n5080) );
  XOR U16767 ( .A(n5790), .B(n5791), .Z(n5078) );
  ANDN U16768 ( .B(n5792), .A(n5793), .Z(n5790) );
  AND U16769 ( .A(a[15]), .B(b[104]), .Z(n5789) );
  XNOR U16770 ( .A(n5794), .B(n5083), .Z(n5085) );
  XOR U16771 ( .A(n5795), .B(n5796), .Z(n5083) );
  ANDN U16772 ( .B(n5797), .A(n5798), .Z(n5795) );
  AND U16773 ( .A(a[16]), .B(b[103]), .Z(n5794) );
  XNOR U16774 ( .A(n5799), .B(n5088), .Z(n5090) );
  XOR U16775 ( .A(n5800), .B(n5801), .Z(n5088) );
  ANDN U16776 ( .B(n5802), .A(n5803), .Z(n5800) );
  AND U16777 ( .A(a[17]), .B(b[102]), .Z(n5799) );
  XNOR U16778 ( .A(n5804), .B(n5093), .Z(n5095) );
  XOR U16779 ( .A(n5805), .B(n5806), .Z(n5093) );
  ANDN U16780 ( .B(n5807), .A(n5808), .Z(n5805) );
  AND U16781 ( .A(a[18]), .B(b[101]), .Z(n5804) );
  XNOR U16782 ( .A(n5809), .B(n5098), .Z(n5100) );
  XOR U16783 ( .A(n5810), .B(n5811), .Z(n5098) );
  ANDN U16784 ( .B(n5812), .A(n5813), .Z(n5810) );
  AND U16785 ( .A(a[19]), .B(b[100]), .Z(n5809) );
  XNOR U16786 ( .A(n5814), .B(n5103), .Z(n5105) );
  XOR U16787 ( .A(n5815), .B(n5816), .Z(n5103) );
  ANDN U16788 ( .B(n5817), .A(n5818), .Z(n5815) );
  AND U16789 ( .A(a[20]), .B(b[99]), .Z(n5814) );
  XNOR U16790 ( .A(n5819), .B(n5108), .Z(n5110) );
  XOR U16791 ( .A(n5820), .B(n5821), .Z(n5108) );
  ANDN U16792 ( .B(n5822), .A(n5823), .Z(n5820) );
  AND U16793 ( .A(a[21]), .B(b[98]), .Z(n5819) );
  XNOR U16794 ( .A(n5824), .B(n5113), .Z(n5115) );
  XOR U16795 ( .A(n5825), .B(n5826), .Z(n5113) );
  ANDN U16796 ( .B(n5827), .A(n5828), .Z(n5825) );
  AND U16797 ( .A(a[22]), .B(b[97]), .Z(n5824) );
  XNOR U16798 ( .A(n5829), .B(n5118), .Z(n5120) );
  XOR U16799 ( .A(n5830), .B(n5831), .Z(n5118) );
  ANDN U16800 ( .B(n5832), .A(n5833), .Z(n5830) );
  AND U16801 ( .A(a[23]), .B(b[96]), .Z(n5829) );
  XNOR U16802 ( .A(n5834), .B(n5123), .Z(n5125) );
  XOR U16803 ( .A(n5835), .B(n5836), .Z(n5123) );
  ANDN U16804 ( .B(n5837), .A(n5838), .Z(n5835) );
  AND U16805 ( .A(a[24]), .B(b[95]), .Z(n5834) );
  XNOR U16806 ( .A(n5839), .B(n5128), .Z(n5130) );
  XOR U16807 ( .A(n5840), .B(n5841), .Z(n5128) );
  ANDN U16808 ( .B(n5842), .A(n5843), .Z(n5840) );
  AND U16809 ( .A(a[25]), .B(b[94]), .Z(n5839) );
  XNOR U16810 ( .A(n5844), .B(n5133), .Z(n5135) );
  XOR U16811 ( .A(n5845), .B(n5846), .Z(n5133) );
  ANDN U16812 ( .B(n5847), .A(n5848), .Z(n5845) );
  AND U16813 ( .A(a[26]), .B(b[93]), .Z(n5844) );
  XNOR U16814 ( .A(n5849), .B(n5138), .Z(n5140) );
  XOR U16815 ( .A(n5850), .B(n5851), .Z(n5138) );
  ANDN U16816 ( .B(n5852), .A(n5853), .Z(n5850) );
  AND U16817 ( .A(a[27]), .B(b[92]), .Z(n5849) );
  XNOR U16818 ( .A(n5854), .B(n5143), .Z(n5145) );
  XOR U16819 ( .A(n5855), .B(n5856), .Z(n5143) );
  ANDN U16820 ( .B(n5857), .A(n5858), .Z(n5855) );
  AND U16821 ( .A(a[28]), .B(b[91]), .Z(n5854) );
  XNOR U16822 ( .A(n5859), .B(n5148), .Z(n5150) );
  XOR U16823 ( .A(n5860), .B(n5861), .Z(n5148) );
  ANDN U16824 ( .B(n5862), .A(n5863), .Z(n5860) );
  AND U16825 ( .A(a[29]), .B(b[90]), .Z(n5859) );
  XNOR U16826 ( .A(n5864), .B(n5153), .Z(n5155) );
  XOR U16827 ( .A(n5865), .B(n5866), .Z(n5153) );
  ANDN U16828 ( .B(n5867), .A(n5868), .Z(n5865) );
  AND U16829 ( .A(a[30]), .B(b[89]), .Z(n5864) );
  XNOR U16830 ( .A(n5869), .B(n5158), .Z(n5160) );
  XOR U16831 ( .A(n5870), .B(n5871), .Z(n5158) );
  ANDN U16832 ( .B(n5872), .A(n5873), .Z(n5870) );
  AND U16833 ( .A(a[31]), .B(b[88]), .Z(n5869) );
  XNOR U16834 ( .A(n5874), .B(n5163), .Z(n5165) );
  XOR U16835 ( .A(n5875), .B(n5876), .Z(n5163) );
  ANDN U16836 ( .B(n5877), .A(n5878), .Z(n5875) );
  AND U16837 ( .A(a[32]), .B(b[87]), .Z(n5874) );
  XNOR U16838 ( .A(n5879), .B(n5168), .Z(n5170) );
  XOR U16839 ( .A(n5880), .B(n5881), .Z(n5168) );
  ANDN U16840 ( .B(n5882), .A(n5883), .Z(n5880) );
  AND U16841 ( .A(a[33]), .B(b[86]), .Z(n5879) );
  XNOR U16842 ( .A(n5884), .B(n5173), .Z(n5175) );
  XOR U16843 ( .A(n5885), .B(n5886), .Z(n5173) );
  ANDN U16844 ( .B(n5887), .A(n5888), .Z(n5885) );
  AND U16845 ( .A(a[34]), .B(b[85]), .Z(n5884) );
  XNOR U16846 ( .A(n5889), .B(n5178), .Z(n5180) );
  XOR U16847 ( .A(n5890), .B(n5891), .Z(n5178) );
  ANDN U16848 ( .B(n5892), .A(n5893), .Z(n5890) );
  AND U16849 ( .A(a[35]), .B(b[84]), .Z(n5889) );
  XNOR U16850 ( .A(n5894), .B(n5183), .Z(n5185) );
  XOR U16851 ( .A(n5895), .B(n5896), .Z(n5183) );
  ANDN U16852 ( .B(n5897), .A(n5898), .Z(n5895) );
  AND U16853 ( .A(a[36]), .B(b[83]), .Z(n5894) );
  XNOR U16854 ( .A(n5899), .B(n5188), .Z(n5190) );
  XOR U16855 ( .A(n5900), .B(n5901), .Z(n5188) );
  ANDN U16856 ( .B(n5902), .A(n5903), .Z(n5900) );
  AND U16857 ( .A(a[37]), .B(b[82]), .Z(n5899) );
  XNOR U16858 ( .A(n5904), .B(n5193), .Z(n5195) );
  XOR U16859 ( .A(n5905), .B(n5906), .Z(n5193) );
  ANDN U16860 ( .B(n5907), .A(n5908), .Z(n5905) );
  AND U16861 ( .A(a[38]), .B(b[81]), .Z(n5904) );
  XNOR U16862 ( .A(n5909), .B(n5198), .Z(n5200) );
  XOR U16863 ( .A(n5910), .B(n5911), .Z(n5198) );
  ANDN U16864 ( .B(n5912), .A(n5913), .Z(n5910) );
  AND U16865 ( .A(a[39]), .B(b[80]), .Z(n5909) );
  XNOR U16866 ( .A(n5914), .B(n5203), .Z(n5205) );
  XOR U16867 ( .A(n5915), .B(n5916), .Z(n5203) );
  ANDN U16868 ( .B(n5917), .A(n5918), .Z(n5915) );
  AND U16869 ( .A(a[40]), .B(b[79]), .Z(n5914) );
  XNOR U16870 ( .A(n5919), .B(n5208), .Z(n5210) );
  XOR U16871 ( .A(n5920), .B(n5921), .Z(n5208) );
  ANDN U16872 ( .B(n5922), .A(n5923), .Z(n5920) );
  AND U16873 ( .A(a[41]), .B(b[78]), .Z(n5919) );
  XNOR U16874 ( .A(n5924), .B(n5213), .Z(n5215) );
  XOR U16875 ( .A(n5925), .B(n5926), .Z(n5213) );
  ANDN U16876 ( .B(n5927), .A(n5928), .Z(n5925) );
  AND U16877 ( .A(a[42]), .B(b[77]), .Z(n5924) );
  XNOR U16878 ( .A(n5929), .B(n5218), .Z(n5220) );
  XOR U16879 ( .A(n5930), .B(n5931), .Z(n5218) );
  ANDN U16880 ( .B(n5932), .A(n5933), .Z(n5930) );
  AND U16881 ( .A(a[43]), .B(b[76]), .Z(n5929) );
  XNOR U16882 ( .A(n5934), .B(n5223), .Z(n5225) );
  XOR U16883 ( .A(n5935), .B(n5936), .Z(n5223) );
  ANDN U16884 ( .B(n5937), .A(n5938), .Z(n5935) );
  AND U16885 ( .A(a[44]), .B(b[75]), .Z(n5934) );
  XNOR U16886 ( .A(n5939), .B(n5228), .Z(n5230) );
  XOR U16887 ( .A(n5940), .B(n5941), .Z(n5228) );
  ANDN U16888 ( .B(n5942), .A(n5943), .Z(n5940) );
  AND U16889 ( .A(a[45]), .B(b[74]), .Z(n5939) );
  XNOR U16890 ( .A(n5944), .B(n5233), .Z(n5235) );
  XOR U16891 ( .A(n5945), .B(n5946), .Z(n5233) );
  ANDN U16892 ( .B(n5947), .A(n5948), .Z(n5945) );
  AND U16893 ( .A(a[46]), .B(b[73]), .Z(n5944) );
  XNOR U16894 ( .A(n5949), .B(n5238), .Z(n5240) );
  XOR U16895 ( .A(n5950), .B(n5951), .Z(n5238) );
  ANDN U16896 ( .B(n5952), .A(n5953), .Z(n5950) );
  AND U16897 ( .A(a[47]), .B(b[72]), .Z(n5949) );
  XNOR U16898 ( .A(n5954), .B(n5243), .Z(n5245) );
  XOR U16899 ( .A(n5955), .B(n5956), .Z(n5243) );
  ANDN U16900 ( .B(n5957), .A(n5958), .Z(n5955) );
  AND U16901 ( .A(a[48]), .B(b[71]), .Z(n5954) );
  XNOR U16902 ( .A(n5959), .B(n5248), .Z(n5250) );
  XOR U16903 ( .A(n5960), .B(n5961), .Z(n5248) );
  ANDN U16904 ( .B(n5962), .A(n5963), .Z(n5960) );
  AND U16905 ( .A(a[49]), .B(b[70]), .Z(n5959) );
  XNOR U16906 ( .A(n5964), .B(n5253), .Z(n5255) );
  XOR U16907 ( .A(n5965), .B(n5966), .Z(n5253) );
  ANDN U16908 ( .B(n5967), .A(n5968), .Z(n5965) );
  AND U16909 ( .A(a[50]), .B(b[69]), .Z(n5964) );
  XNOR U16910 ( .A(n5969), .B(n5258), .Z(n5260) );
  XOR U16911 ( .A(n5970), .B(n5971), .Z(n5258) );
  ANDN U16912 ( .B(n5972), .A(n5973), .Z(n5970) );
  AND U16913 ( .A(a[51]), .B(b[68]), .Z(n5969) );
  XNOR U16914 ( .A(n5974), .B(n5263), .Z(n5265) );
  XOR U16915 ( .A(n5975), .B(n5976), .Z(n5263) );
  ANDN U16916 ( .B(n5977), .A(n5978), .Z(n5975) );
  AND U16917 ( .A(a[52]), .B(b[67]), .Z(n5974) );
  XNOR U16918 ( .A(n5979), .B(n5268), .Z(n5270) );
  XOR U16919 ( .A(n5980), .B(n5981), .Z(n5268) );
  ANDN U16920 ( .B(n5982), .A(n5983), .Z(n5980) );
  AND U16921 ( .A(a[53]), .B(b[66]), .Z(n5979) );
  XNOR U16922 ( .A(n5984), .B(n5273), .Z(n5275) );
  XOR U16923 ( .A(n5985), .B(n5986), .Z(n5273) );
  ANDN U16924 ( .B(n5987), .A(n5988), .Z(n5985) );
  AND U16925 ( .A(a[54]), .B(b[65]), .Z(n5984) );
  XNOR U16926 ( .A(n5989), .B(n5278), .Z(n5280) );
  XOR U16927 ( .A(n5990), .B(n5991), .Z(n5278) );
  ANDN U16928 ( .B(n5992), .A(n5993), .Z(n5990) );
  AND U16929 ( .A(a[55]), .B(b[64]), .Z(n5989) );
  XNOR U16930 ( .A(n5994), .B(n5283), .Z(n5285) );
  XOR U16931 ( .A(n5995), .B(n5996), .Z(n5283) );
  ANDN U16932 ( .B(n5997), .A(n5998), .Z(n5995) );
  AND U16933 ( .A(a[56]), .B(b[63]), .Z(n5994) );
  XNOR U16934 ( .A(n5999), .B(n5288), .Z(n5290) );
  XOR U16935 ( .A(n6000), .B(n6001), .Z(n5288) );
  ANDN U16936 ( .B(n6002), .A(n6003), .Z(n6000) );
  AND U16937 ( .A(a[57]), .B(b[62]), .Z(n5999) );
  XNOR U16938 ( .A(n6004), .B(n5293), .Z(n5295) );
  XOR U16939 ( .A(n6005), .B(n6006), .Z(n5293) );
  ANDN U16940 ( .B(n6007), .A(n6008), .Z(n6005) );
  AND U16941 ( .A(a[58]), .B(b[61]), .Z(n6004) );
  XNOR U16942 ( .A(n6009), .B(n5298), .Z(n5300) );
  XOR U16943 ( .A(n6010), .B(n6011), .Z(n5298) );
  ANDN U16944 ( .B(n6012), .A(n6013), .Z(n6010) );
  AND U16945 ( .A(a[59]), .B(b[60]), .Z(n6009) );
  XNOR U16946 ( .A(n6014), .B(n5303), .Z(n5305) );
  XOR U16947 ( .A(n6015), .B(n6016), .Z(n5303) );
  ANDN U16948 ( .B(n6017), .A(n6018), .Z(n6015) );
  AND U16949 ( .A(a[60]), .B(b[59]), .Z(n6014) );
  XNOR U16950 ( .A(n6019), .B(n5308), .Z(n5310) );
  XOR U16951 ( .A(n6020), .B(n6021), .Z(n5308) );
  ANDN U16952 ( .B(n6022), .A(n6023), .Z(n6020) );
  AND U16953 ( .A(a[61]), .B(b[58]), .Z(n6019) );
  XNOR U16954 ( .A(n6024), .B(n5313), .Z(n5315) );
  XOR U16955 ( .A(n6025), .B(n6026), .Z(n5313) );
  ANDN U16956 ( .B(n6027), .A(n6028), .Z(n6025) );
  AND U16957 ( .A(a[62]), .B(b[57]), .Z(n6024) );
  XNOR U16958 ( .A(n6029), .B(n5318), .Z(n5320) );
  XOR U16959 ( .A(n6030), .B(n6031), .Z(n5318) );
  ANDN U16960 ( .B(n6032), .A(n6033), .Z(n6030) );
  AND U16961 ( .A(a[63]), .B(b[56]), .Z(n6029) );
  XNOR U16962 ( .A(n6034), .B(n5323), .Z(n5325) );
  XOR U16963 ( .A(n6035), .B(n6036), .Z(n5323) );
  ANDN U16964 ( .B(n6037), .A(n6038), .Z(n6035) );
  AND U16965 ( .A(a[64]), .B(b[55]), .Z(n6034) );
  XNOR U16966 ( .A(n6039), .B(n5328), .Z(n5330) );
  XOR U16967 ( .A(n6040), .B(n6041), .Z(n5328) );
  ANDN U16968 ( .B(n6042), .A(n6043), .Z(n6040) );
  AND U16969 ( .A(a[65]), .B(b[54]), .Z(n6039) );
  XNOR U16970 ( .A(n6044), .B(n5333), .Z(n5335) );
  XOR U16971 ( .A(n6045), .B(n6046), .Z(n5333) );
  ANDN U16972 ( .B(n6047), .A(n6048), .Z(n6045) );
  AND U16973 ( .A(a[66]), .B(b[53]), .Z(n6044) );
  XNOR U16974 ( .A(n6049), .B(n5338), .Z(n5340) );
  XOR U16975 ( .A(n6050), .B(n6051), .Z(n5338) );
  ANDN U16976 ( .B(n6052), .A(n6053), .Z(n6050) );
  AND U16977 ( .A(a[67]), .B(b[52]), .Z(n6049) );
  XNOR U16978 ( .A(n6054), .B(n5343), .Z(n5345) );
  XOR U16979 ( .A(n6055), .B(n6056), .Z(n5343) );
  ANDN U16980 ( .B(n6057), .A(n6058), .Z(n6055) );
  AND U16981 ( .A(a[68]), .B(b[51]), .Z(n6054) );
  XNOR U16982 ( .A(n6059), .B(n5348), .Z(n5350) );
  XOR U16983 ( .A(n6060), .B(n6061), .Z(n5348) );
  ANDN U16984 ( .B(n6062), .A(n6063), .Z(n6060) );
  AND U16985 ( .A(a[69]), .B(b[50]), .Z(n6059) );
  XNOR U16986 ( .A(n6064), .B(n5353), .Z(n5355) );
  XOR U16987 ( .A(n6065), .B(n6066), .Z(n5353) );
  ANDN U16988 ( .B(n6067), .A(n6068), .Z(n6065) );
  AND U16989 ( .A(a[70]), .B(b[49]), .Z(n6064) );
  XNOR U16990 ( .A(n6069), .B(n5358), .Z(n5360) );
  XOR U16991 ( .A(n6070), .B(n6071), .Z(n5358) );
  ANDN U16992 ( .B(n6072), .A(n6073), .Z(n6070) );
  AND U16993 ( .A(a[71]), .B(b[48]), .Z(n6069) );
  XNOR U16994 ( .A(n6074), .B(n5363), .Z(n5365) );
  XOR U16995 ( .A(n6075), .B(n6076), .Z(n5363) );
  ANDN U16996 ( .B(n6077), .A(n6078), .Z(n6075) );
  AND U16997 ( .A(a[72]), .B(b[47]), .Z(n6074) );
  XNOR U16998 ( .A(n6079), .B(n5368), .Z(n5370) );
  XOR U16999 ( .A(n6080), .B(n6081), .Z(n5368) );
  ANDN U17000 ( .B(n6082), .A(n6083), .Z(n6080) );
  AND U17001 ( .A(a[73]), .B(b[46]), .Z(n6079) );
  XNOR U17002 ( .A(n6084), .B(n5373), .Z(n5375) );
  XOR U17003 ( .A(n6085), .B(n6086), .Z(n5373) );
  ANDN U17004 ( .B(n6087), .A(n6088), .Z(n6085) );
  AND U17005 ( .A(a[74]), .B(b[45]), .Z(n6084) );
  XNOR U17006 ( .A(n6089), .B(n5378), .Z(n5380) );
  XOR U17007 ( .A(n6090), .B(n6091), .Z(n5378) );
  ANDN U17008 ( .B(n6092), .A(n6093), .Z(n6090) );
  AND U17009 ( .A(a[75]), .B(b[44]), .Z(n6089) );
  XNOR U17010 ( .A(n6094), .B(n5383), .Z(n5385) );
  XOR U17011 ( .A(n6095), .B(n6096), .Z(n5383) );
  ANDN U17012 ( .B(n6097), .A(n6098), .Z(n6095) );
  AND U17013 ( .A(a[76]), .B(b[43]), .Z(n6094) );
  XNOR U17014 ( .A(n6099), .B(n5388), .Z(n5390) );
  XOR U17015 ( .A(n6100), .B(n6101), .Z(n5388) );
  ANDN U17016 ( .B(n6102), .A(n6103), .Z(n6100) );
  AND U17017 ( .A(a[77]), .B(b[42]), .Z(n6099) );
  XNOR U17018 ( .A(n6104), .B(n5393), .Z(n5395) );
  XOR U17019 ( .A(n6105), .B(n6106), .Z(n5393) );
  ANDN U17020 ( .B(n6107), .A(n6108), .Z(n6105) );
  AND U17021 ( .A(a[78]), .B(b[41]), .Z(n6104) );
  XNOR U17022 ( .A(n6109), .B(n5398), .Z(n5400) );
  XOR U17023 ( .A(n6110), .B(n6111), .Z(n5398) );
  ANDN U17024 ( .B(n6112), .A(n6113), .Z(n6110) );
  AND U17025 ( .A(a[79]), .B(b[40]), .Z(n6109) );
  XNOR U17026 ( .A(n6114), .B(n5403), .Z(n5405) );
  XOR U17027 ( .A(n6115), .B(n6116), .Z(n5403) );
  ANDN U17028 ( .B(n6117), .A(n6118), .Z(n6115) );
  AND U17029 ( .A(a[80]), .B(b[39]), .Z(n6114) );
  XNOR U17030 ( .A(n6119), .B(n5408), .Z(n5410) );
  XOR U17031 ( .A(n6120), .B(n6121), .Z(n5408) );
  ANDN U17032 ( .B(n6122), .A(n6123), .Z(n6120) );
  AND U17033 ( .A(a[81]), .B(b[38]), .Z(n6119) );
  XNOR U17034 ( .A(n6124), .B(n5413), .Z(n5415) );
  XOR U17035 ( .A(n6125), .B(n6126), .Z(n5413) );
  ANDN U17036 ( .B(n6127), .A(n6128), .Z(n6125) );
  AND U17037 ( .A(a[82]), .B(b[37]), .Z(n6124) );
  XNOR U17038 ( .A(n6129), .B(n5418), .Z(n5420) );
  XOR U17039 ( .A(n6130), .B(n6131), .Z(n5418) );
  ANDN U17040 ( .B(n6132), .A(n6133), .Z(n6130) );
  AND U17041 ( .A(a[83]), .B(b[36]), .Z(n6129) );
  XNOR U17042 ( .A(n6134), .B(n5423), .Z(n5425) );
  XOR U17043 ( .A(n6135), .B(n6136), .Z(n5423) );
  ANDN U17044 ( .B(n6137), .A(n6138), .Z(n6135) );
  AND U17045 ( .A(a[84]), .B(b[35]), .Z(n6134) );
  XNOR U17046 ( .A(n6139), .B(n5428), .Z(n5430) );
  XOR U17047 ( .A(n6140), .B(n6141), .Z(n5428) );
  ANDN U17048 ( .B(n6142), .A(n6143), .Z(n6140) );
  AND U17049 ( .A(a[85]), .B(b[34]), .Z(n6139) );
  XNOR U17050 ( .A(n6144), .B(n5433), .Z(n5435) );
  XOR U17051 ( .A(n6145), .B(n6146), .Z(n5433) );
  ANDN U17052 ( .B(n6147), .A(n6148), .Z(n6145) );
  AND U17053 ( .A(a[86]), .B(b[33]), .Z(n6144) );
  XNOR U17054 ( .A(n6149), .B(n5438), .Z(n5440) );
  XOR U17055 ( .A(n6150), .B(n6151), .Z(n5438) );
  ANDN U17056 ( .B(n6152), .A(n6153), .Z(n6150) );
  AND U17057 ( .A(a[87]), .B(b[32]), .Z(n6149) );
  XNOR U17058 ( .A(n6154), .B(n5443), .Z(n5445) );
  XOR U17059 ( .A(n6155), .B(n6156), .Z(n5443) );
  ANDN U17060 ( .B(n6157), .A(n6158), .Z(n6155) );
  AND U17061 ( .A(a[88]), .B(b[31]), .Z(n6154) );
  XNOR U17062 ( .A(n6159), .B(n5448), .Z(n5450) );
  XOR U17063 ( .A(n6160), .B(n6161), .Z(n5448) );
  ANDN U17064 ( .B(n6162), .A(n6163), .Z(n6160) );
  AND U17065 ( .A(a[89]), .B(b[30]), .Z(n6159) );
  XNOR U17066 ( .A(n6164), .B(n5453), .Z(n5455) );
  XOR U17067 ( .A(n6165), .B(n6166), .Z(n5453) );
  ANDN U17068 ( .B(n6167), .A(n6168), .Z(n6165) );
  AND U17069 ( .A(a[90]), .B(b[29]), .Z(n6164) );
  XNOR U17070 ( .A(n6169), .B(n5458), .Z(n5460) );
  XOR U17071 ( .A(n6170), .B(n6171), .Z(n5458) );
  ANDN U17072 ( .B(n6172), .A(n6173), .Z(n6170) );
  AND U17073 ( .A(a[91]), .B(b[28]), .Z(n6169) );
  XNOR U17074 ( .A(n6174), .B(n5463), .Z(n5465) );
  XOR U17075 ( .A(n6175), .B(n6176), .Z(n5463) );
  ANDN U17076 ( .B(n6177), .A(n6178), .Z(n6175) );
  AND U17077 ( .A(a[92]), .B(b[27]), .Z(n6174) );
  XNOR U17078 ( .A(n6179), .B(n5468), .Z(n5470) );
  XOR U17079 ( .A(n6180), .B(n6181), .Z(n5468) );
  ANDN U17080 ( .B(n6182), .A(n6183), .Z(n6180) );
  AND U17081 ( .A(a[93]), .B(b[26]), .Z(n6179) );
  XNOR U17082 ( .A(n6184), .B(n5473), .Z(n5475) );
  XOR U17083 ( .A(n6185), .B(n6186), .Z(n5473) );
  ANDN U17084 ( .B(n6187), .A(n6188), .Z(n6185) );
  AND U17085 ( .A(a[94]), .B(b[25]), .Z(n6184) );
  XNOR U17086 ( .A(n6189), .B(n5478), .Z(n5480) );
  XOR U17087 ( .A(n6190), .B(n6191), .Z(n5478) );
  ANDN U17088 ( .B(n6192), .A(n6193), .Z(n6190) );
  AND U17089 ( .A(a[95]), .B(b[24]), .Z(n6189) );
  XNOR U17090 ( .A(n6194), .B(n5483), .Z(n5485) );
  XOR U17091 ( .A(n6195), .B(n6196), .Z(n5483) );
  ANDN U17092 ( .B(n6197), .A(n6198), .Z(n6195) );
  AND U17093 ( .A(a[96]), .B(b[23]), .Z(n6194) );
  XNOR U17094 ( .A(n6199), .B(n5488), .Z(n5490) );
  XOR U17095 ( .A(n6200), .B(n6201), .Z(n5488) );
  ANDN U17096 ( .B(n6202), .A(n6203), .Z(n6200) );
  AND U17097 ( .A(a[97]), .B(b[22]), .Z(n6199) );
  XNOR U17098 ( .A(n6204), .B(n5493), .Z(n5495) );
  XOR U17099 ( .A(n6205), .B(n6206), .Z(n5493) );
  ANDN U17100 ( .B(n6207), .A(n6208), .Z(n6205) );
  AND U17101 ( .A(a[98]), .B(b[21]), .Z(n6204) );
  XNOR U17102 ( .A(n6209), .B(n5498), .Z(n5500) );
  XOR U17103 ( .A(n6210), .B(n6211), .Z(n5498) );
  ANDN U17104 ( .B(n6212), .A(n6213), .Z(n6210) );
  AND U17105 ( .A(a[99]), .B(b[20]), .Z(n6209) );
  XNOR U17106 ( .A(n6214), .B(n5503), .Z(n5505) );
  XOR U17107 ( .A(n6215), .B(n6216), .Z(n5503) );
  ANDN U17108 ( .B(n6217), .A(n6218), .Z(n6215) );
  AND U17109 ( .A(b[19]), .B(a[100]), .Z(n6214) );
  XNOR U17110 ( .A(n6219), .B(n5508), .Z(n5510) );
  XOR U17111 ( .A(n6220), .B(n6221), .Z(n5508) );
  ANDN U17112 ( .B(n6222), .A(n6223), .Z(n6220) );
  AND U17113 ( .A(b[18]), .B(a[101]), .Z(n6219) );
  XNOR U17114 ( .A(n6224), .B(n5513), .Z(n5515) );
  XOR U17115 ( .A(n6225), .B(n6226), .Z(n5513) );
  ANDN U17116 ( .B(n6227), .A(n6228), .Z(n6225) );
  AND U17117 ( .A(b[17]), .B(a[102]), .Z(n6224) );
  XNOR U17118 ( .A(n6229), .B(n5518), .Z(n5520) );
  XOR U17119 ( .A(n6230), .B(n6231), .Z(n5518) );
  ANDN U17120 ( .B(n6232), .A(n6233), .Z(n6230) );
  AND U17121 ( .A(b[16]), .B(a[103]), .Z(n6229) );
  XNOR U17122 ( .A(n6234), .B(n5523), .Z(n5525) );
  XOR U17123 ( .A(n6235), .B(n6236), .Z(n5523) );
  ANDN U17124 ( .B(n6237), .A(n6238), .Z(n6235) );
  AND U17125 ( .A(b[15]), .B(a[104]), .Z(n6234) );
  XNOR U17126 ( .A(n6239), .B(n5528), .Z(n5530) );
  XOR U17127 ( .A(n6240), .B(n6241), .Z(n5528) );
  ANDN U17128 ( .B(n6242), .A(n6243), .Z(n6240) );
  AND U17129 ( .A(b[14]), .B(a[105]), .Z(n6239) );
  XNOR U17130 ( .A(n6244), .B(n5533), .Z(n5535) );
  XOR U17131 ( .A(n6245), .B(n6246), .Z(n5533) );
  ANDN U17132 ( .B(n6247), .A(n6248), .Z(n6245) );
  AND U17133 ( .A(b[13]), .B(a[106]), .Z(n6244) );
  XNOR U17134 ( .A(n6249), .B(n5538), .Z(n5540) );
  XOR U17135 ( .A(n6250), .B(n6251), .Z(n5538) );
  ANDN U17136 ( .B(n6252), .A(n6253), .Z(n6250) );
  AND U17137 ( .A(b[12]), .B(a[107]), .Z(n6249) );
  XNOR U17138 ( .A(n6254), .B(n5543), .Z(n5545) );
  XOR U17139 ( .A(n6255), .B(n6256), .Z(n5543) );
  ANDN U17140 ( .B(n6257), .A(n6258), .Z(n6255) );
  AND U17141 ( .A(b[11]), .B(a[108]), .Z(n6254) );
  XNOR U17142 ( .A(n6259), .B(n5548), .Z(n5550) );
  XOR U17143 ( .A(n6260), .B(n6261), .Z(n5548) );
  ANDN U17144 ( .B(n6262), .A(n6263), .Z(n6260) );
  AND U17145 ( .A(b[10]), .B(a[109]), .Z(n6259) );
  XNOR U17146 ( .A(n6264), .B(n5553), .Z(n5555) );
  XOR U17147 ( .A(n6265), .B(n6266), .Z(n5553) );
  ANDN U17148 ( .B(n6267), .A(n6268), .Z(n6265) );
  AND U17149 ( .A(b[9]), .B(a[110]), .Z(n6264) );
  XNOR U17150 ( .A(n6269), .B(n5558), .Z(n5560) );
  XOR U17151 ( .A(n6270), .B(n6271), .Z(n5558) );
  ANDN U17152 ( .B(n6272), .A(n6273), .Z(n6270) );
  AND U17153 ( .A(b[8]), .B(a[111]), .Z(n6269) );
  XNOR U17154 ( .A(n6274), .B(n5563), .Z(n5565) );
  XOR U17155 ( .A(n6275), .B(n6276), .Z(n5563) );
  ANDN U17156 ( .B(n6277), .A(n6278), .Z(n6275) );
  AND U17157 ( .A(b[7]), .B(a[112]), .Z(n6274) );
  XNOR U17158 ( .A(n6279), .B(n5568), .Z(n5570) );
  XOR U17159 ( .A(n6280), .B(n6281), .Z(n5568) );
  ANDN U17160 ( .B(n6282), .A(n6283), .Z(n6280) );
  AND U17161 ( .A(b[6]), .B(a[113]), .Z(n6279) );
  XNOR U17162 ( .A(n6284), .B(n5573), .Z(n5575) );
  XOR U17163 ( .A(n6285), .B(n6286), .Z(n5573) );
  ANDN U17164 ( .B(n6287), .A(n6288), .Z(n6285) );
  AND U17165 ( .A(b[5]), .B(a[114]), .Z(n6284) );
  XNOR U17166 ( .A(n6289), .B(n5578), .Z(n5580) );
  XOR U17167 ( .A(n6290), .B(n6291), .Z(n5578) );
  ANDN U17168 ( .B(n6292), .A(n6293), .Z(n6290) );
  AND U17169 ( .A(b[4]), .B(a[115]), .Z(n6289) );
  XNOR U17170 ( .A(n6294), .B(n6295), .Z(n5592) );
  NANDN U17171 ( .A(n6296), .B(n6297), .Z(n6295) );
  XNOR U17172 ( .A(n6298), .B(n5583), .Z(n5585) );
  XNOR U17173 ( .A(n6299), .B(n6300), .Z(n5583) );
  AND U17174 ( .A(n6301), .B(n6302), .Z(n6299) );
  AND U17175 ( .A(b[3]), .B(a[116]), .Z(n6298) );
  NAND U17176 ( .A(a[119]), .B(b[0]), .Z(n4886) );
  XNOR U17177 ( .A(n5600), .B(n5601), .Z(c[118]) );
  XNOR U17178 ( .A(n6296), .B(n6297), .Z(n5601) );
  XOR U17179 ( .A(n6294), .B(n6303), .Z(n6297) );
  NAND U17180 ( .A(b[1]), .B(a[117]), .Z(n6303) );
  XOR U17181 ( .A(n6302), .B(n6304), .Z(n6296) );
  XOR U17182 ( .A(n6294), .B(n6301), .Z(n6304) );
  XNOR U17183 ( .A(n6305), .B(n6300), .Z(n6301) );
  AND U17184 ( .A(b[2]), .B(a[116]), .Z(n6305) );
  NANDN U17185 ( .A(n6306), .B(n6307), .Z(n6294) );
  XOR U17186 ( .A(n6300), .B(n6292), .Z(n6308) );
  XNOR U17187 ( .A(n6291), .B(n6287), .Z(n6309) );
  XNOR U17188 ( .A(n6286), .B(n6282), .Z(n6310) );
  XNOR U17189 ( .A(n6281), .B(n6277), .Z(n6311) );
  XNOR U17190 ( .A(n6276), .B(n6272), .Z(n6312) );
  XNOR U17191 ( .A(n6271), .B(n6267), .Z(n6313) );
  XNOR U17192 ( .A(n6266), .B(n6262), .Z(n6314) );
  XNOR U17193 ( .A(n6261), .B(n6257), .Z(n6315) );
  XNOR U17194 ( .A(n6256), .B(n6252), .Z(n6316) );
  XNOR U17195 ( .A(n6251), .B(n6247), .Z(n6317) );
  XNOR U17196 ( .A(n6246), .B(n6242), .Z(n6318) );
  XNOR U17197 ( .A(n6241), .B(n6237), .Z(n6319) );
  XNOR U17198 ( .A(n6236), .B(n6232), .Z(n6320) );
  XNOR U17199 ( .A(n6231), .B(n6227), .Z(n6321) );
  XNOR U17200 ( .A(n6226), .B(n6222), .Z(n6322) );
  XNOR U17201 ( .A(n6221), .B(n6217), .Z(n6323) );
  XNOR U17202 ( .A(n6216), .B(n6212), .Z(n6324) );
  XNOR U17203 ( .A(n6211), .B(n6207), .Z(n6325) );
  XNOR U17204 ( .A(n6206), .B(n6202), .Z(n6326) );
  XNOR U17205 ( .A(n6201), .B(n6197), .Z(n6327) );
  XNOR U17206 ( .A(n6196), .B(n6192), .Z(n6328) );
  XNOR U17207 ( .A(n6191), .B(n6187), .Z(n6329) );
  XNOR U17208 ( .A(n6186), .B(n6182), .Z(n6330) );
  XNOR U17209 ( .A(n6181), .B(n6177), .Z(n6331) );
  XNOR U17210 ( .A(n6176), .B(n6172), .Z(n6332) );
  XNOR U17211 ( .A(n6171), .B(n6167), .Z(n6333) );
  XNOR U17212 ( .A(n6166), .B(n6162), .Z(n6334) );
  XNOR U17213 ( .A(n6161), .B(n6157), .Z(n6335) );
  XNOR U17214 ( .A(n6156), .B(n6152), .Z(n6336) );
  XNOR U17215 ( .A(n6151), .B(n6147), .Z(n6337) );
  XNOR U17216 ( .A(n6146), .B(n6142), .Z(n6338) );
  XNOR U17217 ( .A(n6141), .B(n6137), .Z(n6339) );
  XNOR U17218 ( .A(n6136), .B(n6132), .Z(n6340) );
  XNOR U17219 ( .A(n6131), .B(n6127), .Z(n6341) );
  XNOR U17220 ( .A(n6126), .B(n6122), .Z(n6342) );
  XNOR U17221 ( .A(n6121), .B(n6117), .Z(n6343) );
  XNOR U17222 ( .A(n6116), .B(n6112), .Z(n6344) );
  XNOR U17223 ( .A(n6111), .B(n6107), .Z(n6345) );
  XNOR U17224 ( .A(n6106), .B(n6102), .Z(n6346) );
  XNOR U17225 ( .A(n6101), .B(n6097), .Z(n6347) );
  XNOR U17226 ( .A(n6096), .B(n6092), .Z(n6348) );
  XNOR U17227 ( .A(n6091), .B(n6087), .Z(n6349) );
  XNOR U17228 ( .A(n6086), .B(n6082), .Z(n6350) );
  XNOR U17229 ( .A(n6081), .B(n6077), .Z(n6351) );
  XNOR U17230 ( .A(n6076), .B(n6072), .Z(n6352) );
  XNOR U17231 ( .A(n6071), .B(n6067), .Z(n6353) );
  XNOR U17232 ( .A(n6066), .B(n6062), .Z(n6354) );
  XNOR U17233 ( .A(n6061), .B(n6057), .Z(n6355) );
  XNOR U17234 ( .A(n6056), .B(n6052), .Z(n6356) );
  XNOR U17235 ( .A(n6051), .B(n6047), .Z(n6357) );
  XNOR U17236 ( .A(n6046), .B(n6042), .Z(n6358) );
  XNOR U17237 ( .A(n6041), .B(n6037), .Z(n6359) );
  XNOR U17238 ( .A(n6036), .B(n6032), .Z(n6360) );
  XNOR U17239 ( .A(n6031), .B(n6027), .Z(n6361) );
  XNOR U17240 ( .A(n6026), .B(n6022), .Z(n6362) );
  XNOR U17241 ( .A(n6021), .B(n6017), .Z(n6363) );
  XNOR U17242 ( .A(n6016), .B(n6012), .Z(n6364) );
  XNOR U17243 ( .A(n6011), .B(n6007), .Z(n6365) );
  XNOR U17244 ( .A(n6006), .B(n6002), .Z(n6366) );
  XNOR U17245 ( .A(n6001), .B(n5997), .Z(n6367) );
  XNOR U17246 ( .A(n5996), .B(n5992), .Z(n6368) );
  XNOR U17247 ( .A(n5991), .B(n5987), .Z(n6369) );
  XNOR U17248 ( .A(n5986), .B(n5982), .Z(n6370) );
  XNOR U17249 ( .A(n5981), .B(n5977), .Z(n6371) );
  XNOR U17250 ( .A(n5976), .B(n5972), .Z(n6372) );
  XNOR U17251 ( .A(n5971), .B(n5967), .Z(n6373) );
  XNOR U17252 ( .A(n5966), .B(n5962), .Z(n6374) );
  XNOR U17253 ( .A(n5961), .B(n5957), .Z(n6375) );
  XNOR U17254 ( .A(n5956), .B(n5952), .Z(n6376) );
  XNOR U17255 ( .A(n5951), .B(n5947), .Z(n6377) );
  XNOR U17256 ( .A(n5946), .B(n5942), .Z(n6378) );
  XNOR U17257 ( .A(n5941), .B(n5937), .Z(n6379) );
  XNOR U17258 ( .A(n5936), .B(n5932), .Z(n6380) );
  XNOR U17259 ( .A(n5931), .B(n5927), .Z(n6381) );
  XNOR U17260 ( .A(n5926), .B(n5922), .Z(n6382) );
  XNOR U17261 ( .A(n5921), .B(n5917), .Z(n6383) );
  XNOR U17262 ( .A(n5916), .B(n5912), .Z(n6384) );
  XNOR U17263 ( .A(n5911), .B(n5907), .Z(n6385) );
  XNOR U17264 ( .A(n5906), .B(n5902), .Z(n6386) );
  XNOR U17265 ( .A(n5901), .B(n5897), .Z(n6387) );
  XNOR U17266 ( .A(n5896), .B(n5892), .Z(n6388) );
  XNOR U17267 ( .A(n5891), .B(n5887), .Z(n6389) );
  XNOR U17268 ( .A(n5886), .B(n5882), .Z(n6390) );
  XNOR U17269 ( .A(n5881), .B(n5877), .Z(n6391) );
  XNOR U17270 ( .A(n5876), .B(n5872), .Z(n6392) );
  XNOR U17271 ( .A(n5871), .B(n5867), .Z(n6393) );
  XNOR U17272 ( .A(n5866), .B(n5862), .Z(n6394) );
  XNOR U17273 ( .A(n5861), .B(n5857), .Z(n6395) );
  XNOR U17274 ( .A(n5856), .B(n5852), .Z(n6396) );
  XNOR U17275 ( .A(n5851), .B(n5847), .Z(n6397) );
  XNOR U17276 ( .A(n5846), .B(n5842), .Z(n6398) );
  XNOR U17277 ( .A(n5841), .B(n5837), .Z(n6399) );
  XNOR U17278 ( .A(n5836), .B(n5832), .Z(n6400) );
  XNOR U17279 ( .A(n5831), .B(n5827), .Z(n6401) );
  XNOR U17280 ( .A(n5826), .B(n5822), .Z(n6402) );
  XNOR U17281 ( .A(n5821), .B(n5817), .Z(n6403) );
  XNOR U17282 ( .A(n5816), .B(n5812), .Z(n6404) );
  XNOR U17283 ( .A(n5811), .B(n5807), .Z(n6405) );
  XNOR U17284 ( .A(n5806), .B(n5802), .Z(n6406) );
  XNOR U17285 ( .A(n5801), .B(n5797), .Z(n6407) );
  XNOR U17286 ( .A(n5796), .B(n5792), .Z(n6408) );
  XNOR U17287 ( .A(n5791), .B(n5787), .Z(n6409) );
  XNOR U17288 ( .A(n5786), .B(n5782), .Z(n6410) );
  XNOR U17289 ( .A(n5781), .B(n5777), .Z(n6411) );
  XNOR U17290 ( .A(n5776), .B(n5772), .Z(n6412) );
  XNOR U17291 ( .A(n5771), .B(n5767), .Z(n6413) );
  XNOR U17292 ( .A(n5766), .B(n5762), .Z(n6414) );
  XNOR U17293 ( .A(n5761), .B(n5757), .Z(n6415) );
  XNOR U17294 ( .A(n5756), .B(n5752), .Z(n6416) );
  XNOR U17295 ( .A(n5751), .B(n5747), .Z(n6417) );
  XNOR U17296 ( .A(n5746), .B(n5742), .Z(n6418) );
  XNOR U17297 ( .A(n5741), .B(n5737), .Z(n6419) );
  XNOR U17298 ( .A(n5736), .B(n5732), .Z(n6420) );
  XNOR U17299 ( .A(n5731), .B(n5727), .Z(n6421) );
  XNOR U17300 ( .A(n5726), .B(n5722), .Z(n6422) );
  XOR U17301 ( .A(n6423), .B(n5721), .Z(n5722) );
  AND U17302 ( .A(a[0]), .B(b[118]), .Z(n6423) );
  XNOR U17303 ( .A(n6424), .B(n5721), .Z(n5723) );
  XNOR U17304 ( .A(n6425), .B(n6426), .Z(n5721) );
  ANDN U17305 ( .B(n6427), .A(n6428), .Z(n6425) );
  AND U17306 ( .A(a[1]), .B(b[117]), .Z(n6424) );
  XNOR U17307 ( .A(n6429), .B(n5726), .Z(n5728) );
  XOR U17308 ( .A(n6430), .B(n6431), .Z(n5726) );
  ANDN U17309 ( .B(n6432), .A(n6433), .Z(n6430) );
  AND U17310 ( .A(a[2]), .B(b[116]), .Z(n6429) );
  XNOR U17311 ( .A(n6434), .B(n5731), .Z(n5733) );
  XOR U17312 ( .A(n6435), .B(n6436), .Z(n5731) );
  ANDN U17313 ( .B(n6437), .A(n6438), .Z(n6435) );
  AND U17314 ( .A(a[3]), .B(b[115]), .Z(n6434) );
  XNOR U17315 ( .A(n6439), .B(n5736), .Z(n5738) );
  XOR U17316 ( .A(n6440), .B(n6441), .Z(n5736) );
  ANDN U17317 ( .B(n6442), .A(n6443), .Z(n6440) );
  AND U17318 ( .A(a[4]), .B(b[114]), .Z(n6439) );
  XNOR U17319 ( .A(n6444), .B(n5741), .Z(n5743) );
  XOR U17320 ( .A(n6445), .B(n6446), .Z(n5741) );
  ANDN U17321 ( .B(n6447), .A(n6448), .Z(n6445) );
  AND U17322 ( .A(a[5]), .B(b[113]), .Z(n6444) );
  XNOR U17323 ( .A(n6449), .B(n5746), .Z(n5748) );
  XOR U17324 ( .A(n6450), .B(n6451), .Z(n5746) );
  ANDN U17325 ( .B(n6452), .A(n6453), .Z(n6450) );
  AND U17326 ( .A(a[6]), .B(b[112]), .Z(n6449) );
  XNOR U17327 ( .A(n6454), .B(n5751), .Z(n5753) );
  XOR U17328 ( .A(n6455), .B(n6456), .Z(n5751) );
  ANDN U17329 ( .B(n6457), .A(n6458), .Z(n6455) );
  AND U17330 ( .A(a[7]), .B(b[111]), .Z(n6454) );
  XNOR U17331 ( .A(n6459), .B(n5756), .Z(n5758) );
  XOR U17332 ( .A(n6460), .B(n6461), .Z(n5756) );
  ANDN U17333 ( .B(n6462), .A(n6463), .Z(n6460) );
  AND U17334 ( .A(a[8]), .B(b[110]), .Z(n6459) );
  XNOR U17335 ( .A(n6464), .B(n5761), .Z(n5763) );
  XOR U17336 ( .A(n6465), .B(n6466), .Z(n5761) );
  ANDN U17337 ( .B(n6467), .A(n6468), .Z(n6465) );
  AND U17338 ( .A(a[9]), .B(b[109]), .Z(n6464) );
  XNOR U17339 ( .A(n6469), .B(n5766), .Z(n5768) );
  XOR U17340 ( .A(n6470), .B(n6471), .Z(n5766) );
  ANDN U17341 ( .B(n6472), .A(n6473), .Z(n6470) );
  AND U17342 ( .A(a[10]), .B(b[108]), .Z(n6469) );
  XNOR U17343 ( .A(n6474), .B(n5771), .Z(n5773) );
  XOR U17344 ( .A(n6475), .B(n6476), .Z(n5771) );
  ANDN U17345 ( .B(n6477), .A(n6478), .Z(n6475) );
  AND U17346 ( .A(a[11]), .B(b[107]), .Z(n6474) );
  XNOR U17347 ( .A(n6479), .B(n5776), .Z(n5778) );
  XOR U17348 ( .A(n6480), .B(n6481), .Z(n5776) );
  ANDN U17349 ( .B(n6482), .A(n6483), .Z(n6480) );
  AND U17350 ( .A(a[12]), .B(b[106]), .Z(n6479) );
  XNOR U17351 ( .A(n6484), .B(n5781), .Z(n5783) );
  XOR U17352 ( .A(n6485), .B(n6486), .Z(n5781) );
  ANDN U17353 ( .B(n6487), .A(n6488), .Z(n6485) );
  AND U17354 ( .A(a[13]), .B(b[105]), .Z(n6484) );
  XNOR U17355 ( .A(n6489), .B(n5786), .Z(n5788) );
  XOR U17356 ( .A(n6490), .B(n6491), .Z(n5786) );
  ANDN U17357 ( .B(n6492), .A(n6493), .Z(n6490) );
  AND U17358 ( .A(a[14]), .B(b[104]), .Z(n6489) );
  XNOR U17359 ( .A(n6494), .B(n5791), .Z(n5793) );
  XOR U17360 ( .A(n6495), .B(n6496), .Z(n5791) );
  ANDN U17361 ( .B(n6497), .A(n6498), .Z(n6495) );
  AND U17362 ( .A(a[15]), .B(b[103]), .Z(n6494) );
  XNOR U17363 ( .A(n6499), .B(n5796), .Z(n5798) );
  XOR U17364 ( .A(n6500), .B(n6501), .Z(n5796) );
  ANDN U17365 ( .B(n6502), .A(n6503), .Z(n6500) );
  AND U17366 ( .A(a[16]), .B(b[102]), .Z(n6499) );
  XNOR U17367 ( .A(n6504), .B(n5801), .Z(n5803) );
  XOR U17368 ( .A(n6505), .B(n6506), .Z(n5801) );
  ANDN U17369 ( .B(n6507), .A(n6508), .Z(n6505) );
  AND U17370 ( .A(a[17]), .B(b[101]), .Z(n6504) );
  XNOR U17371 ( .A(n6509), .B(n5806), .Z(n5808) );
  XOR U17372 ( .A(n6510), .B(n6511), .Z(n5806) );
  ANDN U17373 ( .B(n6512), .A(n6513), .Z(n6510) );
  AND U17374 ( .A(a[18]), .B(b[100]), .Z(n6509) );
  XNOR U17375 ( .A(n6514), .B(n5811), .Z(n5813) );
  XOR U17376 ( .A(n6515), .B(n6516), .Z(n5811) );
  ANDN U17377 ( .B(n6517), .A(n6518), .Z(n6515) );
  AND U17378 ( .A(a[19]), .B(b[99]), .Z(n6514) );
  XNOR U17379 ( .A(n6519), .B(n5816), .Z(n5818) );
  XOR U17380 ( .A(n6520), .B(n6521), .Z(n5816) );
  ANDN U17381 ( .B(n6522), .A(n6523), .Z(n6520) );
  AND U17382 ( .A(a[20]), .B(b[98]), .Z(n6519) );
  XNOR U17383 ( .A(n6524), .B(n5821), .Z(n5823) );
  XOR U17384 ( .A(n6525), .B(n6526), .Z(n5821) );
  ANDN U17385 ( .B(n6527), .A(n6528), .Z(n6525) );
  AND U17386 ( .A(a[21]), .B(b[97]), .Z(n6524) );
  XNOR U17387 ( .A(n6529), .B(n5826), .Z(n5828) );
  XOR U17388 ( .A(n6530), .B(n6531), .Z(n5826) );
  ANDN U17389 ( .B(n6532), .A(n6533), .Z(n6530) );
  AND U17390 ( .A(a[22]), .B(b[96]), .Z(n6529) );
  XNOR U17391 ( .A(n6534), .B(n5831), .Z(n5833) );
  XOR U17392 ( .A(n6535), .B(n6536), .Z(n5831) );
  ANDN U17393 ( .B(n6537), .A(n6538), .Z(n6535) );
  AND U17394 ( .A(a[23]), .B(b[95]), .Z(n6534) );
  XNOR U17395 ( .A(n6539), .B(n5836), .Z(n5838) );
  XOR U17396 ( .A(n6540), .B(n6541), .Z(n5836) );
  ANDN U17397 ( .B(n6542), .A(n6543), .Z(n6540) );
  AND U17398 ( .A(a[24]), .B(b[94]), .Z(n6539) );
  XNOR U17399 ( .A(n6544), .B(n5841), .Z(n5843) );
  XOR U17400 ( .A(n6545), .B(n6546), .Z(n5841) );
  ANDN U17401 ( .B(n6547), .A(n6548), .Z(n6545) );
  AND U17402 ( .A(a[25]), .B(b[93]), .Z(n6544) );
  XNOR U17403 ( .A(n6549), .B(n5846), .Z(n5848) );
  XOR U17404 ( .A(n6550), .B(n6551), .Z(n5846) );
  ANDN U17405 ( .B(n6552), .A(n6553), .Z(n6550) );
  AND U17406 ( .A(a[26]), .B(b[92]), .Z(n6549) );
  XNOR U17407 ( .A(n6554), .B(n5851), .Z(n5853) );
  XOR U17408 ( .A(n6555), .B(n6556), .Z(n5851) );
  ANDN U17409 ( .B(n6557), .A(n6558), .Z(n6555) );
  AND U17410 ( .A(a[27]), .B(b[91]), .Z(n6554) );
  XNOR U17411 ( .A(n6559), .B(n5856), .Z(n5858) );
  XOR U17412 ( .A(n6560), .B(n6561), .Z(n5856) );
  ANDN U17413 ( .B(n6562), .A(n6563), .Z(n6560) );
  AND U17414 ( .A(a[28]), .B(b[90]), .Z(n6559) );
  XNOR U17415 ( .A(n6564), .B(n5861), .Z(n5863) );
  XOR U17416 ( .A(n6565), .B(n6566), .Z(n5861) );
  ANDN U17417 ( .B(n6567), .A(n6568), .Z(n6565) );
  AND U17418 ( .A(a[29]), .B(b[89]), .Z(n6564) );
  XNOR U17419 ( .A(n6569), .B(n5866), .Z(n5868) );
  XOR U17420 ( .A(n6570), .B(n6571), .Z(n5866) );
  ANDN U17421 ( .B(n6572), .A(n6573), .Z(n6570) );
  AND U17422 ( .A(a[30]), .B(b[88]), .Z(n6569) );
  XNOR U17423 ( .A(n6574), .B(n5871), .Z(n5873) );
  XOR U17424 ( .A(n6575), .B(n6576), .Z(n5871) );
  ANDN U17425 ( .B(n6577), .A(n6578), .Z(n6575) );
  AND U17426 ( .A(a[31]), .B(b[87]), .Z(n6574) );
  XNOR U17427 ( .A(n6579), .B(n5876), .Z(n5878) );
  XOR U17428 ( .A(n6580), .B(n6581), .Z(n5876) );
  ANDN U17429 ( .B(n6582), .A(n6583), .Z(n6580) );
  AND U17430 ( .A(a[32]), .B(b[86]), .Z(n6579) );
  XNOR U17431 ( .A(n6584), .B(n5881), .Z(n5883) );
  XOR U17432 ( .A(n6585), .B(n6586), .Z(n5881) );
  ANDN U17433 ( .B(n6587), .A(n6588), .Z(n6585) );
  AND U17434 ( .A(a[33]), .B(b[85]), .Z(n6584) );
  XNOR U17435 ( .A(n6589), .B(n5886), .Z(n5888) );
  XOR U17436 ( .A(n6590), .B(n6591), .Z(n5886) );
  ANDN U17437 ( .B(n6592), .A(n6593), .Z(n6590) );
  AND U17438 ( .A(a[34]), .B(b[84]), .Z(n6589) );
  XNOR U17439 ( .A(n6594), .B(n5891), .Z(n5893) );
  XOR U17440 ( .A(n6595), .B(n6596), .Z(n5891) );
  ANDN U17441 ( .B(n6597), .A(n6598), .Z(n6595) );
  AND U17442 ( .A(a[35]), .B(b[83]), .Z(n6594) );
  XNOR U17443 ( .A(n6599), .B(n5896), .Z(n5898) );
  XOR U17444 ( .A(n6600), .B(n6601), .Z(n5896) );
  ANDN U17445 ( .B(n6602), .A(n6603), .Z(n6600) );
  AND U17446 ( .A(a[36]), .B(b[82]), .Z(n6599) );
  XNOR U17447 ( .A(n6604), .B(n5901), .Z(n5903) );
  XOR U17448 ( .A(n6605), .B(n6606), .Z(n5901) );
  ANDN U17449 ( .B(n6607), .A(n6608), .Z(n6605) );
  AND U17450 ( .A(a[37]), .B(b[81]), .Z(n6604) );
  XNOR U17451 ( .A(n6609), .B(n5906), .Z(n5908) );
  XOR U17452 ( .A(n6610), .B(n6611), .Z(n5906) );
  ANDN U17453 ( .B(n6612), .A(n6613), .Z(n6610) );
  AND U17454 ( .A(a[38]), .B(b[80]), .Z(n6609) );
  XNOR U17455 ( .A(n6614), .B(n5911), .Z(n5913) );
  XOR U17456 ( .A(n6615), .B(n6616), .Z(n5911) );
  ANDN U17457 ( .B(n6617), .A(n6618), .Z(n6615) );
  AND U17458 ( .A(a[39]), .B(b[79]), .Z(n6614) );
  XNOR U17459 ( .A(n6619), .B(n5916), .Z(n5918) );
  XOR U17460 ( .A(n6620), .B(n6621), .Z(n5916) );
  ANDN U17461 ( .B(n6622), .A(n6623), .Z(n6620) );
  AND U17462 ( .A(a[40]), .B(b[78]), .Z(n6619) );
  XNOR U17463 ( .A(n6624), .B(n5921), .Z(n5923) );
  XOR U17464 ( .A(n6625), .B(n6626), .Z(n5921) );
  ANDN U17465 ( .B(n6627), .A(n6628), .Z(n6625) );
  AND U17466 ( .A(a[41]), .B(b[77]), .Z(n6624) );
  XNOR U17467 ( .A(n6629), .B(n5926), .Z(n5928) );
  XOR U17468 ( .A(n6630), .B(n6631), .Z(n5926) );
  ANDN U17469 ( .B(n6632), .A(n6633), .Z(n6630) );
  AND U17470 ( .A(a[42]), .B(b[76]), .Z(n6629) );
  XNOR U17471 ( .A(n6634), .B(n5931), .Z(n5933) );
  XOR U17472 ( .A(n6635), .B(n6636), .Z(n5931) );
  ANDN U17473 ( .B(n6637), .A(n6638), .Z(n6635) );
  AND U17474 ( .A(a[43]), .B(b[75]), .Z(n6634) );
  XNOR U17475 ( .A(n6639), .B(n5936), .Z(n5938) );
  XOR U17476 ( .A(n6640), .B(n6641), .Z(n5936) );
  ANDN U17477 ( .B(n6642), .A(n6643), .Z(n6640) );
  AND U17478 ( .A(a[44]), .B(b[74]), .Z(n6639) );
  XNOR U17479 ( .A(n6644), .B(n5941), .Z(n5943) );
  XOR U17480 ( .A(n6645), .B(n6646), .Z(n5941) );
  ANDN U17481 ( .B(n6647), .A(n6648), .Z(n6645) );
  AND U17482 ( .A(a[45]), .B(b[73]), .Z(n6644) );
  XNOR U17483 ( .A(n6649), .B(n5946), .Z(n5948) );
  XOR U17484 ( .A(n6650), .B(n6651), .Z(n5946) );
  ANDN U17485 ( .B(n6652), .A(n6653), .Z(n6650) );
  AND U17486 ( .A(a[46]), .B(b[72]), .Z(n6649) );
  XNOR U17487 ( .A(n6654), .B(n5951), .Z(n5953) );
  XOR U17488 ( .A(n6655), .B(n6656), .Z(n5951) );
  ANDN U17489 ( .B(n6657), .A(n6658), .Z(n6655) );
  AND U17490 ( .A(a[47]), .B(b[71]), .Z(n6654) );
  XNOR U17491 ( .A(n6659), .B(n5956), .Z(n5958) );
  XOR U17492 ( .A(n6660), .B(n6661), .Z(n5956) );
  ANDN U17493 ( .B(n6662), .A(n6663), .Z(n6660) );
  AND U17494 ( .A(a[48]), .B(b[70]), .Z(n6659) );
  XNOR U17495 ( .A(n6664), .B(n5961), .Z(n5963) );
  XOR U17496 ( .A(n6665), .B(n6666), .Z(n5961) );
  ANDN U17497 ( .B(n6667), .A(n6668), .Z(n6665) );
  AND U17498 ( .A(a[49]), .B(b[69]), .Z(n6664) );
  XNOR U17499 ( .A(n6669), .B(n5966), .Z(n5968) );
  XOR U17500 ( .A(n6670), .B(n6671), .Z(n5966) );
  ANDN U17501 ( .B(n6672), .A(n6673), .Z(n6670) );
  AND U17502 ( .A(a[50]), .B(b[68]), .Z(n6669) );
  XNOR U17503 ( .A(n6674), .B(n5971), .Z(n5973) );
  XOR U17504 ( .A(n6675), .B(n6676), .Z(n5971) );
  ANDN U17505 ( .B(n6677), .A(n6678), .Z(n6675) );
  AND U17506 ( .A(a[51]), .B(b[67]), .Z(n6674) );
  XNOR U17507 ( .A(n6679), .B(n5976), .Z(n5978) );
  XOR U17508 ( .A(n6680), .B(n6681), .Z(n5976) );
  ANDN U17509 ( .B(n6682), .A(n6683), .Z(n6680) );
  AND U17510 ( .A(a[52]), .B(b[66]), .Z(n6679) );
  XNOR U17511 ( .A(n6684), .B(n5981), .Z(n5983) );
  XOR U17512 ( .A(n6685), .B(n6686), .Z(n5981) );
  ANDN U17513 ( .B(n6687), .A(n6688), .Z(n6685) );
  AND U17514 ( .A(a[53]), .B(b[65]), .Z(n6684) );
  XNOR U17515 ( .A(n6689), .B(n5986), .Z(n5988) );
  XOR U17516 ( .A(n6690), .B(n6691), .Z(n5986) );
  ANDN U17517 ( .B(n6692), .A(n6693), .Z(n6690) );
  AND U17518 ( .A(a[54]), .B(b[64]), .Z(n6689) );
  XNOR U17519 ( .A(n6694), .B(n5991), .Z(n5993) );
  XOR U17520 ( .A(n6695), .B(n6696), .Z(n5991) );
  ANDN U17521 ( .B(n6697), .A(n6698), .Z(n6695) );
  AND U17522 ( .A(a[55]), .B(b[63]), .Z(n6694) );
  XNOR U17523 ( .A(n6699), .B(n5996), .Z(n5998) );
  XOR U17524 ( .A(n6700), .B(n6701), .Z(n5996) );
  ANDN U17525 ( .B(n6702), .A(n6703), .Z(n6700) );
  AND U17526 ( .A(a[56]), .B(b[62]), .Z(n6699) );
  XNOR U17527 ( .A(n6704), .B(n6001), .Z(n6003) );
  XOR U17528 ( .A(n6705), .B(n6706), .Z(n6001) );
  ANDN U17529 ( .B(n6707), .A(n6708), .Z(n6705) );
  AND U17530 ( .A(a[57]), .B(b[61]), .Z(n6704) );
  XNOR U17531 ( .A(n6709), .B(n6006), .Z(n6008) );
  XOR U17532 ( .A(n6710), .B(n6711), .Z(n6006) );
  ANDN U17533 ( .B(n6712), .A(n6713), .Z(n6710) );
  AND U17534 ( .A(a[58]), .B(b[60]), .Z(n6709) );
  XNOR U17535 ( .A(n6714), .B(n6011), .Z(n6013) );
  XOR U17536 ( .A(n6715), .B(n6716), .Z(n6011) );
  ANDN U17537 ( .B(n6717), .A(n6718), .Z(n6715) );
  AND U17538 ( .A(a[59]), .B(b[59]), .Z(n6714) );
  XNOR U17539 ( .A(n6719), .B(n6016), .Z(n6018) );
  XOR U17540 ( .A(n6720), .B(n6721), .Z(n6016) );
  ANDN U17541 ( .B(n6722), .A(n6723), .Z(n6720) );
  AND U17542 ( .A(a[60]), .B(b[58]), .Z(n6719) );
  XNOR U17543 ( .A(n6724), .B(n6021), .Z(n6023) );
  XOR U17544 ( .A(n6725), .B(n6726), .Z(n6021) );
  ANDN U17545 ( .B(n6727), .A(n6728), .Z(n6725) );
  AND U17546 ( .A(a[61]), .B(b[57]), .Z(n6724) );
  XNOR U17547 ( .A(n6729), .B(n6026), .Z(n6028) );
  XOR U17548 ( .A(n6730), .B(n6731), .Z(n6026) );
  ANDN U17549 ( .B(n6732), .A(n6733), .Z(n6730) );
  AND U17550 ( .A(a[62]), .B(b[56]), .Z(n6729) );
  XNOR U17551 ( .A(n6734), .B(n6031), .Z(n6033) );
  XOR U17552 ( .A(n6735), .B(n6736), .Z(n6031) );
  ANDN U17553 ( .B(n6737), .A(n6738), .Z(n6735) );
  AND U17554 ( .A(a[63]), .B(b[55]), .Z(n6734) );
  XNOR U17555 ( .A(n6739), .B(n6036), .Z(n6038) );
  XOR U17556 ( .A(n6740), .B(n6741), .Z(n6036) );
  ANDN U17557 ( .B(n6742), .A(n6743), .Z(n6740) );
  AND U17558 ( .A(a[64]), .B(b[54]), .Z(n6739) );
  XNOR U17559 ( .A(n6744), .B(n6041), .Z(n6043) );
  XOR U17560 ( .A(n6745), .B(n6746), .Z(n6041) );
  ANDN U17561 ( .B(n6747), .A(n6748), .Z(n6745) );
  AND U17562 ( .A(a[65]), .B(b[53]), .Z(n6744) );
  XNOR U17563 ( .A(n6749), .B(n6046), .Z(n6048) );
  XOR U17564 ( .A(n6750), .B(n6751), .Z(n6046) );
  ANDN U17565 ( .B(n6752), .A(n6753), .Z(n6750) );
  AND U17566 ( .A(a[66]), .B(b[52]), .Z(n6749) );
  XNOR U17567 ( .A(n6754), .B(n6051), .Z(n6053) );
  XOR U17568 ( .A(n6755), .B(n6756), .Z(n6051) );
  ANDN U17569 ( .B(n6757), .A(n6758), .Z(n6755) );
  AND U17570 ( .A(a[67]), .B(b[51]), .Z(n6754) );
  XNOR U17571 ( .A(n6759), .B(n6056), .Z(n6058) );
  XOR U17572 ( .A(n6760), .B(n6761), .Z(n6056) );
  ANDN U17573 ( .B(n6762), .A(n6763), .Z(n6760) );
  AND U17574 ( .A(a[68]), .B(b[50]), .Z(n6759) );
  XNOR U17575 ( .A(n6764), .B(n6061), .Z(n6063) );
  XOR U17576 ( .A(n6765), .B(n6766), .Z(n6061) );
  ANDN U17577 ( .B(n6767), .A(n6768), .Z(n6765) );
  AND U17578 ( .A(a[69]), .B(b[49]), .Z(n6764) );
  XNOR U17579 ( .A(n6769), .B(n6066), .Z(n6068) );
  XOR U17580 ( .A(n6770), .B(n6771), .Z(n6066) );
  ANDN U17581 ( .B(n6772), .A(n6773), .Z(n6770) );
  AND U17582 ( .A(a[70]), .B(b[48]), .Z(n6769) );
  XNOR U17583 ( .A(n6774), .B(n6071), .Z(n6073) );
  XOR U17584 ( .A(n6775), .B(n6776), .Z(n6071) );
  ANDN U17585 ( .B(n6777), .A(n6778), .Z(n6775) );
  AND U17586 ( .A(a[71]), .B(b[47]), .Z(n6774) );
  XNOR U17587 ( .A(n6779), .B(n6076), .Z(n6078) );
  XOR U17588 ( .A(n6780), .B(n6781), .Z(n6076) );
  ANDN U17589 ( .B(n6782), .A(n6783), .Z(n6780) );
  AND U17590 ( .A(a[72]), .B(b[46]), .Z(n6779) );
  XNOR U17591 ( .A(n6784), .B(n6081), .Z(n6083) );
  XOR U17592 ( .A(n6785), .B(n6786), .Z(n6081) );
  ANDN U17593 ( .B(n6787), .A(n6788), .Z(n6785) );
  AND U17594 ( .A(a[73]), .B(b[45]), .Z(n6784) );
  XNOR U17595 ( .A(n6789), .B(n6086), .Z(n6088) );
  XOR U17596 ( .A(n6790), .B(n6791), .Z(n6086) );
  ANDN U17597 ( .B(n6792), .A(n6793), .Z(n6790) );
  AND U17598 ( .A(a[74]), .B(b[44]), .Z(n6789) );
  XNOR U17599 ( .A(n6794), .B(n6091), .Z(n6093) );
  XOR U17600 ( .A(n6795), .B(n6796), .Z(n6091) );
  ANDN U17601 ( .B(n6797), .A(n6798), .Z(n6795) );
  AND U17602 ( .A(a[75]), .B(b[43]), .Z(n6794) );
  XNOR U17603 ( .A(n6799), .B(n6096), .Z(n6098) );
  XOR U17604 ( .A(n6800), .B(n6801), .Z(n6096) );
  ANDN U17605 ( .B(n6802), .A(n6803), .Z(n6800) );
  AND U17606 ( .A(a[76]), .B(b[42]), .Z(n6799) );
  XNOR U17607 ( .A(n6804), .B(n6101), .Z(n6103) );
  XOR U17608 ( .A(n6805), .B(n6806), .Z(n6101) );
  ANDN U17609 ( .B(n6807), .A(n6808), .Z(n6805) );
  AND U17610 ( .A(a[77]), .B(b[41]), .Z(n6804) );
  XNOR U17611 ( .A(n6809), .B(n6106), .Z(n6108) );
  XOR U17612 ( .A(n6810), .B(n6811), .Z(n6106) );
  ANDN U17613 ( .B(n6812), .A(n6813), .Z(n6810) );
  AND U17614 ( .A(a[78]), .B(b[40]), .Z(n6809) );
  XNOR U17615 ( .A(n6814), .B(n6111), .Z(n6113) );
  XOR U17616 ( .A(n6815), .B(n6816), .Z(n6111) );
  ANDN U17617 ( .B(n6817), .A(n6818), .Z(n6815) );
  AND U17618 ( .A(a[79]), .B(b[39]), .Z(n6814) );
  XNOR U17619 ( .A(n6819), .B(n6116), .Z(n6118) );
  XOR U17620 ( .A(n6820), .B(n6821), .Z(n6116) );
  ANDN U17621 ( .B(n6822), .A(n6823), .Z(n6820) );
  AND U17622 ( .A(a[80]), .B(b[38]), .Z(n6819) );
  XNOR U17623 ( .A(n6824), .B(n6121), .Z(n6123) );
  XOR U17624 ( .A(n6825), .B(n6826), .Z(n6121) );
  ANDN U17625 ( .B(n6827), .A(n6828), .Z(n6825) );
  AND U17626 ( .A(a[81]), .B(b[37]), .Z(n6824) );
  XNOR U17627 ( .A(n6829), .B(n6126), .Z(n6128) );
  XOR U17628 ( .A(n6830), .B(n6831), .Z(n6126) );
  ANDN U17629 ( .B(n6832), .A(n6833), .Z(n6830) );
  AND U17630 ( .A(a[82]), .B(b[36]), .Z(n6829) );
  XNOR U17631 ( .A(n6834), .B(n6131), .Z(n6133) );
  XOR U17632 ( .A(n6835), .B(n6836), .Z(n6131) );
  ANDN U17633 ( .B(n6837), .A(n6838), .Z(n6835) );
  AND U17634 ( .A(a[83]), .B(b[35]), .Z(n6834) );
  XNOR U17635 ( .A(n6839), .B(n6136), .Z(n6138) );
  XOR U17636 ( .A(n6840), .B(n6841), .Z(n6136) );
  ANDN U17637 ( .B(n6842), .A(n6843), .Z(n6840) );
  AND U17638 ( .A(a[84]), .B(b[34]), .Z(n6839) );
  XNOR U17639 ( .A(n6844), .B(n6141), .Z(n6143) );
  XOR U17640 ( .A(n6845), .B(n6846), .Z(n6141) );
  ANDN U17641 ( .B(n6847), .A(n6848), .Z(n6845) );
  AND U17642 ( .A(a[85]), .B(b[33]), .Z(n6844) );
  XNOR U17643 ( .A(n6849), .B(n6146), .Z(n6148) );
  XOR U17644 ( .A(n6850), .B(n6851), .Z(n6146) );
  ANDN U17645 ( .B(n6852), .A(n6853), .Z(n6850) );
  AND U17646 ( .A(a[86]), .B(b[32]), .Z(n6849) );
  XNOR U17647 ( .A(n6854), .B(n6151), .Z(n6153) );
  XOR U17648 ( .A(n6855), .B(n6856), .Z(n6151) );
  ANDN U17649 ( .B(n6857), .A(n6858), .Z(n6855) );
  AND U17650 ( .A(a[87]), .B(b[31]), .Z(n6854) );
  XNOR U17651 ( .A(n6859), .B(n6156), .Z(n6158) );
  XOR U17652 ( .A(n6860), .B(n6861), .Z(n6156) );
  ANDN U17653 ( .B(n6862), .A(n6863), .Z(n6860) );
  AND U17654 ( .A(a[88]), .B(b[30]), .Z(n6859) );
  XNOR U17655 ( .A(n6864), .B(n6161), .Z(n6163) );
  XOR U17656 ( .A(n6865), .B(n6866), .Z(n6161) );
  ANDN U17657 ( .B(n6867), .A(n6868), .Z(n6865) );
  AND U17658 ( .A(a[89]), .B(b[29]), .Z(n6864) );
  XNOR U17659 ( .A(n6869), .B(n6166), .Z(n6168) );
  XOR U17660 ( .A(n6870), .B(n6871), .Z(n6166) );
  ANDN U17661 ( .B(n6872), .A(n6873), .Z(n6870) );
  AND U17662 ( .A(a[90]), .B(b[28]), .Z(n6869) );
  XNOR U17663 ( .A(n6874), .B(n6171), .Z(n6173) );
  XOR U17664 ( .A(n6875), .B(n6876), .Z(n6171) );
  ANDN U17665 ( .B(n6877), .A(n6878), .Z(n6875) );
  AND U17666 ( .A(a[91]), .B(b[27]), .Z(n6874) );
  XNOR U17667 ( .A(n6879), .B(n6176), .Z(n6178) );
  XOR U17668 ( .A(n6880), .B(n6881), .Z(n6176) );
  ANDN U17669 ( .B(n6882), .A(n6883), .Z(n6880) );
  AND U17670 ( .A(a[92]), .B(b[26]), .Z(n6879) );
  XNOR U17671 ( .A(n6884), .B(n6181), .Z(n6183) );
  XOR U17672 ( .A(n6885), .B(n6886), .Z(n6181) );
  ANDN U17673 ( .B(n6887), .A(n6888), .Z(n6885) );
  AND U17674 ( .A(a[93]), .B(b[25]), .Z(n6884) );
  XNOR U17675 ( .A(n6889), .B(n6186), .Z(n6188) );
  XOR U17676 ( .A(n6890), .B(n6891), .Z(n6186) );
  ANDN U17677 ( .B(n6892), .A(n6893), .Z(n6890) );
  AND U17678 ( .A(a[94]), .B(b[24]), .Z(n6889) );
  XNOR U17679 ( .A(n6894), .B(n6191), .Z(n6193) );
  XOR U17680 ( .A(n6895), .B(n6896), .Z(n6191) );
  ANDN U17681 ( .B(n6897), .A(n6898), .Z(n6895) );
  AND U17682 ( .A(a[95]), .B(b[23]), .Z(n6894) );
  XNOR U17683 ( .A(n6899), .B(n6196), .Z(n6198) );
  XOR U17684 ( .A(n6900), .B(n6901), .Z(n6196) );
  ANDN U17685 ( .B(n6902), .A(n6903), .Z(n6900) );
  AND U17686 ( .A(a[96]), .B(b[22]), .Z(n6899) );
  XNOR U17687 ( .A(n6904), .B(n6201), .Z(n6203) );
  XOR U17688 ( .A(n6905), .B(n6906), .Z(n6201) );
  ANDN U17689 ( .B(n6907), .A(n6908), .Z(n6905) );
  AND U17690 ( .A(a[97]), .B(b[21]), .Z(n6904) );
  XNOR U17691 ( .A(n6909), .B(n6206), .Z(n6208) );
  XOR U17692 ( .A(n6910), .B(n6911), .Z(n6206) );
  ANDN U17693 ( .B(n6912), .A(n6913), .Z(n6910) );
  AND U17694 ( .A(a[98]), .B(b[20]), .Z(n6909) );
  XNOR U17695 ( .A(n6914), .B(n6211), .Z(n6213) );
  XOR U17696 ( .A(n6915), .B(n6916), .Z(n6211) );
  ANDN U17697 ( .B(n6917), .A(n6918), .Z(n6915) );
  AND U17698 ( .A(a[99]), .B(b[19]), .Z(n6914) );
  XNOR U17699 ( .A(n6919), .B(n6216), .Z(n6218) );
  XOR U17700 ( .A(n6920), .B(n6921), .Z(n6216) );
  ANDN U17701 ( .B(n6922), .A(n6923), .Z(n6920) );
  AND U17702 ( .A(b[18]), .B(a[100]), .Z(n6919) );
  XNOR U17703 ( .A(n6924), .B(n6221), .Z(n6223) );
  XOR U17704 ( .A(n6925), .B(n6926), .Z(n6221) );
  ANDN U17705 ( .B(n6927), .A(n6928), .Z(n6925) );
  AND U17706 ( .A(b[17]), .B(a[101]), .Z(n6924) );
  XNOR U17707 ( .A(n6929), .B(n6226), .Z(n6228) );
  XOR U17708 ( .A(n6930), .B(n6931), .Z(n6226) );
  ANDN U17709 ( .B(n6932), .A(n6933), .Z(n6930) );
  AND U17710 ( .A(b[16]), .B(a[102]), .Z(n6929) );
  XNOR U17711 ( .A(n6934), .B(n6231), .Z(n6233) );
  XOR U17712 ( .A(n6935), .B(n6936), .Z(n6231) );
  ANDN U17713 ( .B(n6937), .A(n6938), .Z(n6935) );
  AND U17714 ( .A(b[15]), .B(a[103]), .Z(n6934) );
  XNOR U17715 ( .A(n6939), .B(n6236), .Z(n6238) );
  XOR U17716 ( .A(n6940), .B(n6941), .Z(n6236) );
  ANDN U17717 ( .B(n6942), .A(n6943), .Z(n6940) );
  AND U17718 ( .A(b[14]), .B(a[104]), .Z(n6939) );
  XNOR U17719 ( .A(n6944), .B(n6241), .Z(n6243) );
  XOR U17720 ( .A(n6945), .B(n6946), .Z(n6241) );
  ANDN U17721 ( .B(n6947), .A(n6948), .Z(n6945) );
  AND U17722 ( .A(b[13]), .B(a[105]), .Z(n6944) );
  XNOR U17723 ( .A(n6949), .B(n6246), .Z(n6248) );
  XOR U17724 ( .A(n6950), .B(n6951), .Z(n6246) );
  ANDN U17725 ( .B(n6952), .A(n6953), .Z(n6950) );
  AND U17726 ( .A(b[12]), .B(a[106]), .Z(n6949) );
  XNOR U17727 ( .A(n6954), .B(n6251), .Z(n6253) );
  XOR U17728 ( .A(n6955), .B(n6956), .Z(n6251) );
  ANDN U17729 ( .B(n6957), .A(n6958), .Z(n6955) );
  AND U17730 ( .A(b[11]), .B(a[107]), .Z(n6954) );
  XNOR U17731 ( .A(n6959), .B(n6256), .Z(n6258) );
  XOR U17732 ( .A(n6960), .B(n6961), .Z(n6256) );
  ANDN U17733 ( .B(n6962), .A(n6963), .Z(n6960) );
  AND U17734 ( .A(b[10]), .B(a[108]), .Z(n6959) );
  XNOR U17735 ( .A(n6964), .B(n6261), .Z(n6263) );
  XOR U17736 ( .A(n6965), .B(n6966), .Z(n6261) );
  ANDN U17737 ( .B(n6967), .A(n6968), .Z(n6965) );
  AND U17738 ( .A(b[9]), .B(a[109]), .Z(n6964) );
  XNOR U17739 ( .A(n6969), .B(n6266), .Z(n6268) );
  XOR U17740 ( .A(n6970), .B(n6971), .Z(n6266) );
  ANDN U17741 ( .B(n6972), .A(n6973), .Z(n6970) );
  AND U17742 ( .A(b[8]), .B(a[110]), .Z(n6969) );
  XNOR U17743 ( .A(n6974), .B(n6271), .Z(n6273) );
  XOR U17744 ( .A(n6975), .B(n6976), .Z(n6271) );
  ANDN U17745 ( .B(n6977), .A(n6978), .Z(n6975) );
  AND U17746 ( .A(b[7]), .B(a[111]), .Z(n6974) );
  XNOR U17747 ( .A(n6979), .B(n6276), .Z(n6278) );
  XOR U17748 ( .A(n6980), .B(n6981), .Z(n6276) );
  ANDN U17749 ( .B(n6982), .A(n6983), .Z(n6980) );
  AND U17750 ( .A(b[6]), .B(a[112]), .Z(n6979) );
  XNOR U17751 ( .A(n6984), .B(n6281), .Z(n6283) );
  XOR U17752 ( .A(n6985), .B(n6986), .Z(n6281) );
  ANDN U17753 ( .B(n6987), .A(n6988), .Z(n6985) );
  AND U17754 ( .A(b[5]), .B(a[113]), .Z(n6984) );
  XNOR U17755 ( .A(n6989), .B(n6286), .Z(n6288) );
  XOR U17756 ( .A(n6990), .B(n6991), .Z(n6286) );
  ANDN U17757 ( .B(n6992), .A(n6993), .Z(n6990) );
  AND U17758 ( .A(b[4]), .B(a[114]), .Z(n6989) );
  XNOR U17759 ( .A(n6994), .B(n6995), .Z(n6300) );
  NANDN U17760 ( .A(n6996), .B(n6997), .Z(n6995) );
  XNOR U17761 ( .A(n6998), .B(n6291), .Z(n6293) );
  XNOR U17762 ( .A(n6999), .B(n7000), .Z(n6291) );
  AND U17763 ( .A(n7001), .B(n7002), .Z(n6999) );
  AND U17764 ( .A(b[3]), .B(a[115]), .Z(n6998) );
  NAND U17765 ( .A(a[118]), .B(b[0]), .Z(n5600) );
  XNOR U17766 ( .A(n6306), .B(n6307), .Z(c[117]) );
  XNOR U17767 ( .A(n6996), .B(n6997), .Z(n6307) );
  XOR U17768 ( .A(n6994), .B(n7003), .Z(n6997) );
  NAND U17769 ( .A(b[1]), .B(a[116]), .Z(n7003) );
  XOR U17770 ( .A(n7002), .B(n7004), .Z(n6996) );
  XOR U17771 ( .A(n6994), .B(n7001), .Z(n7004) );
  XNOR U17772 ( .A(n7005), .B(n7000), .Z(n7001) );
  AND U17773 ( .A(b[2]), .B(a[115]), .Z(n7005) );
  NANDN U17774 ( .A(n7006), .B(n7007), .Z(n6994) );
  XOR U17775 ( .A(n7000), .B(n6992), .Z(n7008) );
  XNOR U17776 ( .A(n6991), .B(n6987), .Z(n7009) );
  XNOR U17777 ( .A(n6986), .B(n6982), .Z(n7010) );
  XNOR U17778 ( .A(n6981), .B(n6977), .Z(n7011) );
  XNOR U17779 ( .A(n6976), .B(n6972), .Z(n7012) );
  XNOR U17780 ( .A(n6971), .B(n6967), .Z(n7013) );
  XNOR U17781 ( .A(n6966), .B(n6962), .Z(n7014) );
  XNOR U17782 ( .A(n6961), .B(n6957), .Z(n7015) );
  XNOR U17783 ( .A(n6956), .B(n6952), .Z(n7016) );
  XNOR U17784 ( .A(n6951), .B(n6947), .Z(n7017) );
  XNOR U17785 ( .A(n6946), .B(n6942), .Z(n7018) );
  XNOR U17786 ( .A(n6941), .B(n6937), .Z(n7019) );
  XNOR U17787 ( .A(n6936), .B(n6932), .Z(n7020) );
  XNOR U17788 ( .A(n6931), .B(n6927), .Z(n7021) );
  XNOR U17789 ( .A(n6926), .B(n6922), .Z(n7022) );
  XNOR U17790 ( .A(n6921), .B(n6917), .Z(n7023) );
  XNOR U17791 ( .A(n6916), .B(n6912), .Z(n7024) );
  XNOR U17792 ( .A(n6911), .B(n6907), .Z(n7025) );
  XNOR U17793 ( .A(n6906), .B(n6902), .Z(n7026) );
  XNOR U17794 ( .A(n6901), .B(n6897), .Z(n7027) );
  XNOR U17795 ( .A(n6896), .B(n6892), .Z(n7028) );
  XNOR U17796 ( .A(n6891), .B(n6887), .Z(n7029) );
  XNOR U17797 ( .A(n6886), .B(n6882), .Z(n7030) );
  XNOR U17798 ( .A(n6881), .B(n6877), .Z(n7031) );
  XNOR U17799 ( .A(n6876), .B(n6872), .Z(n7032) );
  XNOR U17800 ( .A(n6871), .B(n6867), .Z(n7033) );
  XNOR U17801 ( .A(n6866), .B(n6862), .Z(n7034) );
  XNOR U17802 ( .A(n6861), .B(n6857), .Z(n7035) );
  XNOR U17803 ( .A(n6856), .B(n6852), .Z(n7036) );
  XNOR U17804 ( .A(n6851), .B(n6847), .Z(n7037) );
  XNOR U17805 ( .A(n6846), .B(n6842), .Z(n7038) );
  XNOR U17806 ( .A(n6841), .B(n6837), .Z(n7039) );
  XNOR U17807 ( .A(n6836), .B(n6832), .Z(n7040) );
  XNOR U17808 ( .A(n6831), .B(n6827), .Z(n7041) );
  XNOR U17809 ( .A(n6826), .B(n6822), .Z(n7042) );
  XNOR U17810 ( .A(n6821), .B(n6817), .Z(n7043) );
  XNOR U17811 ( .A(n6816), .B(n6812), .Z(n7044) );
  XNOR U17812 ( .A(n6811), .B(n6807), .Z(n7045) );
  XNOR U17813 ( .A(n6806), .B(n6802), .Z(n7046) );
  XNOR U17814 ( .A(n6801), .B(n6797), .Z(n7047) );
  XNOR U17815 ( .A(n6796), .B(n6792), .Z(n7048) );
  XNOR U17816 ( .A(n6791), .B(n6787), .Z(n7049) );
  XNOR U17817 ( .A(n6786), .B(n6782), .Z(n7050) );
  XNOR U17818 ( .A(n6781), .B(n6777), .Z(n7051) );
  XNOR U17819 ( .A(n6776), .B(n6772), .Z(n7052) );
  XNOR U17820 ( .A(n6771), .B(n6767), .Z(n7053) );
  XNOR U17821 ( .A(n6766), .B(n6762), .Z(n7054) );
  XNOR U17822 ( .A(n6761), .B(n6757), .Z(n7055) );
  XNOR U17823 ( .A(n6756), .B(n6752), .Z(n7056) );
  XNOR U17824 ( .A(n6751), .B(n6747), .Z(n7057) );
  XNOR U17825 ( .A(n6746), .B(n6742), .Z(n7058) );
  XNOR U17826 ( .A(n6741), .B(n6737), .Z(n7059) );
  XNOR U17827 ( .A(n6736), .B(n6732), .Z(n7060) );
  XNOR U17828 ( .A(n6731), .B(n6727), .Z(n7061) );
  XNOR U17829 ( .A(n6726), .B(n6722), .Z(n7062) );
  XNOR U17830 ( .A(n6721), .B(n6717), .Z(n7063) );
  XNOR U17831 ( .A(n6716), .B(n6712), .Z(n7064) );
  XNOR U17832 ( .A(n6711), .B(n6707), .Z(n7065) );
  XNOR U17833 ( .A(n6706), .B(n6702), .Z(n7066) );
  XNOR U17834 ( .A(n6701), .B(n6697), .Z(n7067) );
  XNOR U17835 ( .A(n6696), .B(n6692), .Z(n7068) );
  XNOR U17836 ( .A(n6691), .B(n6687), .Z(n7069) );
  XNOR U17837 ( .A(n6686), .B(n6682), .Z(n7070) );
  XNOR U17838 ( .A(n6681), .B(n6677), .Z(n7071) );
  XNOR U17839 ( .A(n6676), .B(n6672), .Z(n7072) );
  XNOR U17840 ( .A(n6671), .B(n6667), .Z(n7073) );
  XNOR U17841 ( .A(n6666), .B(n6662), .Z(n7074) );
  XNOR U17842 ( .A(n6661), .B(n6657), .Z(n7075) );
  XNOR U17843 ( .A(n6656), .B(n6652), .Z(n7076) );
  XNOR U17844 ( .A(n6651), .B(n6647), .Z(n7077) );
  XNOR U17845 ( .A(n6646), .B(n6642), .Z(n7078) );
  XNOR U17846 ( .A(n6641), .B(n6637), .Z(n7079) );
  XNOR U17847 ( .A(n6636), .B(n6632), .Z(n7080) );
  XNOR U17848 ( .A(n6631), .B(n6627), .Z(n7081) );
  XNOR U17849 ( .A(n6626), .B(n6622), .Z(n7082) );
  XNOR U17850 ( .A(n6621), .B(n6617), .Z(n7083) );
  XNOR U17851 ( .A(n6616), .B(n6612), .Z(n7084) );
  XNOR U17852 ( .A(n6611), .B(n6607), .Z(n7085) );
  XNOR U17853 ( .A(n6606), .B(n6602), .Z(n7086) );
  XNOR U17854 ( .A(n6601), .B(n6597), .Z(n7087) );
  XNOR U17855 ( .A(n6596), .B(n6592), .Z(n7088) );
  XNOR U17856 ( .A(n6591), .B(n6587), .Z(n7089) );
  XNOR U17857 ( .A(n6586), .B(n6582), .Z(n7090) );
  XNOR U17858 ( .A(n6581), .B(n6577), .Z(n7091) );
  XNOR U17859 ( .A(n6576), .B(n6572), .Z(n7092) );
  XNOR U17860 ( .A(n6571), .B(n6567), .Z(n7093) );
  XNOR U17861 ( .A(n6566), .B(n6562), .Z(n7094) );
  XNOR U17862 ( .A(n6561), .B(n6557), .Z(n7095) );
  XNOR U17863 ( .A(n6556), .B(n6552), .Z(n7096) );
  XNOR U17864 ( .A(n6551), .B(n6547), .Z(n7097) );
  XNOR U17865 ( .A(n6546), .B(n6542), .Z(n7098) );
  XNOR U17866 ( .A(n6541), .B(n6537), .Z(n7099) );
  XNOR U17867 ( .A(n6536), .B(n6532), .Z(n7100) );
  XNOR U17868 ( .A(n6531), .B(n6527), .Z(n7101) );
  XNOR U17869 ( .A(n6526), .B(n6522), .Z(n7102) );
  XNOR U17870 ( .A(n6521), .B(n6517), .Z(n7103) );
  XNOR U17871 ( .A(n6516), .B(n6512), .Z(n7104) );
  XNOR U17872 ( .A(n6511), .B(n6507), .Z(n7105) );
  XNOR U17873 ( .A(n6506), .B(n6502), .Z(n7106) );
  XNOR U17874 ( .A(n6501), .B(n6497), .Z(n7107) );
  XNOR U17875 ( .A(n6496), .B(n6492), .Z(n7108) );
  XNOR U17876 ( .A(n6491), .B(n6487), .Z(n7109) );
  XNOR U17877 ( .A(n6486), .B(n6482), .Z(n7110) );
  XNOR U17878 ( .A(n6481), .B(n6477), .Z(n7111) );
  XNOR U17879 ( .A(n6476), .B(n6472), .Z(n7112) );
  XNOR U17880 ( .A(n6471), .B(n6467), .Z(n7113) );
  XNOR U17881 ( .A(n6466), .B(n6462), .Z(n7114) );
  XNOR U17882 ( .A(n6461), .B(n6457), .Z(n7115) );
  XNOR U17883 ( .A(n6456), .B(n6452), .Z(n7116) );
  XNOR U17884 ( .A(n6451), .B(n6447), .Z(n7117) );
  XNOR U17885 ( .A(n6446), .B(n6442), .Z(n7118) );
  XNOR U17886 ( .A(n6441), .B(n6437), .Z(n7119) );
  XNOR U17887 ( .A(n6436), .B(n6432), .Z(n7120) );
  XNOR U17888 ( .A(n6431), .B(n6427), .Z(n7121) );
  XNOR U17889 ( .A(n7122), .B(n6426), .Z(n6427) );
  AND U17890 ( .A(a[0]), .B(b[117]), .Z(n7122) );
  XOR U17891 ( .A(n7123), .B(n6426), .Z(n6428) );
  XNOR U17892 ( .A(n7124), .B(n7125), .Z(n6426) );
  ANDN U17893 ( .B(n7126), .A(n7127), .Z(n7124) );
  AND U17894 ( .A(a[1]), .B(b[116]), .Z(n7123) );
  XNOR U17895 ( .A(n7128), .B(n6431), .Z(n6433) );
  XOR U17896 ( .A(n7129), .B(n7130), .Z(n6431) );
  ANDN U17897 ( .B(n7131), .A(n7132), .Z(n7129) );
  AND U17898 ( .A(a[2]), .B(b[115]), .Z(n7128) );
  XNOR U17899 ( .A(n7133), .B(n6436), .Z(n6438) );
  XOR U17900 ( .A(n7134), .B(n7135), .Z(n6436) );
  ANDN U17901 ( .B(n7136), .A(n7137), .Z(n7134) );
  AND U17902 ( .A(a[3]), .B(b[114]), .Z(n7133) );
  XNOR U17903 ( .A(n7138), .B(n6441), .Z(n6443) );
  XOR U17904 ( .A(n7139), .B(n7140), .Z(n6441) );
  ANDN U17905 ( .B(n7141), .A(n7142), .Z(n7139) );
  AND U17906 ( .A(a[4]), .B(b[113]), .Z(n7138) );
  XNOR U17907 ( .A(n7143), .B(n6446), .Z(n6448) );
  XOR U17908 ( .A(n7144), .B(n7145), .Z(n6446) );
  ANDN U17909 ( .B(n7146), .A(n7147), .Z(n7144) );
  AND U17910 ( .A(a[5]), .B(b[112]), .Z(n7143) );
  XNOR U17911 ( .A(n7148), .B(n6451), .Z(n6453) );
  XOR U17912 ( .A(n7149), .B(n7150), .Z(n6451) );
  ANDN U17913 ( .B(n7151), .A(n7152), .Z(n7149) );
  AND U17914 ( .A(a[6]), .B(b[111]), .Z(n7148) );
  XNOR U17915 ( .A(n7153), .B(n6456), .Z(n6458) );
  XOR U17916 ( .A(n7154), .B(n7155), .Z(n6456) );
  ANDN U17917 ( .B(n7156), .A(n7157), .Z(n7154) );
  AND U17918 ( .A(a[7]), .B(b[110]), .Z(n7153) );
  XNOR U17919 ( .A(n7158), .B(n6461), .Z(n6463) );
  XOR U17920 ( .A(n7159), .B(n7160), .Z(n6461) );
  ANDN U17921 ( .B(n7161), .A(n7162), .Z(n7159) );
  AND U17922 ( .A(a[8]), .B(b[109]), .Z(n7158) );
  XNOR U17923 ( .A(n7163), .B(n6466), .Z(n6468) );
  XOR U17924 ( .A(n7164), .B(n7165), .Z(n6466) );
  ANDN U17925 ( .B(n7166), .A(n7167), .Z(n7164) );
  AND U17926 ( .A(a[9]), .B(b[108]), .Z(n7163) );
  XNOR U17927 ( .A(n7168), .B(n6471), .Z(n6473) );
  XOR U17928 ( .A(n7169), .B(n7170), .Z(n6471) );
  ANDN U17929 ( .B(n7171), .A(n7172), .Z(n7169) );
  AND U17930 ( .A(a[10]), .B(b[107]), .Z(n7168) );
  XNOR U17931 ( .A(n7173), .B(n6476), .Z(n6478) );
  XOR U17932 ( .A(n7174), .B(n7175), .Z(n6476) );
  ANDN U17933 ( .B(n7176), .A(n7177), .Z(n7174) );
  AND U17934 ( .A(a[11]), .B(b[106]), .Z(n7173) );
  XNOR U17935 ( .A(n7178), .B(n6481), .Z(n6483) );
  XOR U17936 ( .A(n7179), .B(n7180), .Z(n6481) );
  ANDN U17937 ( .B(n7181), .A(n7182), .Z(n7179) );
  AND U17938 ( .A(a[12]), .B(b[105]), .Z(n7178) );
  XNOR U17939 ( .A(n7183), .B(n6486), .Z(n6488) );
  XOR U17940 ( .A(n7184), .B(n7185), .Z(n6486) );
  ANDN U17941 ( .B(n7186), .A(n7187), .Z(n7184) );
  AND U17942 ( .A(a[13]), .B(b[104]), .Z(n7183) );
  XNOR U17943 ( .A(n7188), .B(n6491), .Z(n6493) );
  XOR U17944 ( .A(n7189), .B(n7190), .Z(n6491) );
  ANDN U17945 ( .B(n7191), .A(n7192), .Z(n7189) );
  AND U17946 ( .A(a[14]), .B(b[103]), .Z(n7188) );
  XNOR U17947 ( .A(n7193), .B(n6496), .Z(n6498) );
  XOR U17948 ( .A(n7194), .B(n7195), .Z(n6496) );
  ANDN U17949 ( .B(n7196), .A(n7197), .Z(n7194) );
  AND U17950 ( .A(a[15]), .B(b[102]), .Z(n7193) );
  XNOR U17951 ( .A(n7198), .B(n6501), .Z(n6503) );
  XOR U17952 ( .A(n7199), .B(n7200), .Z(n6501) );
  ANDN U17953 ( .B(n7201), .A(n7202), .Z(n7199) );
  AND U17954 ( .A(a[16]), .B(b[101]), .Z(n7198) );
  XNOR U17955 ( .A(n7203), .B(n6506), .Z(n6508) );
  XOR U17956 ( .A(n7204), .B(n7205), .Z(n6506) );
  ANDN U17957 ( .B(n7206), .A(n7207), .Z(n7204) );
  AND U17958 ( .A(a[17]), .B(b[100]), .Z(n7203) );
  XNOR U17959 ( .A(n7208), .B(n6511), .Z(n6513) );
  XOR U17960 ( .A(n7209), .B(n7210), .Z(n6511) );
  ANDN U17961 ( .B(n7211), .A(n7212), .Z(n7209) );
  AND U17962 ( .A(a[18]), .B(b[99]), .Z(n7208) );
  XNOR U17963 ( .A(n7213), .B(n6516), .Z(n6518) );
  XOR U17964 ( .A(n7214), .B(n7215), .Z(n6516) );
  ANDN U17965 ( .B(n7216), .A(n7217), .Z(n7214) );
  AND U17966 ( .A(a[19]), .B(b[98]), .Z(n7213) );
  XNOR U17967 ( .A(n7218), .B(n6521), .Z(n6523) );
  XOR U17968 ( .A(n7219), .B(n7220), .Z(n6521) );
  ANDN U17969 ( .B(n7221), .A(n7222), .Z(n7219) );
  AND U17970 ( .A(a[20]), .B(b[97]), .Z(n7218) );
  XNOR U17971 ( .A(n7223), .B(n6526), .Z(n6528) );
  XOR U17972 ( .A(n7224), .B(n7225), .Z(n6526) );
  ANDN U17973 ( .B(n7226), .A(n7227), .Z(n7224) );
  AND U17974 ( .A(a[21]), .B(b[96]), .Z(n7223) );
  XNOR U17975 ( .A(n7228), .B(n6531), .Z(n6533) );
  XOR U17976 ( .A(n7229), .B(n7230), .Z(n6531) );
  ANDN U17977 ( .B(n7231), .A(n7232), .Z(n7229) );
  AND U17978 ( .A(a[22]), .B(b[95]), .Z(n7228) );
  XNOR U17979 ( .A(n7233), .B(n6536), .Z(n6538) );
  XOR U17980 ( .A(n7234), .B(n7235), .Z(n6536) );
  ANDN U17981 ( .B(n7236), .A(n7237), .Z(n7234) );
  AND U17982 ( .A(a[23]), .B(b[94]), .Z(n7233) );
  XNOR U17983 ( .A(n7238), .B(n6541), .Z(n6543) );
  XOR U17984 ( .A(n7239), .B(n7240), .Z(n6541) );
  ANDN U17985 ( .B(n7241), .A(n7242), .Z(n7239) );
  AND U17986 ( .A(a[24]), .B(b[93]), .Z(n7238) );
  XNOR U17987 ( .A(n7243), .B(n6546), .Z(n6548) );
  XOR U17988 ( .A(n7244), .B(n7245), .Z(n6546) );
  ANDN U17989 ( .B(n7246), .A(n7247), .Z(n7244) );
  AND U17990 ( .A(a[25]), .B(b[92]), .Z(n7243) );
  XNOR U17991 ( .A(n7248), .B(n6551), .Z(n6553) );
  XOR U17992 ( .A(n7249), .B(n7250), .Z(n6551) );
  ANDN U17993 ( .B(n7251), .A(n7252), .Z(n7249) );
  AND U17994 ( .A(a[26]), .B(b[91]), .Z(n7248) );
  XNOR U17995 ( .A(n7253), .B(n6556), .Z(n6558) );
  XOR U17996 ( .A(n7254), .B(n7255), .Z(n6556) );
  ANDN U17997 ( .B(n7256), .A(n7257), .Z(n7254) );
  AND U17998 ( .A(a[27]), .B(b[90]), .Z(n7253) );
  XNOR U17999 ( .A(n7258), .B(n6561), .Z(n6563) );
  XOR U18000 ( .A(n7259), .B(n7260), .Z(n6561) );
  ANDN U18001 ( .B(n7261), .A(n7262), .Z(n7259) );
  AND U18002 ( .A(a[28]), .B(b[89]), .Z(n7258) );
  XNOR U18003 ( .A(n7263), .B(n6566), .Z(n6568) );
  XOR U18004 ( .A(n7264), .B(n7265), .Z(n6566) );
  ANDN U18005 ( .B(n7266), .A(n7267), .Z(n7264) );
  AND U18006 ( .A(a[29]), .B(b[88]), .Z(n7263) );
  XNOR U18007 ( .A(n7268), .B(n6571), .Z(n6573) );
  XOR U18008 ( .A(n7269), .B(n7270), .Z(n6571) );
  ANDN U18009 ( .B(n7271), .A(n7272), .Z(n7269) );
  AND U18010 ( .A(a[30]), .B(b[87]), .Z(n7268) );
  XNOR U18011 ( .A(n7273), .B(n6576), .Z(n6578) );
  XOR U18012 ( .A(n7274), .B(n7275), .Z(n6576) );
  ANDN U18013 ( .B(n7276), .A(n7277), .Z(n7274) );
  AND U18014 ( .A(a[31]), .B(b[86]), .Z(n7273) );
  XNOR U18015 ( .A(n7278), .B(n6581), .Z(n6583) );
  XOR U18016 ( .A(n7279), .B(n7280), .Z(n6581) );
  ANDN U18017 ( .B(n7281), .A(n7282), .Z(n7279) );
  AND U18018 ( .A(a[32]), .B(b[85]), .Z(n7278) );
  XNOR U18019 ( .A(n7283), .B(n6586), .Z(n6588) );
  XOR U18020 ( .A(n7284), .B(n7285), .Z(n6586) );
  ANDN U18021 ( .B(n7286), .A(n7287), .Z(n7284) );
  AND U18022 ( .A(a[33]), .B(b[84]), .Z(n7283) );
  XNOR U18023 ( .A(n7288), .B(n6591), .Z(n6593) );
  XOR U18024 ( .A(n7289), .B(n7290), .Z(n6591) );
  ANDN U18025 ( .B(n7291), .A(n7292), .Z(n7289) );
  AND U18026 ( .A(a[34]), .B(b[83]), .Z(n7288) );
  XNOR U18027 ( .A(n7293), .B(n6596), .Z(n6598) );
  XOR U18028 ( .A(n7294), .B(n7295), .Z(n6596) );
  ANDN U18029 ( .B(n7296), .A(n7297), .Z(n7294) );
  AND U18030 ( .A(a[35]), .B(b[82]), .Z(n7293) );
  XNOR U18031 ( .A(n7298), .B(n6601), .Z(n6603) );
  XOR U18032 ( .A(n7299), .B(n7300), .Z(n6601) );
  ANDN U18033 ( .B(n7301), .A(n7302), .Z(n7299) );
  AND U18034 ( .A(a[36]), .B(b[81]), .Z(n7298) );
  XNOR U18035 ( .A(n7303), .B(n6606), .Z(n6608) );
  XOR U18036 ( .A(n7304), .B(n7305), .Z(n6606) );
  ANDN U18037 ( .B(n7306), .A(n7307), .Z(n7304) );
  AND U18038 ( .A(a[37]), .B(b[80]), .Z(n7303) );
  XNOR U18039 ( .A(n7308), .B(n6611), .Z(n6613) );
  XOR U18040 ( .A(n7309), .B(n7310), .Z(n6611) );
  ANDN U18041 ( .B(n7311), .A(n7312), .Z(n7309) );
  AND U18042 ( .A(a[38]), .B(b[79]), .Z(n7308) );
  XNOR U18043 ( .A(n7313), .B(n6616), .Z(n6618) );
  XOR U18044 ( .A(n7314), .B(n7315), .Z(n6616) );
  ANDN U18045 ( .B(n7316), .A(n7317), .Z(n7314) );
  AND U18046 ( .A(a[39]), .B(b[78]), .Z(n7313) );
  XNOR U18047 ( .A(n7318), .B(n6621), .Z(n6623) );
  XOR U18048 ( .A(n7319), .B(n7320), .Z(n6621) );
  ANDN U18049 ( .B(n7321), .A(n7322), .Z(n7319) );
  AND U18050 ( .A(a[40]), .B(b[77]), .Z(n7318) );
  XNOR U18051 ( .A(n7323), .B(n6626), .Z(n6628) );
  XOR U18052 ( .A(n7324), .B(n7325), .Z(n6626) );
  ANDN U18053 ( .B(n7326), .A(n7327), .Z(n7324) );
  AND U18054 ( .A(a[41]), .B(b[76]), .Z(n7323) );
  XNOR U18055 ( .A(n7328), .B(n6631), .Z(n6633) );
  XOR U18056 ( .A(n7329), .B(n7330), .Z(n6631) );
  ANDN U18057 ( .B(n7331), .A(n7332), .Z(n7329) );
  AND U18058 ( .A(a[42]), .B(b[75]), .Z(n7328) );
  XNOR U18059 ( .A(n7333), .B(n6636), .Z(n6638) );
  XOR U18060 ( .A(n7334), .B(n7335), .Z(n6636) );
  ANDN U18061 ( .B(n7336), .A(n7337), .Z(n7334) );
  AND U18062 ( .A(a[43]), .B(b[74]), .Z(n7333) );
  XNOR U18063 ( .A(n7338), .B(n6641), .Z(n6643) );
  XOR U18064 ( .A(n7339), .B(n7340), .Z(n6641) );
  ANDN U18065 ( .B(n7341), .A(n7342), .Z(n7339) );
  AND U18066 ( .A(a[44]), .B(b[73]), .Z(n7338) );
  XNOR U18067 ( .A(n7343), .B(n6646), .Z(n6648) );
  XOR U18068 ( .A(n7344), .B(n7345), .Z(n6646) );
  ANDN U18069 ( .B(n7346), .A(n7347), .Z(n7344) );
  AND U18070 ( .A(a[45]), .B(b[72]), .Z(n7343) );
  XNOR U18071 ( .A(n7348), .B(n6651), .Z(n6653) );
  XOR U18072 ( .A(n7349), .B(n7350), .Z(n6651) );
  ANDN U18073 ( .B(n7351), .A(n7352), .Z(n7349) );
  AND U18074 ( .A(a[46]), .B(b[71]), .Z(n7348) );
  XNOR U18075 ( .A(n7353), .B(n6656), .Z(n6658) );
  XOR U18076 ( .A(n7354), .B(n7355), .Z(n6656) );
  ANDN U18077 ( .B(n7356), .A(n7357), .Z(n7354) );
  AND U18078 ( .A(a[47]), .B(b[70]), .Z(n7353) );
  XNOR U18079 ( .A(n7358), .B(n6661), .Z(n6663) );
  XOR U18080 ( .A(n7359), .B(n7360), .Z(n6661) );
  ANDN U18081 ( .B(n7361), .A(n7362), .Z(n7359) );
  AND U18082 ( .A(a[48]), .B(b[69]), .Z(n7358) );
  XNOR U18083 ( .A(n7363), .B(n6666), .Z(n6668) );
  XOR U18084 ( .A(n7364), .B(n7365), .Z(n6666) );
  ANDN U18085 ( .B(n7366), .A(n7367), .Z(n7364) );
  AND U18086 ( .A(a[49]), .B(b[68]), .Z(n7363) );
  XNOR U18087 ( .A(n7368), .B(n6671), .Z(n6673) );
  XOR U18088 ( .A(n7369), .B(n7370), .Z(n6671) );
  ANDN U18089 ( .B(n7371), .A(n7372), .Z(n7369) );
  AND U18090 ( .A(a[50]), .B(b[67]), .Z(n7368) );
  XNOR U18091 ( .A(n7373), .B(n6676), .Z(n6678) );
  XOR U18092 ( .A(n7374), .B(n7375), .Z(n6676) );
  ANDN U18093 ( .B(n7376), .A(n7377), .Z(n7374) );
  AND U18094 ( .A(a[51]), .B(b[66]), .Z(n7373) );
  XNOR U18095 ( .A(n7378), .B(n6681), .Z(n6683) );
  XOR U18096 ( .A(n7379), .B(n7380), .Z(n6681) );
  ANDN U18097 ( .B(n7381), .A(n7382), .Z(n7379) );
  AND U18098 ( .A(a[52]), .B(b[65]), .Z(n7378) );
  XNOR U18099 ( .A(n7383), .B(n6686), .Z(n6688) );
  XOR U18100 ( .A(n7384), .B(n7385), .Z(n6686) );
  ANDN U18101 ( .B(n7386), .A(n7387), .Z(n7384) );
  AND U18102 ( .A(a[53]), .B(b[64]), .Z(n7383) );
  XNOR U18103 ( .A(n7388), .B(n6691), .Z(n6693) );
  XOR U18104 ( .A(n7389), .B(n7390), .Z(n6691) );
  ANDN U18105 ( .B(n7391), .A(n7392), .Z(n7389) );
  AND U18106 ( .A(a[54]), .B(b[63]), .Z(n7388) );
  XNOR U18107 ( .A(n7393), .B(n6696), .Z(n6698) );
  XOR U18108 ( .A(n7394), .B(n7395), .Z(n6696) );
  ANDN U18109 ( .B(n7396), .A(n7397), .Z(n7394) );
  AND U18110 ( .A(a[55]), .B(b[62]), .Z(n7393) );
  XNOR U18111 ( .A(n7398), .B(n6701), .Z(n6703) );
  XOR U18112 ( .A(n7399), .B(n7400), .Z(n6701) );
  ANDN U18113 ( .B(n7401), .A(n7402), .Z(n7399) );
  AND U18114 ( .A(a[56]), .B(b[61]), .Z(n7398) );
  XNOR U18115 ( .A(n7403), .B(n6706), .Z(n6708) );
  XOR U18116 ( .A(n7404), .B(n7405), .Z(n6706) );
  ANDN U18117 ( .B(n7406), .A(n7407), .Z(n7404) );
  AND U18118 ( .A(a[57]), .B(b[60]), .Z(n7403) );
  XNOR U18119 ( .A(n7408), .B(n6711), .Z(n6713) );
  XOR U18120 ( .A(n7409), .B(n7410), .Z(n6711) );
  ANDN U18121 ( .B(n7411), .A(n7412), .Z(n7409) );
  AND U18122 ( .A(a[58]), .B(b[59]), .Z(n7408) );
  XNOR U18123 ( .A(n7413), .B(n6716), .Z(n6718) );
  XOR U18124 ( .A(n7414), .B(n7415), .Z(n6716) );
  ANDN U18125 ( .B(n7416), .A(n7417), .Z(n7414) );
  AND U18126 ( .A(a[59]), .B(b[58]), .Z(n7413) );
  XNOR U18127 ( .A(n7418), .B(n6721), .Z(n6723) );
  XOR U18128 ( .A(n7419), .B(n7420), .Z(n6721) );
  ANDN U18129 ( .B(n7421), .A(n7422), .Z(n7419) );
  AND U18130 ( .A(a[60]), .B(b[57]), .Z(n7418) );
  XNOR U18131 ( .A(n7423), .B(n6726), .Z(n6728) );
  XOR U18132 ( .A(n7424), .B(n7425), .Z(n6726) );
  ANDN U18133 ( .B(n7426), .A(n7427), .Z(n7424) );
  AND U18134 ( .A(a[61]), .B(b[56]), .Z(n7423) );
  XNOR U18135 ( .A(n7428), .B(n6731), .Z(n6733) );
  XOR U18136 ( .A(n7429), .B(n7430), .Z(n6731) );
  ANDN U18137 ( .B(n7431), .A(n7432), .Z(n7429) );
  AND U18138 ( .A(a[62]), .B(b[55]), .Z(n7428) );
  XNOR U18139 ( .A(n7433), .B(n6736), .Z(n6738) );
  XOR U18140 ( .A(n7434), .B(n7435), .Z(n6736) );
  ANDN U18141 ( .B(n7436), .A(n7437), .Z(n7434) );
  AND U18142 ( .A(a[63]), .B(b[54]), .Z(n7433) );
  XNOR U18143 ( .A(n7438), .B(n6741), .Z(n6743) );
  XOR U18144 ( .A(n7439), .B(n7440), .Z(n6741) );
  ANDN U18145 ( .B(n7441), .A(n7442), .Z(n7439) );
  AND U18146 ( .A(a[64]), .B(b[53]), .Z(n7438) );
  XNOR U18147 ( .A(n7443), .B(n6746), .Z(n6748) );
  XOR U18148 ( .A(n7444), .B(n7445), .Z(n6746) );
  ANDN U18149 ( .B(n7446), .A(n7447), .Z(n7444) );
  AND U18150 ( .A(a[65]), .B(b[52]), .Z(n7443) );
  XNOR U18151 ( .A(n7448), .B(n6751), .Z(n6753) );
  XOR U18152 ( .A(n7449), .B(n7450), .Z(n6751) );
  ANDN U18153 ( .B(n7451), .A(n7452), .Z(n7449) );
  AND U18154 ( .A(a[66]), .B(b[51]), .Z(n7448) );
  XNOR U18155 ( .A(n7453), .B(n6756), .Z(n6758) );
  XOR U18156 ( .A(n7454), .B(n7455), .Z(n6756) );
  ANDN U18157 ( .B(n7456), .A(n7457), .Z(n7454) );
  AND U18158 ( .A(a[67]), .B(b[50]), .Z(n7453) );
  XNOR U18159 ( .A(n7458), .B(n6761), .Z(n6763) );
  XOR U18160 ( .A(n7459), .B(n7460), .Z(n6761) );
  ANDN U18161 ( .B(n7461), .A(n7462), .Z(n7459) );
  AND U18162 ( .A(a[68]), .B(b[49]), .Z(n7458) );
  XNOR U18163 ( .A(n7463), .B(n6766), .Z(n6768) );
  XOR U18164 ( .A(n7464), .B(n7465), .Z(n6766) );
  ANDN U18165 ( .B(n7466), .A(n7467), .Z(n7464) );
  AND U18166 ( .A(a[69]), .B(b[48]), .Z(n7463) );
  XNOR U18167 ( .A(n7468), .B(n6771), .Z(n6773) );
  XOR U18168 ( .A(n7469), .B(n7470), .Z(n6771) );
  ANDN U18169 ( .B(n7471), .A(n7472), .Z(n7469) );
  AND U18170 ( .A(a[70]), .B(b[47]), .Z(n7468) );
  XNOR U18171 ( .A(n7473), .B(n6776), .Z(n6778) );
  XOR U18172 ( .A(n7474), .B(n7475), .Z(n6776) );
  ANDN U18173 ( .B(n7476), .A(n7477), .Z(n7474) );
  AND U18174 ( .A(a[71]), .B(b[46]), .Z(n7473) );
  XNOR U18175 ( .A(n7478), .B(n6781), .Z(n6783) );
  XOR U18176 ( .A(n7479), .B(n7480), .Z(n6781) );
  ANDN U18177 ( .B(n7481), .A(n7482), .Z(n7479) );
  AND U18178 ( .A(a[72]), .B(b[45]), .Z(n7478) );
  XNOR U18179 ( .A(n7483), .B(n6786), .Z(n6788) );
  XOR U18180 ( .A(n7484), .B(n7485), .Z(n6786) );
  ANDN U18181 ( .B(n7486), .A(n7487), .Z(n7484) );
  AND U18182 ( .A(a[73]), .B(b[44]), .Z(n7483) );
  XNOR U18183 ( .A(n7488), .B(n6791), .Z(n6793) );
  XOR U18184 ( .A(n7489), .B(n7490), .Z(n6791) );
  ANDN U18185 ( .B(n7491), .A(n7492), .Z(n7489) );
  AND U18186 ( .A(a[74]), .B(b[43]), .Z(n7488) );
  XNOR U18187 ( .A(n7493), .B(n6796), .Z(n6798) );
  XOR U18188 ( .A(n7494), .B(n7495), .Z(n6796) );
  ANDN U18189 ( .B(n7496), .A(n7497), .Z(n7494) );
  AND U18190 ( .A(a[75]), .B(b[42]), .Z(n7493) );
  XNOR U18191 ( .A(n7498), .B(n6801), .Z(n6803) );
  XOR U18192 ( .A(n7499), .B(n7500), .Z(n6801) );
  ANDN U18193 ( .B(n7501), .A(n7502), .Z(n7499) );
  AND U18194 ( .A(a[76]), .B(b[41]), .Z(n7498) );
  XNOR U18195 ( .A(n7503), .B(n6806), .Z(n6808) );
  XOR U18196 ( .A(n7504), .B(n7505), .Z(n6806) );
  ANDN U18197 ( .B(n7506), .A(n7507), .Z(n7504) );
  AND U18198 ( .A(a[77]), .B(b[40]), .Z(n7503) );
  XNOR U18199 ( .A(n7508), .B(n6811), .Z(n6813) );
  XOR U18200 ( .A(n7509), .B(n7510), .Z(n6811) );
  ANDN U18201 ( .B(n7511), .A(n7512), .Z(n7509) );
  AND U18202 ( .A(a[78]), .B(b[39]), .Z(n7508) );
  XNOR U18203 ( .A(n7513), .B(n6816), .Z(n6818) );
  XOR U18204 ( .A(n7514), .B(n7515), .Z(n6816) );
  ANDN U18205 ( .B(n7516), .A(n7517), .Z(n7514) );
  AND U18206 ( .A(a[79]), .B(b[38]), .Z(n7513) );
  XNOR U18207 ( .A(n7518), .B(n6821), .Z(n6823) );
  XOR U18208 ( .A(n7519), .B(n7520), .Z(n6821) );
  ANDN U18209 ( .B(n7521), .A(n7522), .Z(n7519) );
  AND U18210 ( .A(a[80]), .B(b[37]), .Z(n7518) );
  XNOR U18211 ( .A(n7523), .B(n6826), .Z(n6828) );
  XOR U18212 ( .A(n7524), .B(n7525), .Z(n6826) );
  ANDN U18213 ( .B(n7526), .A(n7527), .Z(n7524) );
  AND U18214 ( .A(a[81]), .B(b[36]), .Z(n7523) );
  XNOR U18215 ( .A(n7528), .B(n6831), .Z(n6833) );
  XOR U18216 ( .A(n7529), .B(n7530), .Z(n6831) );
  ANDN U18217 ( .B(n7531), .A(n7532), .Z(n7529) );
  AND U18218 ( .A(a[82]), .B(b[35]), .Z(n7528) );
  XNOR U18219 ( .A(n7533), .B(n6836), .Z(n6838) );
  XOR U18220 ( .A(n7534), .B(n7535), .Z(n6836) );
  ANDN U18221 ( .B(n7536), .A(n7537), .Z(n7534) );
  AND U18222 ( .A(a[83]), .B(b[34]), .Z(n7533) );
  XNOR U18223 ( .A(n7538), .B(n6841), .Z(n6843) );
  XOR U18224 ( .A(n7539), .B(n7540), .Z(n6841) );
  ANDN U18225 ( .B(n7541), .A(n7542), .Z(n7539) );
  AND U18226 ( .A(a[84]), .B(b[33]), .Z(n7538) );
  XNOR U18227 ( .A(n7543), .B(n6846), .Z(n6848) );
  XOR U18228 ( .A(n7544), .B(n7545), .Z(n6846) );
  ANDN U18229 ( .B(n7546), .A(n7547), .Z(n7544) );
  AND U18230 ( .A(a[85]), .B(b[32]), .Z(n7543) );
  XNOR U18231 ( .A(n7548), .B(n6851), .Z(n6853) );
  XOR U18232 ( .A(n7549), .B(n7550), .Z(n6851) );
  ANDN U18233 ( .B(n7551), .A(n7552), .Z(n7549) );
  AND U18234 ( .A(a[86]), .B(b[31]), .Z(n7548) );
  XNOR U18235 ( .A(n7553), .B(n6856), .Z(n6858) );
  XOR U18236 ( .A(n7554), .B(n7555), .Z(n6856) );
  ANDN U18237 ( .B(n7556), .A(n7557), .Z(n7554) );
  AND U18238 ( .A(a[87]), .B(b[30]), .Z(n7553) );
  XNOR U18239 ( .A(n7558), .B(n6861), .Z(n6863) );
  XOR U18240 ( .A(n7559), .B(n7560), .Z(n6861) );
  ANDN U18241 ( .B(n7561), .A(n7562), .Z(n7559) );
  AND U18242 ( .A(a[88]), .B(b[29]), .Z(n7558) );
  XNOR U18243 ( .A(n7563), .B(n6866), .Z(n6868) );
  XOR U18244 ( .A(n7564), .B(n7565), .Z(n6866) );
  ANDN U18245 ( .B(n7566), .A(n7567), .Z(n7564) );
  AND U18246 ( .A(a[89]), .B(b[28]), .Z(n7563) );
  XNOR U18247 ( .A(n7568), .B(n6871), .Z(n6873) );
  XOR U18248 ( .A(n7569), .B(n7570), .Z(n6871) );
  ANDN U18249 ( .B(n7571), .A(n7572), .Z(n7569) );
  AND U18250 ( .A(a[90]), .B(b[27]), .Z(n7568) );
  XNOR U18251 ( .A(n7573), .B(n6876), .Z(n6878) );
  XOR U18252 ( .A(n7574), .B(n7575), .Z(n6876) );
  ANDN U18253 ( .B(n7576), .A(n7577), .Z(n7574) );
  AND U18254 ( .A(a[91]), .B(b[26]), .Z(n7573) );
  XNOR U18255 ( .A(n7578), .B(n6881), .Z(n6883) );
  XOR U18256 ( .A(n7579), .B(n7580), .Z(n6881) );
  ANDN U18257 ( .B(n7581), .A(n7582), .Z(n7579) );
  AND U18258 ( .A(a[92]), .B(b[25]), .Z(n7578) );
  XNOR U18259 ( .A(n7583), .B(n6886), .Z(n6888) );
  XOR U18260 ( .A(n7584), .B(n7585), .Z(n6886) );
  ANDN U18261 ( .B(n7586), .A(n7587), .Z(n7584) );
  AND U18262 ( .A(a[93]), .B(b[24]), .Z(n7583) );
  XNOR U18263 ( .A(n7588), .B(n6891), .Z(n6893) );
  XOR U18264 ( .A(n7589), .B(n7590), .Z(n6891) );
  ANDN U18265 ( .B(n7591), .A(n7592), .Z(n7589) );
  AND U18266 ( .A(a[94]), .B(b[23]), .Z(n7588) );
  XNOR U18267 ( .A(n7593), .B(n6896), .Z(n6898) );
  XOR U18268 ( .A(n7594), .B(n7595), .Z(n6896) );
  ANDN U18269 ( .B(n7596), .A(n7597), .Z(n7594) );
  AND U18270 ( .A(a[95]), .B(b[22]), .Z(n7593) );
  XNOR U18271 ( .A(n7598), .B(n6901), .Z(n6903) );
  XOR U18272 ( .A(n7599), .B(n7600), .Z(n6901) );
  ANDN U18273 ( .B(n7601), .A(n7602), .Z(n7599) );
  AND U18274 ( .A(a[96]), .B(b[21]), .Z(n7598) );
  XNOR U18275 ( .A(n7603), .B(n6906), .Z(n6908) );
  XOR U18276 ( .A(n7604), .B(n7605), .Z(n6906) );
  ANDN U18277 ( .B(n7606), .A(n7607), .Z(n7604) );
  AND U18278 ( .A(a[97]), .B(b[20]), .Z(n7603) );
  XNOR U18279 ( .A(n7608), .B(n6911), .Z(n6913) );
  XOR U18280 ( .A(n7609), .B(n7610), .Z(n6911) );
  ANDN U18281 ( .B(n7611), .A(n7612), .Z(n7609) );
  AND U18282 ( .A(a[98]), .B(b[19]), .Z(n7608) );
  XNOR U18283 ( .A(n7613), .B(n6916), .Z(n6918) );
  XOR U18284 ( .A(n7614), .B(n7615), .Z(n6916) );
  ANDN U18285 ( .B(n7616), .A(n7617), .Z(n7614) );
  AND U18286 ( .A(a[99]), .B(b[18]), .Z(n7613) );
  XNOR U18287 ( .A(n7618), .B(n6921), .Z(n6923) );
  XOR U18288 ( .A(n7619), .B(n7620), .Z(n6921) );
  ANDN U18289 ( .B(n7621), .A(n7622), .Z(n7619) );
  AND U18290 ( .A(b[17]), .B(a[100]), .Z(n7618) );
  XNOR U18291 ( .A(n7623), .B(n6926), .Z(n6928) );
  XOR U18292 ( .A(n7624), .B(n7625), .Z(n6926) );
  ANDN U18293 ( .B(n7626), .A(n7627), .Z(n7624) );
  AND U18294 ( .A(b[16]), .B(a[101]), .Z(n7623) );
  XNOR U18295 ( .A(n7628), .B(n6931), .Z(n6933) );
  XOR U18296 ( .A(n7629), .B(n7630), .Z(n6931) );
  ANDN U18297 ( .B(n7631), .A(n7632), .Z(n7629) );
  AND U18298 ( .A(b[15]), .B(a[102]), .Z(n7628) );
  XNOR U18299 ( .A(n7633), .B(n6936), .Z(n6938) );
  XOR U18300 ( .A(n7634), .B(n7635), .Z(n6936) );
  ANDN U18301 ( .B(n7636), .A(n7637), .Z(n7634) );
  AND U18302 ( .A(b[14]), .B(a[103]), .Z(n7633) );
  XNOR U18303 ( .A(n7638), .B(n6941), .Z(n6943) );
  XOR U18304 ( .A(n7639), .B(n7640), .Z(n6941) );
  ANDN U18305 ( .B(n7641), .A(n7642), .Z(n7639) );
  AND U18306 ( .A(b[13]), .B(a[104]), .Z(n7638) );
  XNOR U18307 ( .A(n7643), .B(n6946), .Z(n6948) );
  XOR U18308 ( .A(n7644), .B(n7645), .Z(n6946) );
  ANDN U18309 ( .B(n7646), .A(n7647), .Z(n7644) );
  AND U18310 ( .A(b[12]), .B(a[105]), .Z(n7643) );
  XNOR U18311 ( .A(n7648), .B(n6951), .Z(n6953) );
  XOR U18312 ( .A(n7649), .B(n7650), .Z(n6951) );
  ANDN U18313 ( .B(n7651), .A(n7652), .Z(n7649) );
  AND U18314 ( .A(b[11]), .B(a[106]), .Z(n7648) );
  XNOR U18315 ( .A(n7653), .B(n6956), .Z(n6958) );
  XOR U18316 ( .A(n7654), .B(n7655), .Z(n6956) );
  ANDN U18317 ( .B(n7656), .A(n7657), .Z(n7654) );
  AND U18318 ( .A(b[10]), .B(a[107]), .Z(n7653) );
  XNOR U18319 ( .A(n7658), .B(n6961), .Z(n6963) );
  XOR U18320 ( .A(n7659), .B(n7660), .Z(n6961) );
  ANDN U18321 ( .B(n7661), .A(n7662), .Z(n7659) );
  AND U18322 ( .A(b[9]), .B(a[108]), .Z(n7658) );
  XNOR U18323 ( .A(n7663), .B(n6966), .Z(n6968) );
  XOR U18324 ( .A(n7664), .B(n7665), .Z(n6966) );
  ANDN U18325 ( .B(n7666), .A(n7667), .Z(n7664) );
  AND U18326 ( .A(b[8]), .B(a[109]), .Z(n7663) );
  XNOR U18327 ( .A(n7668), .B(n6971), .Z(n6973) );
  XOR U18328 ( .A(n7669), .B(n7670), .Z(n6971) );
  ANDN U18329 ( .B(n7671), .A(n7672), .Z(n7669) );
  AND U18330 ( .A(b[7]), .B(a[110]), .Z(n7668) );
  XNOR U18331 ( .A(n7673), .B(n6976), .Z(n6978) );
  XOR U18332 ( .A(n7674), .B(n7675), .Z(n6976) );
  ANDN U18333 ( .B(n7676), .A(n7677), .Z(n7674) );
  AND U18334 ( .A(b[6]), .B(a[111]), .Z(n7673) );
  XNOR U18335 ( .A(n7678), .B(n6981), .Z(n6983) );
  XOR U18336 ( .A(n7679), .B(n7680), .Z(n6981) );
  ANDN U18337 ( .B(n7681), .A(n7682), .Z(n7679) );
  AND U18338 ( .A(b[5]), .B(a[112]), .Z(n7678) );
  XNOR U18339 ( .A(n7683), .B(n6986), .Z(n6988) );
  XOR U18340 ( .A(n7684), .B(n7685), .Z(n6986) );
  ANDN U18341 ( .B(n7686), .A(n7687), .Z(n7684) );
  AND U18342 ( .A(b[4]), .B(a[113]), .Z(n7683) );
  XNOR U18343 ( .A(n7688), .B(n7689), .Z(n7000) );
  NANDN U18344 ( .A(n7690), .B(n7691), .Z(n7689) );
  XNOR U18345 ( .A(n7692), .B(n6991), .Z(n6993) );
  XNOR U18346 ( .A(n7693), .B(n7694), .Z(n6991) );
  AND U18347 ( .A(n7695), .B(n7696), .Z(n7693) );
  AND U18348 ( .A(b[3]), .B(a[114]), .Z(n7692) );
  NAND U18349 ( .A(a[117]), .B(b[0]), .Z(n6306) );
  XNOR U18350 ( .A(n7006), .B(n7007), .Z(c[116]) );
  XNOR U18351 ( .A(n7690), .B(n7691), .Z(n7007) );
  XOR U18352 ( .A(n7688), .B(n7697), .Z(n7691) );
  NAND U18353 ( .A(b[1]), .B(a[115]), .Z(n7697) );
  XOR U18354 ( .A(n7696), .B(n7698), .Z(n7690) );
  XOR U18355 ( .A(n7688), .B(n7695), .Z(n7698) );
  XNOR U18356 ( .A(n7699), .B(n7694), .Z(n7695) );
  AND U18357 ( .A(b[2]), .B(a[114]), .Z(n7699) );
  NANDN U18358 ( .A(n7700), .B(n7701), .Z(n7688) );
  XOR U18359 ( .A(n7694), .B(n7686), .Z(n7702) );
  XNOR U18360 ( .A(n7685), .B(n7681), .Z(n7703) );
  XNOR U18361 ( .A(n7680), .B(n7676), .Z(n7704) );
  XNOR U18362 ( .A(n7675), .B(n7671), .Z(n7705) );
  XNOR U18363 ( .A(n7670), .B(n7666), .Z(n7706) );
  XNOR U18364 ( .A(n7665), .B(n7661), .Z(n7707) );
  XNOR U18365 ( .A(n7660), .B(n7656), .Z(n7708) );
  XNOR U18366 ( .A(n7655), .B(n7651), .Z(n7709) );
  XNOR U18367 ( .A(n7650), .B(n7646), .Z(n7710) );
  XNOR U18368 ( .A(n7645), .B(n7641), .Z(n7711) );
  XNOR U18369 ( .A(n7640), .B(n7636), .Z(n7712) );
  XNOR U18370 ( .A(n7635), .B(n7631), .Z(n7713) );
  XNOR U18371 ( .A(n7630), .B(n7626), .Z(n7714) );
  XNOR U18372 ( .A(n7625), .B(n7621), .Z(n7715) );
  XNOR U18373 ( .A(n7620), .B(n7616), .Z(n7716) );
  XNOR U18374 ( .A(n7615), .B(n7611), .Z(n7717) );
  XNOR U18375 ( .A(n7610), .B(n7606), .Z(n7718) );
  XNOR U18376 ( .A(n7605), .B(n7601), .Z(n7719) );
  XNOR U18377 ( .A(n7600), .B(n7596), .Z(n7720) );
  XNOR U18378 ( .A(n7595), .B(n7591), .Z(n7721) );
  XNOR U18379 ( .A(n7590), .B(n7586), .Z(n7722) );
  XNOR U18380 ( .A(n7585), .B(n7581), .Z(n7723) );
  XNOR U18381 ( .A(n7580), .B(n7576), .Z(n7724) );
  XNOR U18382 ( .A(n7575), .B(n7571), .Z(n7725) );
  XNOR U18383 ( .A(n7570), .B(n7566), .Z(n7726) );
  XNOR U18384 ( .A(n7565), .B(n7561), .Z(n7727) );
  XNOR U18385 ( .A(n7560), .B(n7556), .Z(n7728) );
  XNOR U18386 ( .A(n7555), .B(n7551), .Z(n7729) );
  XNOR U18387 ( .A(n7550), .B(n7546), .Z(n7730) );
  XNOR U18388 ( .A(n7545), .B(n7541), .Z(n7731) );
  XNOR U18389 ( .A(n7540), .B(n7536), .Z(n7732) );
  XNOR U18390 ( .A(n7535), .B(n7531), .Z(n7733) );
  XNOR U18391 ( .A(n7530), .B(n7526), .Z(n7734) );
  XNOR U18392 ( .A(n7525), .B(n7521), .Z(n7735) );
  XNOR U18393 ( .A(n7520), .B(n7516), .Z(n7736) );
  XNOR U18394 ( .A(n7515), .B(n7511), .Z(n7737) );
  XNOR U18395 ( .A(n7510), .B(n7506), .Z(n7738) );
  XNOR U18396 ( .A(n7505), .B(n7501), .Z(n7739) );
  XNOR U18397 ( .A(n7500), .B(n7496), .Z(n7740) );
  XNOR U18398 ( .A(n7495), .B(n7491), .Z(n7741) );
  XNOR U18399 ( .A(n7490), .B(n7486), .Z(n7742) );
  XNOR U18400 ( .A(n7485), .B(n7481), .Z(n7743) );
  XNOR U18401 ( .A(n7480), .B(n7476), .Z(n7744) );
  XNOR U18402 ( .A(n7475), .B(n7471), .Z(n7745) );
  XNOR U18403 ( .A(n7470), .B(n7466), .Z(n7746) );
  XNOR U18404 ( .A(n7465), .B(n7461), .Z(n7747) );
  XNOR U18405 ( .A(n7460), .B(n7456), .Z(n7748) );
  XNOR U18406 ( .A(n7455), .B(n7451), .Z(n7749) );
  XNOR U18407 ( .A(n7450), .B(n7446), .Z(n7750) );
  XNOR U18408 ( .A(n7445), .B(n7441), .Z(n7751) );
  XNOR U18409 ( .A(n7440), .B(n7436), .Z(n7752) );
  XNOR U18410 ( .A(n7435), .B(n7431), .Z(n7753) );
  XNOR U18411 ( .A(n7430), .B(n7426), .Z(n7754) );
  XNOR U18412 ( .A(n7425), .B(n7421), .Z(n7755) );
  XNOR U18413 ( .A(n7420), .B(n7416), .Z(n7756) );
  XNOR U18414 ( .A(n7415), .B(n7411), .Z(n7757) );
  XNOR U18415 ( .A(n7410), .B(n7406), .Z(n7758) );
  XNOR U18416 ( .A(n7405), .B(n7401), .Z(n7759) );
  XNOR U18417 ( .A(n7400), .B(n7396), .Z(n7760) );
  XNOR U18418 ( .A(n7395), .B(n7391), .Z(n7761) );
  XNOR U18419 ( .A(n7390), .B(n7386), .Z(n7762) );
  XNOR U18420 ( .A(n7385), .B(n7381), .Z(n7763) );
  XNOR U18421 ( .A(n7380), .B(n7376), .Z(n7764) );
  XNOR U18422 ( .A(n7375), .B(n7371), .Z(n7765) );
  XNOR U18423 ( .A(n7370), .B(n7366), .Z(n7766) );
  XNOR U18424 ( .A(n7365), .B(n7361), .Z(n7767) );
  XNOR U18425 ( .A(n7360), .B(n7356), .Z(n7768) );
  XNOR U18426 ( .A(n7355), .B(n7351), .Z(n7769) );
  XNOR U18427 ( .A(n7350), .B(n7346), .Z(n7770) );
  XNOR U18428 ( .A(n7345), .B(n7341), .Z(n7771) );
  XNOR U18429 ( .A(n7340), .B(n7336), .Z(n7772) );
  XNOR U18430 ( .A(n7335), .B(n7331), .Z(n7773) );
  XNOR U18431 ( .A(n7330), .B(n7326), .Z(n7774) );
  XNOR U18432 ( .A(n7325), .B(n7321), .Z(n7775) );
  XNOR U18433 ( .A(n7320), .B(n7316), .Z(n7776) );
  XNOR U18434 ( .A(n7315), .B(n7311), .Z(n7777) );
  XNOR U18435 ( .A(n7310), .B(n7306), .Z(n7778) );
  XNOR U18436 ( .A(n7305), .B(n7301), .Z(n7779) );
  XNOR U18437 ( .A(n7300), .B(n7296), .Z(n7780) );
  XNOR U18438 ( .A(n7295), .B(n7291), .Z(n7781) );
  XNOR U18439 ( .A(n7290), .B(n7286), .Z(n7782) );
  XNOR U18440 ( .A(n7285), .B(n7281), .Z(n7783) );
  XNOR U18441 ( .A(n7280), .B(n7276), .Z(n7784) );
  XNOR U18442 ( .A(n7275), .B(n7271), .Z(n7785) );
  XNOR U18443 ( .A(n7270), .B(n7266), .Z(n7786) );
  XNOR U18444 ( .A(n7265), .B(n7261), .Z(n7787) );
  XNOR U18445 ( .A(n7260), .B(n7256), .Z(n7788) );
  XNOR U18446 ( .A(n7255), .B(n7251), .Z(n7789) );
  XNOR U18447 ( .A(n7250), .B(n7246), .Z(n7790) );
  XNOR U18448 ( .A(n7245), .B(n7241), .Z(n7791) );
  XNOR U18449 ( .A(n7240), .B(n7236), .Z(n7792) );
  XNOR U18450 ( .A(n7235), .B(n7231), .Z(n7793) );
  XNOR U18451 ( .A(n7230), .B(n7226), .Z(n7794) );
  XNOR U18452 ( .A(n7225), .B(n7221), .Z(n7795) );
  XNOR U18453 ( .A(n7220), .B(n7216), .Z(n7796) );
  XNOR U18454 ( .A(n7215), .B(n7211), .Z(n7797) );
  XNOR U18455 ( .A(n7210), .B(n7206), .Z(n7798) );
  XNOR U18456 ( .A(n7205), .B(n7201), .Z(n7799) );
  XNOR U18457 ( .A(n7200), .B(n7196), .Z(n7800) );
  XNOR U18458 ( .A(n7195), .B(n7191), .Z(n7801) );
  XNOR U18459 ( .A(n7190), .B(n7186), .Z(n7802) );
  XNOR U18460 ( .A(n7185), .B(n7181), .Z(n7803) );
  XNOR U18461 ( .A(n7180), .B(n7176), .Z(n7804) );
  XNOR U18462 ( .A(n7175), .B(n7171), .Z(n7805) );
  XNOR U18463 ( .A(n7170), .B(n7166), .Z(n7806) );
  XNOR U18464 ( .A(n7165), .B(n7161), .Z(n7807) );
  XNOR U18465 ( .A(n7160), .B(n7156), .Z(n7808) );
  XNOR U18466 ( .A(n7155), .B(n7151), .Z(n7809) );
  XNOR U18467 ( .A(n7150), .B(n7146), .Z(n7810) );
  XNOR U18468 ( .A(n7145), .B(n7141), .Z(n7811) );
  XNOR U18469 ( .A(n7140), .B(n7136), .Z(n7812) );
  XNOR U18470 ( .A(n7135), .B(n7131), .Z(n7813) );
  XNOR U18471 ( .A(n7130), .B(n7126), .Z(n7814) );
  XOR U18472 ( .A(n7815), .B(n7125), .Z(n7126) );
  AND U18473 ( .A(a[0]), .B(b[116]), .Z(n7815) );
  XNOR U18474 ( .A(n7816), .B(n7125), .Z(n7127) );
  XNOR U18475 ( .A(n7817), .B(n7818), .Z(n7125) );
  ANDN U18476 ( .B(n7819), .A(n7820), .Z(n7817) );
  AND U18477 ( .A(a[1]), .B(b[115]), .Z(n7816) );
  XNOR U18478 ( .A(n7821), .B(n7130), .Z(n7132) );
  XOR U18479 ( .A(n7822), .B(n7823), .Z(n7130) );
  ANDN U18480 ( .B(n7824), .A(n7825), .Z(n7822) );
  AND U18481 ( .A(a[2]), .B(b[114]), .Z(n7821) );
  XNOR U18482 ( .A(n7826), .B(n7135), .Z(n7137) );
  XOR U18483 ( .A(n7827), .B(n7828), .Z(n7135) );
  ANDN U18484 ( .B(n7829), .A(n7830), .Z(n7827) );
  AND U18485 ( .A(a[3]), .B(b[113]), .Z(n7826) );
  XNOR U18486 ( .A(n7831), .B(n7140), .Z(n7142) );
  XOR U18487 ( .A(n7832), .B(n7833), .Z(n7140) );
  ANDN U18488 ( .B(n7834), .A(n7835), .Z(n7832) );
  AND U18489 ( .A(a[4]), .B(b[112]), .Z(n7831) );
  XNOR U18490 ( .A(n7836), .B(n7145), .Z(n7147) );
  XOR U18491 ( .A(n7837), .B(n7838), .Z(n7145) );
  ANDN U18492 ( .B(n7839), .A(n7840), .Z(n7837) );
  AND U18493 ( .A(a[5]), .B(b[111]), .Z(n7836) );
  XNOR U18494 ( .A(n7841), .B(n7150), .Z(n7152) );
  XOR U18495 ( .A(n7842), .B(n7843), .Z(n7150) );
  ANDN U18496 ( .B(n7844), .A(n7845), .Z(n7842) );
  AND U18497 ( .A(a[6]), .B(b[110]), .Z(n7841) );
  XNOR U18498 ( .A(n7846), .B(n7155), .Z(n7157) );
  XOR U18499 ( .A(n7847), .B(n7848), .Z(n7155) );
  ANDN U18500 ( .B(n7849), .A(n7850), .Z(n7847) );
  AND U18501 ( .A(a[7]), .B(b[109]), .Z(n7846) );
  XNOR U18502 ( .A(n7851), .B(n7160), .Z(n7162) );
  XOR U18503 ( .A(n7852), .B(n7853), .Z(n7160) );
  ANDN U18504 ( .B(n7854), .A(n7855), .Z(n7852) );
  AND U18505 ( .A(a[8]), .B(b[108]), .Z(n7851) );
  XNOR U18506 ( .A(n7856), .B(n7165), .Z(n7167) );
  XOR U18507 ( .A(n7857), .B(n7858), .Z(n7165) );
  ANDN U18508 ( .B(n7859), .A(n7860), .Z(n7857) );
  AND U18509 ( .A(a[9]), .B(b[107]), .Z(n7856) );
  XNOR U18510 ( .A(n7861), .B(n7170), .Z(n7172) );
  XOR U18511 ( .A(n7862), .B(n7863), .Z(n7170) );
  ANDN U18512 ( .B(n7864), .A(n7865), .Z(n7862) );
  AND U18513 ( .A(a[10]), .B(b[106]), .Z(n7861) );
  XNOR U18514 ( .A(n7866), .B(n7175), .Z(n7177) );
  XOR U18515 ( .A(n7867), .B(n7868), .Z(n7175) );
  ANDN U18516 ( .B(n7869), .A(n7870), .Z(n7867) );
  AND U18517 ( .A(a[11]), .B(b[105]), .Z(n7866) );
  XNOR U18518 ( .A(n7871), .B(n7180), .Z(n7182) );
  XOR U18519 ( .A(n7872), .B(n7873), .Z(n7180) );
  ANDN U18520 ( .B(n7874), .A(n7875), .Z(n7872) );
  AND U18521 ( .A(a[12]), .B(b[104]), .Z(n7871) );
  XNOR U18522 ( .A(n7876), .B(n7185), .Z(n7187) );
  XOR U18523 ( .A(n7877), .B(n7878), .Z(n7185) );
  ANDN U18524 ( .B(n7879), .A(n7880), .Z(n7877) );
  AND U18525 ( .A(a[13]), .B(b[103]), .Z(n7876) );
  XNOR U18526 ( .A(n7881), .B(n7190), .Z(n7192) );
  XOR U18527 ( .A(n7882), .B(n7883), .Z(n7190) );
  ANDN U18528 ( .B(n7884), .A(n7885), .Z(n7882) );
  AND U18529 ( .A(a[14]), .B(b[102]), .Z(n7881) );
  XNOR U18530 ( .A(n7886), .B(n7195), .Z(n7197) );
  XOR U18531 ( .A(n7887), .B(n7888), .Z(n7195) );
  ANDN U18532 ( .B(n7889), .A(n7890), .Z(n7887) );
  AND U18533 ( .A(a[15]), .B(b[101]), .Z(n7886) );
  XNOR U18534 ( .A(n7891), .B(n7200), .Z(n7202) );
  XOR U18535 ( .A(n7892), .B(n7893), .Z(n7200) );
  ANDN U18536 ( .B(n7894), .A(n7895), .Z(n7892) );
  AND U18537 ( .A(a[16]), .B(b[100]), .Z(n7891) );
  XNOR U18538 ( .A(n7896), .B(n7205), .Z(n7207) );
  XOR U18539 ( .A(n7897), .B(n7898), .Z(n7205) );
  ANDN U18540 ( .B(n7899), .A(n7900), .Z(n7897) );
  AND U18541 ( .A(a[17]), .B(b[99]), .Z(n7896) );
  XNOR U18542 ( .A(n7901), .B(n7210), .Z(n7212) );
  XOR U18543 ( .A(n7902), .B(n7903), .Z(n7210) );
  ANDN U18544 ( .B(n7904), .A(n7905), .Z(n7902) );
  AND U18545 ( .A(a[18]), .B(b[98]), .Z(n7901) );
  XNOR U18546 ( .A(n7906), .B(n7215), .Z(n7217) );
  XOR U18547 ( .A(n7907), .B(n7908), .Z(n7215) );
  ANDN U18548 ( .B(n7909), .A(n7910), .Z(n7907) );
  AND U18549 ( .A(a[19]), .B(b[97]), .Z(n7906) );
  XNOR U18550 ( .A(n7911), .B(n7220), .Z(n7222) );
  XOR U18551 ( .A(n7912), .B(n7913), .Z(n7220) );
  ANDN U18552 ( .B(n7914), .A(n7915), .Z(n7912) );
  AND U18553 ( .A(a[20]), .B(b[96]), .Z(n7911) );
  XNOR U18554 ( .A(n7916), .B(n7225), .Z(n7227) );
  XOR U18555 ( .A(n7917), .B(n7918), .Z(n7225) );
  ANDN U18556 ( .B(n7919), .A(n7920), .Z(n7917) );
  AND U18557 ( .A(a[21]), .B(b[95]), .Z(n7916) );
  XNOR U18558 ( .A(n7921), .B(n7230), .Z(n7232) );
  XOR U18559 ( .A(n7922), .B(n7923), .Z(n7230) );
  ANDN U18560 ( .B(n7924), .A(n7925), .Z(n7922) );
  AND U18561 ( .A(a[22]), .B(b[94]), .Z(n7921) );
  XNOR U18562 ( .A(n7926), .B(n7235), .Z(n7237) );
  XOR U18563 ( .A(n7927), .B(n7928), .Z(n7235) );
  ANDN U18564 ( .B(n7929), .A(n7930), .Z(n7927) );
  AND U18565 ( .A(a[23]), .B(b[93]), .Z(n7926) );
  XNOR U18566 ( .A(n7931), .B(n7240), .Z(n7242) );
  XOR U18567 ( .A(n7932), .B(n7933), .Z(n7240) );
  ANDN U18568 ( .B(n7934), .A(n7935), .Z(n7932) );
  AND U18569 ( .A(a[24]), .B(b[92]), .Z(n7931) );
  XNOR U18570 ( .A(n7936), .B(n7245), .Z(n7247) );
  XOR U18571 ( .A(n7937), .B(n7938), .Z(n7245) );
  ANDN U18572 ( .B(n7939), .A(n7940), .Z(n7937) );
  AND U18573 ( .A(a[25]), .B(b[91]), .Z(n7936) );
  XNOR U18574 ( .A(n7941), .B(n7250), .Z(n7252) );
  XOR U18575 ( .A(n7942), .B(n7943), .Z(n7250) );
  ANDN U18576 ( .B(n7944), .A(n7945), .Z(n7942) );
  AND U18577 ( .A(a[26]), .B(b[90]), .Z(n7941) );
  XNOR U18578 ( .A(n7946), .B(n7255), .Z(n7257) );
  XOR U18579 ( .A(n7947), .B(n7948), .Z(n7255) );
  ANDN U18580 ( .B(n7949), .A(n7950), .Z(n7947) );
  AND U18581 ( .A(a[27]), .B(b[89]), .Z(n7946) );
  XNOR U18582 ( .A(n7951), .B(n7260), .Z(n7262) );
  XOR U18583 ( .A(n7952), .B(n7953), .Z(n7260) );
  ANDN U18584 ( .B(n7954), .A(n7955), .Z(n7952) );
  AND U18585 ( .A(a[28]), .B(b[88]), .Z(n7951) );
  XNOR U18586 ( .A(n7956), .B(n7265), .Z(n7267) );
  XOR U18587 ( .A(n7957), .B(n7958), .Z(n7265) );
  ANDN U18588 ( .B(n7959), .A(n7960), .Z(n7957) );
  AND U18589 ( .A(a[29]), .B(b[87]), .Z(n7956) );
  XNOR U18590 ( .A(n7961), .B(n7270), .Z(n7272) );
  XOR U18591 ( .A(n7962), .B(n7963), .Z(n7270) );
  ANDN U18592 ( .B(n7964), .A(n7965), .Z(n7962) );
  AND U18593 ( .A(a[30]), .B(b[86]), .Z(n7961) );
  XNOR U18594 ( .A(n7966), .B(n7275), .Z(n7277) );
  XOR U18595 ( .A(n7967), .B(n7968), .Z(n7275) );
  ANDN U18596 ( .B(n7969), .A(n7970), .Z(n7967) );
  AND U18597 ( .A(a[31]), .B(b[85]), .Z(n7966) );
  XNOR U18598 ( .A(n7971), .B(n7280), .Z(n7282) );
  XOR U18599 ( .A(n7972), .B(n7973), .Z(n7280) );
  ANDN U18600 ( .B(n7974), .A(n7975), .Z(n7972) );
  AND U18601 ( .A(a[32]), .B(b[84]), .Z(n7971) );
  XNOR U18602 ( .A(n7976), .B(n7285), .Z(n7287) );
  XOR U18603 ( .A(n7977), .B(n7978), .Z(n7285) );
  ANDN U18604 ( .B(n7979), .A(n7980), .Z(n7977) );
  AND U18605 ( .A(a[33]), .B(b[83]), .Z(n7976) );
  XNOR U18606 ( .A(n7981), .B(n7290), .Z(n7292) );
  XOR U18607 ( .A(n7982), .B(n7983), .Z(n7290) );
  ANDN U18608 ( .B(n7984), .A(n7985), .Z(n7982) );
  AND U18609 ( .A(a[34]), .B(b[82]), .Z(n7981) );
  XNOR U18610 ( .A(n7986), .B(n7295), .Z(n7297) );
  XOR U18611 ( .A(n7987), .B(n7988), .Z(n7295) );
  ANDN U18612 ( .B(n7989), .A(n7990), .Z(n7987) );
  AND U18613 ( .A(a[35]), .B(b[81]), .Z(n7986) );
  XNOR U18614 ( .A(n7991), .B(n7300), .Z(n7302) );
  XOR U18615 ( .A(n7992), .B(n7993), .Z(n7300) );
  ANDN U18616 ( .B(n7994), .A(n7995), .Z(n7992) );
  AND U18617 ( .A(a[36]), .B(b[80]), .Z(n7991) );
  XNOR U18618 ( .A(n7996), .B(n7305), .Z(n7307) );
  XOR U18619 ( .A(n7997), .B(n7998), .Z(n7305) );
  ANDN U18620 ( .B(n7999), .A(n8000), .Z(n7997) );
  AND U18621 ( .A(a[37]), .B(b[79]), .Z(n7996) );
  XNOR U18622 ( .A(n8001), .B(n7310), .Z(n7312) );
  XOR U18623 ( .A(n8002), .B(n8003), .Z(n7310) );
  ANDN U18624 ( .B(n8004), .A(n8005), .Z(n8002) );
  AND U18625 ( .A(a[38]), .B(b[78]), .Z(n8001) );
  XNOR U18626 ( .A(n8006), .B(n7315), .Z(n7317) );
  XOR U18627 ( .A(n8007), .B(n8008), .Z(n7315) );
  ANDN U18628 ( .B(n8009), .A(n8010), .Z(n8007) );
  AND U18629 ( .A(a[39]), .B(b[77]), .Z(n8006) );
  XNOR U18630 ( .A(n8011), .B(n7320), .Z(n7322) );
  XOR U18631 ( .A(n8012), .B(n8013), .Z(n7320) );
  ANDN U18632 ( .B(n8014), .A(n8015), .Z(n8012) );
  AND U18633 ( .A(a[40]), .B(b[76]), .Z(n8011) );
  XNOR U18634 ( .A(n8016), .B(n7325), .Z(n7327) );
  XOR U18635 ( .A(n8017), .B(n8018), .Z(n7325) );
  ANDN U18636 ( .B(n8019), .A(n8020), .Z(n8017) );
  AND U18637 ( .A(a[41]), .B(b[75]), .Z(n8016) );
  XNOR U18638 ( .A(n8021), .B(n7330), .Z(n7332) );
  XOR U18639 ( .A(n8022), .B(n8023), .Z(n7330) );
  ANDN U18640 ( .B(n8024), .A(n8025), .Z(n8022) );
  AND U18641 ( .A(a[42]), .B(b[74]), .Z(n8021) );
  XNOR U18642 ( .A(n8026), .B(n7335), .Z(n7337) );
  XOR U18643 ( .A(n8027), .B(n8028), .Z(n7335) );
  ANDN U18644 ( .B(n8029), .A(n8030), .Z(n8027) );
  AND U18645 ( .A(a[43]), .B(b[73]), .Z(n8026) );
  XNOR U18646 ( .A(n8031), .B(n7340), .Z(n7342) );
  XOR U18647 ( .A(n8032), .B(n8033), .Z(n7340) );
  ANDN U18648 ( .B(n8034), .A(n8035), .Z(n8032) );
  AND U18649 ( .A(a[44]), .B(b[72]), .Z(n8031) );
  XNOR U18650 ( .A(n8036), .B(n7345), .Z(n7347) );
  XOR U18651 ( .A(n8037), .B(n8038), .Z(n7345) );
  ANDN U18652 ( .B(n8039), .A(n8040), .Z(n8037) );
  AND U18653 ( .A(a[45]), .B(b[71]), .Z(n8036) );
  XNOR U18654 ( .A(n8041), .B(n7350), .Z(n7352) );
  XOR U18655 ( .A(n8042), .B(n8043), .Z(n7350) );
  ANDN U18656 ( .B(n8044), .A(n8045), .Z(n8042) );
  AND U18657 ( .A(a[46]), .B(b[70]), .Z(n8041) );
  XNOR U18658 ( .A(n8046), .B(n7355), .Z(n7357) );
  XOR U18659 ( .A(n8047), .B(n8048), .Z(n7355) );
  ANDN U18660 ( .B(n8049), .A(n8050), .Z(n8047) );
  AND U18661 ( .A(a[47]), .B(b[69]), .Z(n8046) );
  XNOR U18662 ( .A(n8051), .B(n7360), .Z(n7362) );
  XOR U18663 ( .A(n8052), .B(n8053), .Z(n7360) );
  ANDN U18664 ( .B(n8054), .A(n8055), .Z(n8052) );
  AND U18665 ( .A(a[48]), .B(b[68]), .Z(n8051) );
  XNOR U18666 ( .A(n8056), .B(n7365), .Z(n7367) );
  XOR U18667 ( .A(n8057), .B(n8058), .Z(n7365) );
  ANDN U18668 ( .B(n8059), .A(n8060), .Z(n8057) );
  AND U18669 ( .A(a[49]), .B(b[67]), .Z(n8056) );
  XNOR U18670 ( .A(n8061), .B(n7370), .Z(n7372) );
  XOR U18671 ( .A(n8062), .B(n8063), .Z(n7370) );
  ANDN U18672 ( .B(n8064), .A(n8065), .Z(n8062) );
  AND U18673 ( .A(a[50]), .B(b[66]), .Z(n8061) );
  XNOR U18674 ( .A(n8066), .B(n7375), .Z(n7377) );
  XOR U18675 ( .A(n8067), .B(n8068), .Z(n7375) );
  ANDN U18676 ( .B(n8069), .A(n8070), .Z(n8067) );
  AND U18677 ( .A(a[51]), .B(b[65]), .Z(n8066) );
  XNOR U18678 ( .A(n8071), .B(n7380), .Z(n7382) );
  XOR U18679 ( .A(n8072), .B(n8073), .Z(n7380) );
  ANDN U18680 ( .B(n8074), .A(n8075), .Z(n8072) );
  AND U18681 ( .A(a[52]), .B(b[64]), .Z(n8071) );
  XNOR U18682 ( .A(n8076), .B(n7385), .Z(n7387) );
  XOR U18683 ( .A(n8077), .B(n8078), .Z(n7385) );
  ANDN U18684 ( .B(n8079), .A(n8080), .Z(n8077) );
  AND U18685 ( .A(a[53]), .B(b[63]), .Z(n8076) );
  XNOR U18686 ( .A(n8081), .B(n7390), .Z(n7392) );
  XOR U18687 ( .A(n8082), .B(n8083), .Z(n7390) );
  ANDN U18688 ( .B(n8084), .A(n8085), .Z(n8082) );
  AND U18689 ( .A(a[54]), .B(b[62]), .Z(n8081) );
  XNOR U18690 ( .A(n8086), .B(n7395), .Z(n7397) );
  XOR U18691 ( .A(n8087), .B(n8088), .Z(n7395) );
  ANDN U18692 ( .B(n8089), .A(n8090), .Z(n8087) );
  AND U18693 ( .A(a[55]), .B(b[61]), .Z(n8086) );
  XNOR U18694 ( .A(n8091), .B(n7400), .Z(n7402) );
  XOR U18695 ( .A(n8092), .B(n8093), .Z(n7400) );
  ANDN U18696 ( .B(n8094), .A(n8095), .Z(n8092) );
  AND U18697 ( .A(a[56]), .B(b[60]), .Z(n8091) );
  XNOR U18698 ( .A(n8096), .B(n7405), .Z(n7407) );
  XOR U18699 ( .A(n8097), .B(n8098), .Z(n7405) );
  ANDN U18700 ( .B(n8099), .A(n8100), .Z(n8097) );
  AND U18701 ( .A(a[57]), .B(b[59]), .Z(n8096) );
  XNOR U18702 ( .A(n8101), .B(n7410), .Z(n7412) );
  XOR U18703 ( .A(n8102), .B(n8103), .Z(n7410) );
  ANDN U18704 ( .B(n8104), .A(n8105), .Z(n8102) );
  AND U18705 ( .A(a[58]), .B(b[58]), .Z(n8101) );
  XNOR U18706 ( .A(n8106), .B(n7415), .Z(n7417) );
  XOR U18707 ( .A(n8107), .B(n8108), .Z(n7415) );
  ANDN U18708 ( .B(n8109), .A(n8110), .Z(n8107) );
  AND U18709 ( .A(a[59]), .B(b[57]), .Z(n8106) );
  XNOR U18710 ( .A(n8111), .B(n7420), .Z(n7422) );
  XOR U18711 ( .A(n8112), .B(n8113), .Z(n7420) );
  ANDN U18712 ( .B(n8114), .A(n8115), .Z(n8112) );
  AND U18713 ( .A(a[60]), .B(b[56]), .Z(n8111) );
  XNOR U18714 ( .A(n8116), .B(n7425), .Z(n7427) );
  XOR U18715 ( .A(n8117), .B(n8118), .Z(n7425) );
  ANDN U18716 ( .B(n8119), .A(n8120), .Z(n8117) );
  AND U18717 ( .A(a[61]), .B(b[55]), .Z(n8116) );
  XNOR U18718 ( .A(n8121), .B(n7430), .Z(n7432) );
  XOR U18719 ( .A(n8122), .B(n8123), .Z(n7430) );
  ANDN U18720 ( .B(n8124), .A(n8125), .Z(n8122) );
  AND U18721 ( .A(a[62]), .B(b[54]), .Z(n8121) );
  XNOR U18722 ( .A(n8126), .B(n7435), .Z(n7437) );
  XOR U18723 ( .A(n8127), .B(n8128), .Z(n7435) );
  ANDN U18724 ( .B(n8129), .A(n8130), .Z(n8127) );
  AND U18725 ( .A(a[63]), .B(b[53]), .Z(n8126) );
  XNOR U18726 ( .A(n8131), .B(n7440), .Z(n7442) );
  XOR U18727 ( .A(n8132), .B(n8133), .Z(n7440) );
  ANDN U18728 ( .B(n8134), .A(n8135), .Z(n8132) );
  AND U18729 ( .A(a[64]), .B(b[52]), .Z(n8131) );
  XNOR U18730 ( .A(n8136), .B(n7445), .Z(n7447) );
  XOR U18731 ( .A(n8137), .B(n8138), .Z(n7445) );
  ANDN U18732 ( .B(n8139), .A(n8140), .Z(n8137) );
  AND U18733 ( .A(a[65]), .B(b[51]), .Z(n8136) );
  XNOR U18734 ( .A(n8141), .B(n7450), .Z(n7452) );
  XOR U18735 ( .A(n8142), .B(n8143), .Z(n7450) );
  ANDN U18736 ( .B(n8144), .A(n8145), .Z(n8142) );
  AND U18737 ( .A(a[66]), .B(b[50]), .Z(n8141) );
  XNOR U18738 ( .A(n8146), .B(n7455), .Z(n7457) );
  XOR U18739 ( .A(n8147), .B(n8148), .Z(n7455) );
  ANDN U18740 ( .B(n8149), .A(n8150), .Z(n8147) );
  AND U18741 ( .A(a[67]), .B(b[49]), .Z(n8146) );
  XNOR U18742 ( .A(n8151), .B(n7460), .Z(n7462) );
  XOR U18743 ( .A(n8152), .B(n8153), .Z(n7460) );
  ANDN U18744 ( .B(n8154), .A(n8155), .Z(n8152) );
  AND U18745 ( .A(a[68]), .B(b[48]), .Z(n8151) );
  XNOR U18746 ( .A(n8156), .B(n7465), .Z(n7467) );
  XOR U18747 ( .A(n8157), .B(n8158), .Z(n7465) );
  ANDN U18748 ( .B(n8159), .A(n8160), .Z(n8157) );
  AND U18749 ( .A(a[69]), .B(b[47]), .Z(n8156) );
  XNOR U18750 ( .A(n8161), .B(n7470), .Z(n7472) );
  XOR U18751 ( .A(n8162), .B(n8163), .Z(n7470) );
  ANDN U18752 ( .B(n8164), .A(n8165), .Z(n8162) );
  AND U18753 ( .A(a[70]), .B(b[46]), .Z(n8161) );
  XNOR U18754 ( .A(n8166), .B(n7475), .Z(n7477) );
  XOR U18755 ( .A(n8167), .B(n8168), .Z(n7475) );
  ANDN U18756 ( .B(n8169), .A(n8170), .Z(n8167) );
  AND U18757 ( .A(a[71]), .B(b[45]), .Z(n8166) );
  XNOR U18758 ( .A(n8171), .B(n7480), .Z(n7482) );
  XOR U18759 ( .A(n8172), .B(n8173), .Z(n7480) );
  ANDN U18760 ( .B(n8174), .A(n8175), .Z(n8172) );
  AND U18761 ( .A(a[72]), .B(b[44]), .Z(n8171) );
  XNOR U18762 ( .A(n8176), .B(n7485), .Z(n7487) );
  XOR U18763 ( .A(n8177), .B(n8178), .Z(n7485) );
  ANDN U18764 ( .B(n8179), .A(n8180), .Z(n8177) );
  AND U18765 ( .A(a[73]), .B(b[43]), .Z(n8176) );
  XNOR U18766 ( .A(n8181), .B(n7490), .Z(n7492) );
  XOR U18767 ( .A(n8182), .B(n8183), .Z(n7490) );
  ANDN U18768 ( .B(n8184), .A(n8185), .Z(n8182) );
  AND U18769 ( .A(a[74]), .B(b[42]), .Z(n8181) );
  XNOR U18770 ( .A(n8186), .B(n7495), .Z(n7497) );
  XOR U18771 ( .A(n8187), .B(n8188), .Z(n7495) );
  ANDN U18772 ( .B(n8189), .A(n8190), .Z(n8187) );
  AND U18773 ( .A(a[75]), .B(b[41]), .Z(n8186) );
  XNOR U18774 ( .A(n8191), .B(n7500), .Z(n7502) );
  XOR U18775 ( .A(n8192), .B(n8193), .Z(n7500) );
  ANDN U18776 ( .B(n8194), .A(n8195), .Z(n8192) );
  AND U18777 ( .A(a[76]), .B(b[40]), .Z(n8191) );
  XNOR U18778 ( .A(n8196), .B(n7505), .Z(n7507) );
  XOR U18779 ( .A(n8197), .B(n8198), .Z(n7505) );
  ANDN U18780 ( .B(n8199), .A(n8200), .Z(n8197) );
  AND U18781 ( .A(a[77]), .B(b[39]), .Z(n8196) );
  XNOR U18782 ( .A(n8201), .B(n7510), .Z(n7512) );
  XOR U18783 ( .A(n8202), .B(n8203), .Z(n7510) );
  ANDN U18784 ( .B(n8204), .A(n8205), .Z(n8202) );
  AND U18785 ( .A(a[78]), .B(b[38]), .Z(n8201) );
  XNOR U18786 ( .A(n8206), .B(n7515), .Z(n7517) );
  XOR U18787 ( .A(n8207), .B(n8208), .Z(n7515) );
  ANDN U18788 ( .B(n8209), .A(n8210), .Z(n8207) );
  AND U18789 ( .A(a[79]), .B(b[37]), .Z(n8206) );
  XNOR U18790 ( .A(n8211), .B(n7520), .Z(n7522) );
  XOR U18791 ( .A(n8212), .B(n8213), .Z(n7520) );
  ANDN U18792 ( .B(n8214), .A(n8215), .Z(n8212) );
  AND U18793 ( .A(a[80]), .B(b[36]), .Z(n8211) );
  XNOR U18794 ( .A(n8216), .B(n7525), .Z(n7527) );
  XOR U18795 ( .A(n8217), .B(n8218), .Z(n7525) );
  ANDN U18796 ( .B(n8219), .A(n8220), .Z(n8217) );
  AND U18797 ( .A(a[81]), .B(b[35]), .Z(n8216) );
  XNOR U18798 ( .A(n8221), .B(n7530), .Z(n7532) );
  XOR U18799 ( .A(n8222), .B(n8223), .Z(n7530) );
  ANDN U18800 ( .B(n8224), .A(n8225), .Z(n8222) );
  AND U18801 ( .A(a[82]), .B(b[34]), .Z(n8221) );
  XNOR U18802 ( .A(n8226), .B(n7535), .Z(n7537) );
  XOR U18803 ( .A(n8227), .B(n8228), .Z(n7535) );
  ANDN U18804 ( .B(n8229), .A(n8230), .Z(n8227) );
  AND U18805 ( .A(a[83]), .B(b[33]), .Z(n8226) );
  XNOR U18806 ( .A(n8231), .B(n7540), .Z(n7542) );
  XOR U18807 ( .A(n8232), .B(n8233), .Z(n7540) );
  ANDN U18808 ( .B(n8234), .A(n8235), .Z(n8232) );
  AND U18809 ( .A(a[84]), .B(b[32]), .Z(n8231) );
  XNOR U18810 ( .A(n8236), .B(n7545), .Z(n7547) );
  XOR U18811 ( .A(n8237), .B(n8238), .Z(n7545) );
  ANDN U18812 ( .B(n8239), .A(n8240), .Z(n8237) );
  AND U18813 ( .A(a[85]), .B(b[31]), .Z(n8236) );
  XNOR U18814 ( .A(n8241), .B(n7550), .Z(n7552) );
  XOR U18815 ( .A(n8242), .B(n8243), .Z(n7550) );
  ANDN U18816 ( .B(n8244), .A(n8245), .Z(n8242) );
  AND U18817 ( .A(a[86]), .B(b[30]), .Z(n8241) );
  XNOR U18818 ( .A(n8246), .B(n7555), .Z(n7557) );
  XOR U18819 ( .A(n8247), .B(n8248), .Z(n7555) );
  ANDN U18820 ( .B(n8249), .A(n8250), .Z(n8247) );
  AND U18821 ( .A(a[87]), .B(b[29]), .Z(n8246) );
  XNOR U18822 ( .A(n8251), .B(n7560), .Z(n7562) );
  XOR U18823 ( .A(n8252), .B(n8253), .Z(n7560) );
  ANDN U18824 ( .B(n8254), .A(n8255), .Z(n8252) );
  AND U18825 ( .A(a[88]), .B(b[28]), .Z(n8251) );
  XNOR U18826 ( .A(n8256), .B(n7565), .Z(n7567) );
  XOR U18827 ( .A(n8257), .B(n8258), .Z(n7565) );
  ANDN U18828 ( .B(n8259), .A(n8260), .Z(n8257) );
  AND U18829 ( .A(a[89]), .B(b[27]), .Z(n8256) );
  XNOR U18830 ( .A(n8261), .B(n7570), .Z(n7572) );
  XOR U18831 ( .A(n8262), .B(n8263), .Z(n7570) );
  ANDN U18832 ( .B(n8264), .A(n8265), .Z(n8262) );
  AND U18833 ( .A(a[90]), .B(b[26]), .Z(n8261) );
  XNOR U18834 ( .A(n8266), .B(n7575), .Z(n7577) );
  XOR U18835 ( .A(n8267), .B(n8268), .Z(n7575) );
  ANDN U18836 ( .B(n8269), .A(n8270), .Z(n8267) );
  AND U18837 ( .A(a[91]), .B(b[25]), .Z(n8266) );
  XNOR U18838 ( .A(n8271), .B(n7580), .Z(n7582) );
  XOR U18839 ( .A(n8272), .B(n8273), .Z(n7580) );
  ANDN U18840 ( .B(n8274), .A(n8275), .Z(n8272) );
  AND U18841 ( .A(a[92]), .B(b[24]), .Z(n8271) );
  XNOR U18842 ( .A(n8276), .B(n7585), .Z(n7587) );
  XOR U18843 ( .A(n8277), .B(n8278), .Z(n7585) );
  ANDN U18844 ( .B(n8279), .A(n8280), .Z(n8277) );
  AND U18845 ( .A(a[93]), .B(b[23]), .Z(n8276) );
  XNOR U18846 ( .A(n8281), .B(n7590), .Z(n7592) );
  XOR U18847 ( .A(n8282), .B(n8283), .Z(n7590) );
  ANDN U18848 ( .B(n8284), .A(n8285), .Z(n8282) );
  AND U18849 ( .A(a[94]), .B(b[22]), .Z(n8281) );
  XNOR U18850 ( .A(n8286), .B(n7595), .Z(n7597) );
  XOR U18851 ( .A(n8287), .B(n8288), .Z(n7595) );
  ANDN U18852 ( .B(n8289), .A(n8290), .Z(n8287) );
  AND U18853 ( .A(a[95]), .B(b[21]), .Z(n8286) );
  XNOR U18854 ( .A(n8291), .B(n7600), .Z(n7602) );
  XOR U18855 ( .A(n8292), .B(n8293), .Z(n7600) );
  ANDN U18856 ( .B(n8294), .A(n8295), .Z(n8292) );
  AND U18857 ( .A(a[96]), .B(b[20]), .Z(n8291) );
  XNOR U18858 ( .A(n8296), .B(n7605), .Z(n7607) );
  XOR U18859 ( .A(n8297), .B(n8298), .Z(n7605) );
  ANDN U18860 ( .B(n8299), .A(n8300), .Z(n8297) );
  AND U18861 ( .A(a[97]), .B(b[19]), .Z(n8296) );
  XNOR U18862 ( .A(n8301), .B(n7610), .Z(n7612) );
  XOR U18863 ( .A(n8302), .B(n8303), .Z(n7610) );
  ANDN U18864 ( .B(n8304), .A(n8305), .Z(n8302) );
  AND U18865 ( .A(a[98]), .B(b[18]), .Z(n8301) );
  XNOR U18866 ( .A(n8306), .B(n7615), .Z(n7617) );
  XOR U18867 ( .A(n8307), .B(n8308), .Z(n7615) );
  ANDN U18868 ( .B(n8309), .A(n8310), .Z(n8307) );
  AND U18869 ( .A(a[99]), .B(b[17]), .Z(n8306) );
  XNOR U18870 ( .A(n8311), .B(n7620), .Z(n7622) );
  XOR U18871 ( .A(n8312), .B(n8313), .Z(n7620) );
  ANDN U18872 ( .B(n8314), .A(n8315), .Z(n8312) );
  AND U18873 ( .A(b[16]), .B(a[100]), .Z(n8311) );
  XNOR U18874 ( .A(n8316), .B(n7625), .Z(n7627) );
  XOR U18875 ( .A(n8317), .B(n8318), .Z(n7625) );
  ANDN U18876 ( .B(n8319), .A(n8320), .Z(n8317) );
  AND U18877 ( .A(b[15]), .B(a[101]), .Z(n8316) );
  XNOR U18878 ( .A(n8321), .B(n7630), .Z(n7632) );
  XOR U18879 ( .A(n8322), .B(n8323), .Z(n7630) );
  ANDN U18880 ( .B(n8324), .A(n8325), .Z(n8322) );
  AND U18881 ( .A(b[14]), .B(a[102]), .Z(n8321) );
  XNOR U18882 ( .A(n8326), .B(n7635), .Z(n7637) );
  XOR U18883 ( .A(n8327), .B(n8328), .Z(n7635) );
  ANDN U18884 ( .B(n8329), .A(n8330), .Z(n8327) );
  AND U18885 ( .A(b[13]), .B(a[103]), .Z(n8326) );
  XNOR U18886 ( .A(n8331), .B(n7640), .Z(n7642) );
  XOR U18887 ( .A(n8332), .B(n8333), .Z(n7640) );
  ANDN U18888 ( .B(n8334), .A(n8335), .Z(n8332) );
  AND U18889 ( .A(b[12]), .B(a[104]), .Z(n8331) );
  XNOR U18890 ( .A(n8336), .B(n7645), .Z(n7647) );
  XOR U18891 ( .A(n8337), .B(n8338), .Z(n7645) );
  ANDN U18892 ( .B(n8339), .A(n8340), .Z(n8337) );
  AND U18893 ( .A(b[11]), .B(a[105]), .Z(n8336) );
  XNOR U18894 ( .A(n8341), .B(n7650), .Z(n7652) );
  XOR U18895 ( .A(n8342), .B(n8343), .Z(n7650) );
  ANDN U18896 ( .B(n8344), .A(n8345), .Z(n8342) );
  AND U18897 ( .A(b[10]), .B(a[106]), .Z(n8341) );
  XNOR U18898 ( .A(n8346), .B(n7655), .Z(n7657) );
  XOR U18899 ( .A(n8347), .B(n8348), .Z(n7655) );
  ANDN U18900 ( .B(n8349), .A(n8350), .Z(n8347) );
  AND U18901 ( .A(b[9]), .B(a[107]), .Z(n8346) );
  XNOR U18902 ( .A(n8351), .B(n7660), .Z(n7662) );
  XOR U18903 ( .A(n8352), .B(n8353), .Z(n7660) );
  ANDN U18904 ( .B(n8354), .A(n8355), .Z(n8352) );
  AND U18905 ( .A(b[8]), .B(a[108]), .Z(n8351) );
  XNOR U18906 ( .A(n8356), .B(n7665), .Z(n7667) );
  XOR U18907 ( .A(n8357), .B(n8358), .Z(n7665) );
  ANDN U18908 ( .B(n8359), .A(n8360), .Z(n8357) );
  AND U18909 ( .A(b[7]), .B(a[109]), .Z(n8356) );
  XNOR U18910 ( .A(n8361), .B(n7670), .Z(n7672) );
  XOR U18911 ( .A(n8362), .B(n8363), .Z(n7670) );
  ANDN U18912 ( .B(n8364), .A(n8365), .Z(n8362) );
  AND U18913 ( .A(b[6]), .B(a[110]), .Z(n8361) );
  XNOR U18914 ( .A(n8366), .B(n7675), .Z(n7677) );
  XOR U18915 ( .A(n8367), .B(n8368), .Z(n7675) );
  ANDN U18916 ( .B(n8369), .A(n8370), .Z(n8367) );
  AND U18917 ( .A(b[5]), .B(a[111]), .Z(n8366) );
  XNOR U18918 ( .A(n8371), .B(n7680), .Z(n7682) );
  XOR U18919 ( .A(n8372), .B(n8373), .Z(n7680) );
  ANDN U18920 ( .B(n8374), .A(n8375), .Z(n8372) );
  AND U18921 ( .A(b[4]), .B(a[112]), .Z(n8371) );
  XNOR U18922 ( .A(n8376), .B(n8377), .Z(n7694) );
  NANDN U18923 ( .A(n8378), .B(n8379), .Z(n8377) );
  XNOR U18924 ( .A(n8380), .B(n7685), .Z(n7687) );
  XNOR U18925 ( .A(n8381), .B(n8382), .Z(n7685) );
  AND U18926 ( .A(n8383), .B(n8384), .Z(n8381) );
  AND U18927 ( .A(b[3]), .B(a[113]), .Z(n8380) );
  NAND U18928 ( .A(a[116]), .B(b[0]), .Z(n7006) );
  XNOR U18929 ( .A(n7700), .B(n7701), .Z(c[115]) );
  XNOR U18930 ( .A(n8378), .B(n8379), .Z(n7701) );
  XOR U18931 ( .A(n8376), .B(n8385), .Z(n8379) );
  NAND U18932 ( .A(b[1]), .B(a[114]), .Z(n8385) );
  XOR U18933 ( .A(n8384), .B(n8386), .Z(n8378) );
  XOR U18934 ( .A(n8376), .B(n8383), .Z(n8386) );
  XNOR U18935 ( .A(n8387), .B(n8382), .Z(n8383) );
  AND U18936 ( .A(b[2]), .B(a[113]), .Z(n8387) );
  NANDN U18937 ( .A(n8388), .B(n8389), .Z(n8376) );
  XOR U18938 ( .A(n8382), .B(n8374), .Z(n8390) );
  XNOR U18939 ( .A(n8373), .B(n8369), .Z(n8391) );
  XNOR U18940 ( .A(n8368), .B(n8364), .Z(n8392) );
  XNOR U18941 ( .A(n8363), .B(n8359), .Z(n8393) );
  XNOR U18942 ( .A(n8358), .B(n8354), .Z(n8394) );
  XNOR U18943 ( .A(n8353), .B(n8349), .Z(n8395) );
  XNOR U18944 ( .A(n8348), .B(n8344), .Z(n8396) );
  XNOR U18945 ( .A(n8343), .B(n8339), .Z(n8397) );
  XNOR U18946 ( .A(n8338), .B(n8334), .Z(n8398) );
  XNOR U18947 ( .A(n8333), .B(n8329), .Z(n8399) );
  XNOR U18948 ( .A(n8328), .B(n8324), .Z(n8400) );
  XNOR U18949 ( .A(n8323), .B(n8319), .Z(n8401) );
  XNOR U18950 ( .A(n8318), .B(n8314), .Z(n8402) );
  XNOR U18951 ( .A(n8313), .B(n8309), .Z(n8403) );
  XNOR U18952 ( .A(n8308), .B(n8304), .Z(n8404) );
  XNOR U18953 ( .A(n8303), .B(n8299), .Z(n8405) );
  XNOR U18954 ( .A(n8298), .B(n8294), .Z(n8406) );
  XNOR U18955 ( .A(n8293), .B(n8289), .Z(n8407) );
  XNOR U18956 ( .A(n8288), .B(n8284), .Z(n8408) );
  XNOR U18957 ( .A(n8283), .B(n8279), .Z(n8409) );
  XNOR U18958 ( .A(n8278), .B(n8274), .Z(n8410) );
  XNOR U18959 ( .A(n8273), .B(n8269), .Z(n8411) );
  XNOR U18960 ( .A(n8268), .B(n8264), .Z(n8412) );
  XNOR U18961 ( .A(n8263), .B(n8259), .Z(n8413) );
  XNOR U18962 ( .A(n8258), .B(n8254), .Z(n8414) );
  XNOR U18963 ( .A(n8253), .B(n8249), .Z(n8415) );
  XNOR U18964 ( .A(n8248), .B(n8244), .Z(n8416) );
  XNOR U18965 ( .A(n8243), .B(n8239), .Z(n8417) );
  XNOR U18966 ( .A(n8238), .B(n8234), .Z(n8418) );
  XNOR U18967 ( .A(n8233), .B(n8229), .Z(n8419) );
  XNOR U18968 ( .A(n8228), .B(n8224), .Z(n8420) );
  XNOR U18969 ( .A(n8223), .B(n8219), .Z(n8421) );
  XNOR U18970 ( .A(n8218), .B(n8214), .Z(n8422) );
  XNOR U18971 ( .A(n8213), .B(n8209), .Z(n8423) );
  XNOR U18972 ( .A(n8208), .B(n8204), .Z(n8424) );
  XNOR U18973 ( .A(n8203), .B(n8199), .Z(n8425) );
  XNOR U18974 ( .A(n8198), .B(n8194), .Z(n8426) );
  XNOR U18975 ( .A(n8193), .B(n8189), .Z(n8427) );
  XNOR U18976 ( .A(n8188), .B(n8184), .Z(n8428) );
  XNOR U18977 ( .A(n8183), .B(n8179), .Z(n8429) );
  XNOR U18978 ( .A(n8178), .B(n8174), .Z(n8430) );
  XNOR U18979 ( .A(n8173), .B(n8169), .Z(n8431) );
  XNOR U18980 ( .A(n8168), .B(n8164), .Z(n8432) );
  XNOR U18981 ( .A(n8163), .B(n8159), .Z(n8433) );
  XNOR U18982 ( .A(n8158), .B(n8154), .Z(n8434) );
  XNOR U18983 ( .A(n8153), .B(n8149), .Z(n8435) );
  XNOR U18984 ( .A(n8148), .B(n8144), .Z(n8436) );
  XNOR U18985 ( .A(n8143), .B(n8139), .Z(n8437) );
  XNOR U18986 ( .A(n8138), .B(n8134), .Z(n8438) );
  XNOR U18987 ( .A(n8133), .B(n8129), .Z(n8439) );
  XNOR U18988 ( .A(n8128), .B(n8124), .Z(n8440) );
  XNOR U18989 ( .A(n8123), .B(n8119), .Z(n8441) );
  XNOR U18990 ( .A(n8118), .B(n8114), .Z(n8442) );
  XNOR U18991 ( .A(n8113), .B(n8109), .Z(n8443) );
  XNOR U18992 ( .A(n8108), .B(n8104), .Z(n8444) );
  XNOR U18993 ( .A(n8103), .B(n8099), .Z(n8445) );
  XNOR U18994 ( .A(n8098), .B(n8094), .Z(n8446) );
  XNOR U18995 ( .A(n8093), .B(n8089), .Z(n8447) );
  XNOR U18996 ( .A(n8088), .B(n8084), .Z(n8448) );
  XNOR U18997 ( .A(n8083), .B(n8079), .Z(n8449) );
  XNOR U18998 ( .A(n8078), .B(n8074), .Z(n8450) );
  XNOR U18999 ( .A(n8073), .B(n8069), .Z(n8451) );
  XNOR U19000 ( .A(n8068), .B(n8064), .Z(n8452) );
  XNOR U19001 ( .A(n8063), .B(n8059), .Z(n8453) );
  XNOR U19002 ( .A(n8058), .B(n8054), .Z(n8454) );
  XNOR U19003 ( .A(n8053), .B(n8049), .Z(n8455) );
  XNOR U19004 ( .A(n8048), .B(n8044), .Z(n8456) );
  XNOR U19005 ( .A(n8043), .B(n8039), .Z(n8457) );
  XNOR U19006 ( .A(n8038), .B(n8034), .Z(n8458) );
  XNOR U19007 ( .A(n8033), .B(n8029), .Z(n8459) );
  XNOR U19008 ( .A(n8028), .B(n8024), .Z(n8460) );
  XNOR U19009 ( .A(n8023), .B(n8019), .Z(n8461) );
  XNOR U19010 ( .A(n8018), .B(n8014), .Z(n8462) );
  XNOR U19011 ( .A(n8013), .B(n8009), .Z(n8463) );
  XNOR U19012 ( .A(n8008), .B(n8004), .Z(n8464) );
  XNOR U19013 ( .A(n8003), .B(n7999), .Z(n8465) );
  XNOR U19014 ( .A(n7998), .B(n7994), .Z(n8466) );
  XNOR U19015 ( .A(n7993), .B(n7989), .Z(n8467) );
  XNOR U19016 ( .A(n7988), .B(n7984), .Z(n8468) );
  XNOR U19017 ( .A(n7983), .B(n7979), .Z(n8469) );
  XNOR U19018 ( .A(n7978), .B(n7974), .Z(n8470) );
  XNOR U19019 ( .A(n7973), .B(n7969), .Z(n8471) );
  XNOR U19020 ( .A(n7968), .B(n7964), .Z(n8472) );
  XNOR U19021 ( .A(n7963), .B(n7959), .Z(n8473) );
  XNOR U19022 ( .A(n7958), .B(n7954), .Z(n8474) );
  XNOR U19023 ( .A(n7953), .B(n7949), .Z(n8475) );
  XNOR U19024 ( .A(n7948), .B(n7944), .Z(n8476) );
  XNOR U19025 ( .A(n7943), .B(n7939), .Z(n8477) );
  XNOR U19026 ( .A(n7938), .B(n7934), .Z(n8478) );
  XNOR U19027 ( .A(n7933), .B(n7929), .Z(n8479) );
  XNOR U19028 ( .A(n7928), .B(n7924), .Z(n8480) );
  XNOR U19029 ( .A(n7923), .B(n7919), .Z(n8481) );
  XNOR U19030 ( .A(n7918), .B(n7914), .Z(n8482) );
  XNOR U19031 ( .A(n7913), .B(n7909), .Z(n8483) );
  XNOR U19032 ( .A(n7908), .B(n7904), .Z(n8484) );
  XNOR U19033 ( .A(n7903), .B(n7899), .Z(n8485) );
  XNOR U19034 ( .A(n7898), .B(n7894), .Z(n8486) );
  XNOR U19035 ( .A(n7893), .B(n7889), .Z(n8487) );
  XNOR U19036 ( .A(n7888), .B(n7884), .Z(n8488) );
  XNOR U19037 ( .A(n7883), .B(n7879), .Z(n8489) );
  XNOR U19038 ( .A(n7878), .B(n7874), .Z(n8490) );
  XNOR U19039 ( .A(n7873), .B(n7869), .Z(n8491) );
  XNOR U19040 ( .A(n7868), .B(n7864), .Z(n8492) );
  XNOR U19041 ( .A(n7863), .B(n7859), .Z(n8493) );
  XNOR U19042 ( .A(n7858), .B(n7854), .Z(n8494) );
  XNOR U19043 ( .A(n7853), .B(n7849), .Z(n8495) );
  XNOR U19044 ( .A(n7848), .B(n7844), .Z(n8496) );
  XNOR U19045 ( .A(n7843), .B(n7839), .Z(n8497) );
  XNOR U19046 ( .A(n7838), .B(n7834), .Z(n8498) );
  XNOR U19047 ( .A(n7833), .B(n7829), .Z(n8499) );
  XNOR U19048 ( .A(n7828), .B(n7824), .Z(n8500) );
  XNOR U19049 ( .A(n7823), .B(n7819), .Z(n8501) );
  XNOR U19050 ( .A(n8502), .B(n7818), .Z(n7819) );
  AND U19051 ( .A(a[0]), .B(b[115]), .Z(n8502) );
  XOR U19052 ( .A(n8503), .B(n7818), .Z(n7820) );
  XNOR U19053 ( .A(n8504), .B(n8505), .Z(n7818) );
  ANDN U19054 ( .B(n8506), .A(n8507), .Z(n8504) );
  AND U19055 ( .A(a[1]), .B(b[114]), .Z(n8503) );
  XNOR U19056 ( .A(n8508), .B(n7823), .Z(n7825) );
  XOR U19057 ( .A(n8509), .B(n8510), .Z(n7823) );
  ANDN U19058 ( .B(n8511), .A(n8512), .Z(n8509) );
  AND U19059 ( .A(a[2]), .B(b[113]), .Z(n8508) );
  XNOR U19060 ( .A(n8513), .B(n7828), .Z(n7830) );
  XOR U19061 ( .A(n8514), .B(n8515), .Z(n7828) );
  ANDN U19062 ( .B(n8516), .A(n8517), .Z(n8514) );
  AND U19063 ( .A(a[3]), .B(b[112]), .Z(n8513) );
  XNOR U19064 ( .A(n8518), .B(n7833), .Z(n7835) );
  XOR U19065 ( .A(n8519), .B(n8520), .Z(n7833) );
  ANDN U19066 ( .B(n8521), .A(n8522), .Z(n8519) );
  AND U19067 ( .A(a[4]), .B(b[111]), .Z(n8518) );
  XNOR U19068 ( .A(n8523), .B(n7838), .Z(n7840) );
  XOR U19069 ( .A(n8524), .B(n8525), .Z(n7838) );
  ANDN U19070 ( .B(n8526), .A(n8527), .Z(n8524) );
  AND U19071 ( .A(a[5]), .B(b[110]), .Z(n8523) );
  XNOR U19072 ( .A(n8528), .B(n7843), .Z(n7845) );
  XOR U19073 ( .A(n8529), .B(n8530), .Z(n7843) );
  ANDN U19074 ( .B(n8531), .A(n8532), .Z(n8529) );
  AND U19075 ( .A(a[6]), .B(b[109]), .Z(n8528) );
  XNOR U19076 ( .A(n8533), .B(n7848), .Z(n7850) );
  XOR U19077 ( .A(n8534), .B(n8535), .Z(n7848) );
  ANDN U19078 ( .B(n8536), .A(n8537), .Z(n8534) );
  AND U19079 ( .A(a[7]), .B(b[108]), .Z(n8533) );
  XNOR U19080 ( .A(n8538), .B(n7853), .Z(n7855) );
  XOR U19081 ( .A(n8539), .B(n8540), .Z(n7853) );
  ANDN U19082 ( .B(n8541), .A(n8542), .Z(n8539) );
  AND U19083 ( .A(a[8]), .B(b[107]), .Z(n8538) );
  XNOR U19084 ( .A(n8543), .B(n7858), .Z(n7860) );
  XOR U19085 ( .A(n8544), .B(n8545), .Z(n7858) );
  ANDN U19086 ( .B(n8546), .A(n8547), .Z(n8544) );
  AND U19087 ( .A(a[9]), .B(b[106]), .Z(n8543) );
  XNOR U19088 ( .A(n8548), .B(n7863), .Z(n7865) );
  XOR U19089 ( .A(n8549), .B(n8550), .Z(n7863) );
  ANDN U19090 ( .B(n8551), .A(n8552), .Z(n8549) );
  AND U19091 ( .A(a[10]), .B(b[105]), .Z(n8548) );
  XNOR U19092 ( .A(n8553), .B(n7868), .Z(n7870) );
  XOR U19093 ( .A(n8554), .B(n8555), .Z(n7868) );
  ANDN U19094 ( .B(n8556), .A(n8557), .Z(n8554) );
  AND U19095 ( .A(a[11]), .B(b[104]), .Z(n8553) );
  XNOR U19096 ( .A(n8558), .B(n7873), .Z(n7875) );
  XOR U19097 ( .A(n8559), .B(n8560), .Z(n7873) );
  ANDN U19098 ( .B(n8561), .A(n8562), .Z(n8559) );
  AND U19099 ( .A(a[12]), .B(b[103]), .Z(n8558) );
  XNOR U19100 ( .A(n8563), .B(n7878), .Z(n7880) );
  XOR U19101 ( .A(n8564), .B(n8565), .Z(n7878) );
  ANDN U19102 ( .B(n8566), .A(n8567), .Z(n8564) );
  AND U19103 ( .A(a[13]), .B(b[102]), .Z(n8563) );
  XNOR U19104 ( .A(n8568), .B(n7883), .Z(n7885) );
  XOR U19105 ( .A(n8569), .B(n8570), .Z(n7883) );
  ANDN U19106 ( .B(n8571), .A(n8572), .Z(n8569) );
  AND U19107 ( .A(a[14]), .B(b[101]), .Z(n8568) );
  XNOR U19108 ( .A(n8573), .B(n7888), .Z(n7890) );
  XOR U19109 ( .A(n8574), .B(n8575), .Z(n7888) );
  ANDN U19110 ( .B(n8576), .A(n8577), .Z(n8574) );
  AND U19111 ( .A(a[15]), .B(b[100]), .Z(n8573) );
  XNOR U19112 ( .A(n8578), .B(n7893), .Z(n7895) );
  XOR U19113 ( .A(n8579), .B(n8580), .Z(n7893) );
  ANDN U19114 ( .B(n8581), .A(n8582), .Z(n8579) );
  AND U19115 ( .A(a[16]), .B(b[99]), .Z(n8578) );
  XNOR U19116 ( .A(n8583), .B(n7898), .Z(n7900) );
  XOR U19117 ( .A(n8584), .B(n8585), .Z(n7898) );
  ANDN U19118 ( .B(n8586), .A(n8587), .Z(n8584) );
  AND U19119 ( .A(a[17]), .B(b[98]), .Z(n8583) );
  XNOR U19120 ( .A(n8588), .B(n7903), .Z(n7905) );
  XOR U19121 ( .A(n8589), .B(n8590), .Z(n7903) );
  ANDN U19122 ( .B(n8591), .A(n8592), .Z(n8589) );
  AND U19123 ( .A(a[18]), .B(b[97]), .Z(n8588) );
  XNOR U19124 ( .A(n8593), .B(n7908), .Z(n7910) );
  XOR U19125 ( .A(n8594), .B(n8595), .Z(n7908) );
  ANDN U19126 ( .B(n8596), .A(n8597), .Z(n8594) );
  AND U19127 ( .A(a[19]), .B(b[96]), .Z(n8593) );
  XNOR U19128 ( .A(n8598), .B(n7913), .Z(n7915) );
  XOR U19129 ( .A(n8599), .B(n8600), .Z(n7913) );
  ANDN U19130 ( .B(n8601), .A(n8602), .Z(n8599) );
  AND U19131 ( .A(a[20]), .B(b[95]), .Z(n8598) );
  XNOR U19132 ( .A(n8603), .B(n7918), .Z(n7920) );
  XOR U19133 ( .A(n8604), .B(n8605), .Z(n7918) );
  ANDN U19134 ( .B(n8606), .A(n8607), .Z(n8604) );
  AND U19135 ( .A(a[21]), .B(b[94]), .Z(n8603) );
  XNOR U19136 ( .A(n8608), .B(n7923), .Z(n7925) );
  XOR U19137 ( .A(n8609), .B(n8610), .Z(n7923) );
  ANDN U19138 ( .B(n8611), .A(n8612), .Z(n8609) );
  AND U19139 ( .A(a[22]), .B(b[93]), .Z(n8608) );
  XNOR U19140 ( .A(n8613), .B(n7928), .Z(n7930) );
  XOR U19141 ( .A(n8614), .B(n8615), .Z(n7928) );
  ANDN U19142 ( .B(n8616), .A(n8617), .Z(n8614) );
  AND U19143 ( .A(a[23]), .B(b[92]), .Z(n8613) );
  XNOR U19144 ( .A(n8618), .B(n7933), .Z(n7935) );
  XOR U19145 ( .A(n8619), .B(n8620), .Z(n7933) );
  ANDN U19146 ( .B(n8621), .A(n8622), .Z(n8619) );
  AND U19147 ( .A(a[24]), .B(b[91]), .Z(n8618) );
  XNOR U19148 ( .A(n8623), .B(n7938), .Z(n7940) );
  XOR U19149 ( .A(n8624), .B(n8625), .Z(n7938) );
  ANDN U19150 ( .B(n8626), .A(n8627), .Z(n8624) );
  AND U19151 ( .A(a[25]), .B(b[90]), .Z(n8623) );
  XNOR U19152 ( .A(n8628), .B(n7943), .Z(n7945) );
  XOR U19153 ( .A(n8629), .B(n8630), .Z(n7943) );
  ANDN U19154 ( .B(n8631), .A(n8632), .Z(n8629) );
  AND U19155 ( .A(a[26]), .B(b[89]), .Z(n8628) );
  XNOR U19156 ( .A(n8633), .B(n7948), .Z(n7950) );
  XOR U19157 ( .A(n8634), .B(n8635), .Z(n7948) );
  ANDN U19158 ( .B(n8636), .A(n8637), .Z(n8634) );
  AND U19159 ( .A(a[27]), .B(b[88]), .Z(n8633) );
  XNOR U19160 ( .A(n8638), .B(n7953), .Z(n7955) );
  XOR U19161 ( .A(n8639), .B(n8640), .Z(n7953) );
  ANDN U19162 ( .B(n8641), .A(n8642), .Z(n8639) );
  AND U19163 ( .A(a[28]), .B(b[87]), .Z(n8638) );
  XNOR U19164 ( .A(n8643), .B(n7958), .Z(n7960) );
  XOR U19165 ( .A(n8644), .B(n8645), .Z(n7958) );
  ANDN U19166 ( .B(n8646), .A(n8647), .Z(n8644) );
  AND U19167 ( .A(a[29]), .B(b[86]), .Z(n8643) );
  XNOR U19168 ( .A(n8648), .B(n7963), .Z(n7965) );
  XOR U19169 ( .A(n8649), .B(n8650), .Z(n7963) );
  ANDN U19170 ( .B(n8651), .A(n8652), .Z(n8649) );
  AND U19171 ( .A(a[30]), .B(b[85]), .Z(n8648) );
  XNOR U19172 ( .A(n8653), .B(n7968), .Z(n7970) );
  XOR U19173 ( .A(n8654), .B(n8655), .Z(n7968) );
  ANDN U19174 ( .B(n8656), .A(n8657), .Z(n8654) );
  AND U19175 ( .A(a[31]), .B(b[84]), .Z(n8653) );
  XNOR U19176 ( .A(n8658), .B(n7973), .Z(n7975) );
  XOR U19177 ( .A(n8659), .B(n8660), .Z(n7973) );
  ANDN U19178 ( .B(n8661), .A(n8662), .Z(n8659) );
  AND U19179 ( .A(a[32]), .B(b[83]), .Z(n8658) );
  XNOR U19180 ( .A(n8663), .B(n7978), .Z(n7980) );
  XOR U19181 ( .A(n8664), .B(n8665), .Z(n7978) );
  ANDN U19182 ( .B(n8666), .A(n8667), .Z(n8664) );
  AND U19183 ( .A(a[33]), .B(b[82]), .Z(n8663) );
  XNOR U19184 ( .A(n8668), .B(n7983), .Z(n7985) );
  XOR U19185 ( .A(n8669), .B(n8670), .Z(n7983) );
  ANDN U19186 ( .B(n8671), .A(n8672), .Z(n8669) );
  AND U19187 ( .A(a[34]), .B(b[81]), .Z(n8668) );
  XNOR U19188 ( .A(n8673), .B(n7988), .Z(n7990) );
  XOR U19189 ( .A(n8674), .B(n8675), .Z(n7988) );
  ANDN U19190 ( .B(n8676), .A(n8677), .Z(n8674) );
  AND U19191 ( .A(a[35]), .B(b[80]), .Z(n8673) );
  XNOR U19192 ( .A(n8678), .B(n7993), .Z(n7995) );
  XOR U19193 ( .A(n8679), .B(n8680), .Z(n7993) );
  ANDN U19194 ( .B(n8681), .A(n8682), .Z(n8679) );
  AND U19195 ( .A(a[36]), .B(b[79]), .Z(n8678) );
  XNOR U19196 ( .A(n8683), .B(n7998), .Z(n8000) );
  XOR U19197 ( .A(n8684), .B(n8685), .Z(n7998) );
  ANDN U19198 ( .B(n8686), .A(n8687), .Z(n8684) );
  AND U19199 ( .A(a[37]), .B(b[78]), .Z(n8683) );
  XNOR U19200 ( .A(n8688), .B(n8003), .Z(n8005) );
  XOR U19201 ( .A(n8689), .B(n8690), .Z(n8003) );
  ANDN U19202 ( .B(n8691), .A(n8692), .Z(n8689) );
  AND U19203 ( .A(a[38]), .B(b[77]), .Z(n8688) );
  XNOR U19204 ( .A(n8693), .B(n8008), .Z(n8010) );
  XOR U19205 ( .A(n8694), .B(n8695), .Z(n8008) );
  ANDN U19206 ( .B(n8696), .A(n8697), .Z(n8694) );
  AND U19207 ( .A(a[39]), .B(b[76]), .Z(n8693) );
  XNOR U19208 ( .A(n8698), .B(n8013), .Z(n8015) );
  XOR U19209 ( .A(n8699), .B(n8700), .Z(n8013) );
  ANDN U19210 ( .B(n8701), .A(n8702), .Z(n8699) );
  AND U19211 ( .A(a[40]), .B(b[75]), .Z(n8698) );
  XNOR U19212 ( .A(n8703), .B(n8018), .Z(n8020) );
  XOR U19213 ( .A(n8704), .B(n8705), .Z(n8018) );
  ANDN U19214 ( .B(n8706), .A(n8707), .Z(n8704) );
  AND U19215 ( .A(a[41]), .B(b[74]), .Z(n8703) );
  XNOR U19216 ( .A(n8708), .B(n8023), .Z(n8025) );
  XOR U19217 ( .A(n8709), .B(n8710), .Z(n8023) );
  ANDN U19218 ( .B(n8711), .A(n8712), .Z(n8709) );
  AND U19219 ( .A(a[42]), .B(b[73]), .Z(n8708) );
  XNOR U19220 ( .A(n8713), .B(n8028), .Z(n8030) );
  XOR U19221 ( .A(n8714), .B(n8715), .Z(n8028) );
  ANDN U19222 ( .B(n8716), .A(n8717), .Z(n8714) );
  AND U19223 ( .A(a[43]), .B(b[72]), .Z(n8713) );
  XNOR U19224 ( .A(n8718), .B(n8033), .Z(n8035) );
  XOR U19225 ( .A(n8719), .B(n8720), .Z(n8033) );
  ANDN U19226 ( .B(n8721), .A(n8722), .Z(n8719) );
  AND U19227 ( .A(a[44]), .B(b[71]), .Z(n8718) );
  XNOR U19228 ( .A(n8723), .B(n8038), .Z(n8040) );
  XOR U19229 ( .A(n8724), .B(n8725), .Z(n8038) );
  ANDN U19230 ( .B(n8726), .A(n8727), .Z(n8724) );
  AND U19231 ( .A(a[45]), .B(b[70]), .Z(n8723) );
  XNOR U19232 ( .A(n8728), .B(n8043), .Z(n8045) );
  XOR U19233 ( .A(n8729), .B(n8730), .Z(n8043) );
  ANDN U19234 ( .B(n8731), .A(n8732), .Z(n8729) );
  AND U19235 ( .A(a[46]), .B(b[69]), .Z(n8728) );
  XNOR U19236 ( .A(n8733), .B(n8048), .Z(n8050) );
  XOR U19237 ( .A(n8734), .B(n8735), .Z(n8048) );
  ANDN U19238 ( .B(n8736), .A(n8737), .Z(n8734) );
  AND U19239 ( .A(a[47]), .B(b[68]), .Z(n8733) );
  XNOR U19240 ( .A(n8738), .B(n8053), .Z(n8055) );
  XOR U19241 ( .A(n8739), .B(n8740), .Z(n8053) );
  ANDN U19242 ( .B(n8741), .A(n8742), .Z(n8739) );
  AND U19243 ( .A(a[48]), .B(b[67]), .Z(n8738) );
  XNOR U19244 ( .A(n8743), .B(n8058), .Z(n8060) );
  XOR U19245 ( .A(n8744), .B(n8745), .Z(n8058) );
  ANDN U19246 ( .B(n8746), .A(n8747), .Z(n8744) );
  AND U19247 ( .A(a[49]), .B(b[66]), .Z(n8743) );
  XNOR U19248 ( .A(n8748), .B(n8063), .Z(n8065) );
  XOR U19249 ( .A(n8749), .B(n8750), .Z(n8063) );
  ANDN U19250 ( .B(n8751), .A(n8752), .Z(n8749) );
  AND U19251 ( .A(a[50]), .B(b[65]), .Z(n8748) );
  XNOR U19252 ( .A(n8753), .B(n8068), .Z(n8070) );
  XOR U19253 ( .A(n8754), .B(n8755), .Z(n8068) );
  ANDN U19254 ( .B(n8756), .A(n8757), .Z(n8754) );
  AND U19255 ( .A(a[51]), .B(b[64]), .Z(n8753) );
  XNOR U19256 ( .A(n8758), .B(n8073), .Z(n8075) );
  XOR U19257 ( .A(n8759), .B(n8760), .Z(n8073) );
  ANDN U19258 ( .B(n8761), .A(n8762), .Z(n8759) );
  AND U19259 ( .A(a[52]), .B(b[63]), .Z(n8758) );
  XNOR U19260 ( .A(n8763), .B(n8078), .Z(n8080) );
  XOR U19261 ( .A(n8764), .B(n8765), .Z(n8078) );
  ANDN U19262 ( .B(n8766), .A(n8767), .Z(n8764) );
  AND U19263 ( .A(a[53]), .B(b[62]), .Z(n8763) );
  XNOR U19264 ( .A(n8768), .B(n8083), .Z(n8085) );
  XOR U19265 ( .A(n8769), .B(n8770), .Z(n8083) );
  ANDN U19266 ( .B(n8771), .A(n8772), .Z(n8769) );
  AND U19267 ( .A(a[54]), .B(b[61]), .Z(n8768) );
  XNOR U19268 ( .A(n8773), .B(n8088), .Z(n8090) );
  XOR U19269 ( .A(n8774), .B(n8775), .Z(n8088) );
  ANDN U19270 ( .B(n8776), .A(n8777), .Z(n8774) );
  AND U19271 ( .A(a[55]), .B(b[60]), .Z(n8773) );
  XNOR U19272 ( .A(n8778), .B(n8093), .Z(n8095) );
  XOR U19273 ( .A(n8779), .B(n8780), .Z(n8093) );
  ANDN U19274 ( .B(n8781), .A(n8782), .Z(n8779) );
  AND U19275 ( .A(a[56]), .B(b[59]), .Z(n8778) );
  XNOR U19276 ( .A(n8783), .B(n8098), .Z(n8100) );
  XOR U19277 ( .A(n8784), .B(n8785), .Z(n8098) );
  ANDN U19278 ( .B(n8786), .A(n8787), .Z(n8784) );
  AND U19279 ( .A(a[57]), .B(b[58]), .Z(n8783) );
  XNOR U19280 ( .A(n8788), .B(n8103), .Z(n8105) );
  XOR U19281 ( .A(n8789), .B(n8790), .Z(n8103) );
  ANDN U19282 ( .B(n8791), .A(n8792), .Z(n8789) );
  AND U19283 ( .A(a[58]), .B(b[57]), .Z(n8788) );
  XNOR U19284 ( .A(n8793), .B(n8108), .Z(n8110) );
  XOR U19285 ( .A(n8794), .B(n8795), .Z(n8108) );
  ANDN U19286 ( .B(n8796), .A(n8797), .Z(n8794) );
  AND U19287 ( .A(a[59]), .B(b[56]), .Z(n8793) );
  XNOR U19288 ( .A(n8798), .B(n8113), .Z(n8115) );
  XOR U19289 ( .A(n8799), .B(n8800), .Z(n8113) );
  ANDN U19290 ( .B(n8801), .A(n8802), .Z(n8799) );
  AND U19291 ( .A(a[60]), .B(b[55]), .Z(n8798) );
  XNOR U19292 ( .A(n8803), .B(n8118), .Z(n8120) );
  XOR U19293 ( .A(n8804), .B(n8805), .Z(n8118) );
  ANDN U19294 ( .B(n8806), .A(n8807), .Z(n8804) );
  AND U19295 ( .A(a[61]), .B(b[54]), .Z(n8803) );
  XNOR U19296 ( .A(n8808), .B(n8123), .Z(n8125) );
  XOR U19297 ( .A(n8809), .B(n8810), .Z(n8123) );
  ANDN U19298 ( .B(n8811), .A(n8812), .Z(n8809) );
  AND U19299 ( .A(a[62]), .B(b[53]), .Z(n8808) );
  XNOR U19300 ( .A(n8813), .B(n8128), .Z(n8130) );
  XOR U19301 ( .A(n8814), .B(n8815), .Z(n8128) );
  ANDN U19302 ( .B(n8816), .A(n8817), .Z(n8814) );
  AND U19303 ( .A(a[63]), .B(b[52]), .Z(n8813) );
  XNOR U19304 ( .A(n8818), .B(n8133), .Z(n8135) );
  XOR U19305 ( .A(n8819), .B(n8820), .Z(n8133) );
  ANDN U19306 ( .B(n8821), .A(n8822), .Z(n8819) );
  AND U19307 ( .A(a[64]), .B(b[51]), .Z(n8818) );
  XNOR U19308 ( .A(n8823), .B(n8138), .Z(n8140) );
  XOR U19309 ( .A(n8824), .B(n8825), .Z(n8138) );
  ANDN U19310 ( .B(n8826), .A(n8827), .Z(n8824) );
  AND U19311 ( .A(a[65]), .B(b[50]), .Z(n8823) );
  XNOR U19312 ( .A(n8828), .B(n8143), .Z(n8145) );
  XOR U19313 ( .A(n8829), .B(n8830), .Z(n8143) );
  ANDN U19314 ( .B(n8831), .A(n8832), .Z(n8829) );
  AND U19315 ( .A(a[66]), .B(b[49]), .Z(n8828) );
  XNOR U19316 ( .A(n8833), .B(n8148), .Z(n8150) );
  XOR U19317 ( .A(n8834), .B(n8835), .Z(n8148) );
  ANDN U19318 ( .B(n8836), .A(n8837), .Z(n8834) );
  AND U19319 ( .A(a[67]), .B(b[48]), .Z(n8833) );
  XNOR U19320 ( .A(n8838), .B(n8153), .Z(n8155) );
  XOR U19321 ( .A(n8839), .B(n8840), .Z(n8153) );
  ANDN U19322 ( .B(n8841), .A(n8842), .Z(n8839) );
  AND U19323 ( .A(a[68]), .B(b[47]), .Z(n8838) );
  XNOR U19324 ( .A(n8843), .B(n8158), .Z(n8160) );
  XOR U19325 ( .A(n8844), .B(n8845), .Z(n8158) );
  ANDN U19326 ( .B(n8846), .A(n8847), .Z(n8844) );
  AND U19327 ( .A(a[69]), .B(b[46]), .Z(n8843) );
  XNOR U19328 ( .A(n8848), .B(n8163), .Z(n8165) );
  XOR U19329 ( .A(n8849), .B(n8850), .Z(n8163) );
  ANDN U19330 ( .B(n8851), .A(n8852), .Z(n8849) );
  AND U19331 ( .A(a[70]), .B(b[45]), .Z(n8848) );
  XNOR U19332 ( .A(n8853), .B(n8168), .Z(n8170) );
  XOR U19333 ( .A(n8854), .B(n8855), .Z(n8168) );
  ANDN U19334 ( .B(n8856), .A(n8857), .Z(n8854) );
  AND U19335 ( .A(a[71]), .B(b[44]), .Z(n8853) );
  XNOR U19336 ( .A(n8858), .B(n8173), .Z(n8175) );
  XOR U19337 ( .A(n8859), .B(n8860), .Z(n8173) );
  ANDN U19338 ( .B(n8861), .A(n8862), .Z(n8859) );
  AND U19339 ( .A(a[72]), .B(b[43]), .Z(n8858) );
  XNOR U19340 ( .A(n8863), .B(n8178), .Z(n8180) );
  XOR U19341 ( .A(n8864), .B(n8865), .Z(n8178) );
  ANDN U19342 ( .B(n8866), .A(n8867), .Z(n8864) );
  AND U19343 ( .A(a[73]), .B(b[42]), .Z(n8863) );
  XNOR U19344 ( .A(n8868), .B(n8183), .Z(n8185) );
  XOR U19345 ( .A(n8869), .B(n8870), .Z(n8183) );
  ANDN U19346 ( .B(n8871), .A(n8872), .Z(n8869) );
  AND U19347 ( .A(a[74]), .B(b[41]), .Z(n8868) );
  XNOR U19348 ( .A(n8873), .B(n8188), .Z(n8190) );
  XOR U19349 ( .A(n8874), .B(n8875), .Z(n8188) );
  ANDN U19350 ( .B(n8876), .A(n8877), .Z(n8874) );
  AND U19351 ( .A(a[75]), .B(b[40]), .Z(n8873) );
  XNOR U19352 ( .A(n8878), .B(n8193), .Z(n8195) );
  XOR U19353 ( .A(n8879), .B(n8880), .Z(n8193) );
  ANDN U19354 ( .B(n8881), .A(n8882), .Z(n8879) );
  AND U19355 ( .A(a[76]), .B(b[39]), .Z(n8878) );
  XNOR U19356 ( .A(n8883), .B(n8198), .Z(n8200) );
  XOR U19357 ( .A(n8884), .B(n8885), .Z(n8198) );
  ANDN U19358 ( .B(n8886), .A(n8887), .Z(n8884) );
  AND U19359 ( .A(a[77]), .B(b[38]), .Z(n8883) );
  XNOR U19360 ( .A(n8888), .B(n8203), .Z(n8205) );
  XOR U19361 ( .A(n8889), .B(n8890), .Z(n8203) );
  ANDN U19362 ( .B(n8891), .A(n8892), .Z(n8889) );
  AND U19363 ( .A(a[78]), .B(b[37]), .Z(n8888) );
  XNOR U19364 ( .A(n8893), .B(n8208), .Z(n8210) );
  XOR U19365 ( .A(n8894), .B(n8895), .Z(n8208) );
  ANDN U19366 ( .B(n8896), .A(n8897), .Z(n8894) );
  AND U19367 ( .A(a[79]), .B(b[36]), .Z(n8893) );
  XNOR U19368 ( .A(n8898), .B(n8213), .Z(n8215) );
  XOR U19369 ( .A(n8899), .B(n8900), .Z(n8213) );
  ANDN U19370 ( .B(n8901), .A(n8902), .Z(n8899) );
  AND U19371 ( .A(a[80]), .B(b[35]), .Z(n8898) );
  XNOR U19372 ( .A(n8903), .B(n8218), .Z(n8220) );
  XOR U19373 ( .A(n8904), .B(n8905), .Z(n8218) );
  ANDN U19374 ( .B(n8906), .A(n8907), .Z(n8904) );
  AND U19375 ( .A(a[81]), .B(b[34]), .Z(n8903) );
  XNOR U19376 ( .A(n8908), .B(n8223), .Z(n8225) );
  XOR U19377 ( .A(n8909), .B(n8910), .Z(n8223) );
  ANDN U19378 ( .B(n8911), .A(n8912), .Z(n8909) );
  AND U19379 ( .A(a[82]), .B(b[33]), .Z(n8908) );
  XNOR U19380 ( .A(n8913), .B(n8228), .Z(n8230) );
  XOR U19381 ( .A(n8914), .B(n8915), .Z(n8228) );
  ANDN U19382 ( .B(n8916), .A(n8917), .Z(n8914) );
  AND U19383 ( .A(a[83]), .B(b[32]), .Z(n8913) );
  XNOR U19384 ( .A(n8918), .B(n8233), .Z(n8235) );
  XOR U19385 ( .A(n8919), .B(n8920), .Z(n8233) );
  ANDN U19386 ( .B(n8921), .A(n8922), .Z(n8919) );
  AND U19387 ( .A(a[84]), .B(b[31]), .Z(n8918) );
  XNOR U19388 ( .A(n8923), .B(n8238), .Z(n8240) );
  XOR U19389 ( .A(n8924), .B(n8925), .Z(n8238) );
  ANDN U19390 ( .B(n8926), .A(n8927), .Z(n8924) );
  AND U19391 ( .A(a[85]), .B(b[30]), .Z(n8923) );
  XNOR U19392 ( .A(n8928), .B(n8243), .Z(n8245) );
  XOR U19393 ( .A(n8929), .B(n8930), .Z(n8243) );
  ANDN U19394 ( .B(n8931), .A(n8932), .Z(n8929) );
  AND U19395 ( .A(a[86]), .B(b[29]), .Z(n8928) );
  XNOR U19396 ( .A(n8933), .B(n8248), .Z(n8250) );
  XOR U19397 ( .A(n8934), .B(n8935), .Z(n8248) );
  ANDN U19398 ( .B(n8936), .A(n8937), .Z(n8934) );
  AND U19399 ( .A(a[87]), .B(b[28]), .Z(n8933) );
  XNOR U19400 ( .A(n8938), .B(n8253), .Z(n8255) );
  XOR U19401 ( .A(n8939), .B(n8940), .Z(n8253) );
  ANDN U19402 ( .B(n8941), .A(n8942), .Z(n8939) );
  AND U19403 ( .A(a[88]), .B(b[27]), .Z(n8938) );
  XNOR U19404 ( .A(n8943), .B(n8258), .Z(n8260) );
  XOR U19405 ( .A(n8944), .B(n8945), .Z(n8258) );
  ANDN U19406 ( .B(n8946), .A(n8947), .Z(n8944) );
  AND U19407 ( .A(a[89]), .B(b[26]), .Z(n8943) );
  XNOR U19408 ( .A(n8948), .B(n8263), .Z(n8265) );
  XOR U19409 ( .A(n8949), .B(n8950), .Z(n8263) );
  ANDN U19410 ( .B(n8951), .A(n8952), .Z(n8949) );
  AND U19411 ( .A(a[90]), .B(b[25]), .Z(n8948) );
  XNOR U19412 ( .A(n8953), .B(n8268), .Z(n8270) );
  XOR U19413 ( .A(n8954), .B(n8955), .Z(n8268) );
  ANDN U19414 ( .B(n8956), .A(n8957), .Z(n8954) );
  AND U19415 ( .A(a[91]), .B(b[24]), .Z(n8953) );
  XNOR U19416 ( .A(n8958), .B(n8273), .Z(n8275) );
  XOR U19417 ( .A(n8959), .B(n8960), .Z(n8273) );
  ANDN U19418 ( .B(n8961), .A(n8962), .Z(n8959) );
  AND U19419 ( .A(a[92]), .B(b[23]), .Z(n8958) );
  XNOR U19420 ( .A(n8963), .B(n8278), .Z(n8280) );
  XOR U19421 ( .A(n8964), .B(n8965), .Z(n8278) );
  ANDN U19422 ( .B(n8966), .A(n8967), .Z(n8964) );
  AND U19423 ( .A(a[93]), .B(b[22]), .Z(n8963) );
  XNOR U19424 ( .A(n8968), .B(n8283), .Z(n8285) );
  XOR U19425 ( .A(n8969), .B(n8970), .Z(n8283) );
  ANDN U19426 ( .B(n8971), .A(n8972), .Z(n8969) );
  AND U19427 ( .A(a[94]), .B(b[21]), .Z(n8968) );
  XNOR U19428 ( .A(n8973), .B(n8288), .Z(n8290) );
  XOR U19429 ( .A(n8974), .B(n8975), .Z(n8288) );
  ANDN U19430 ( .B(n8976), .A(n8977), .Z(n8974) );
  AND U19431 ( .A(a[95]), .B(b[20]), .Z(n8973) );
  XNOR U19432 ( .A(n8978), .B(n8293), .Z(n8295) );
  XOR U19433 ( .A(n8979), .B(n8980), .Z(n8293) );
  ANDN U19434 ( .B(n8981), .A(n8982), .Z(n8979) );
  AND U19435 ( .A(a[96]), .B(b[19]), .Z(n8978) );
  XNOR U19436 ( .A(n8983), .B(n8298), .Z(n8300) );
  XOR U19437 ( .A(n8984), .B(n8985), .Z(n8298) );
  ANDN U19438 ( .B(n8986), .A(n8987), .Z(n8984) );
  AND U19439 ( .A(a[97]), .B(b[18]), .Z(n8983) );
  XNOR U19440 ( .A(n8988), .B(n8303), .Z(n8305) );
  XOR U19441 ( .A(n8989), .B(n8990), .Z(n8303) );
  ANDN U19442 ( .B(n8991), .A(n8992), .Z(n8989) );
  AND U19443 ( .A(a[98]), .B(b[17]), .Z(n8988) );
  XNOR U19444 ( .A(n8993), .B(n8308), .Z(n8310) );
  XOR U19445 ( .A(n8994), .B(n8995), .Z(n8308) );
  ANDN U19446 ( .B(n8996), .A(n8997), .Z(n8994) );
  AND U19447 ( .A(a[99]), .B(b[16]), .Z(n8993) );
  XNOR U19448 ( .A(n8998), .B(n8313), .Z(n8315) );
  XOR U19449 ( .A(n8999), .B(n9000), .Z(n8313) );
  ANDN U19450 ( .B(n9001), .A(n9002), .Z(n8999) );
  AND U19451 ( .A(b[15]), .B(a[100]), .Z(n8998) );
  XNOR U19452 ( .A(n9003), .B(n8318), .Z(n8320) );
  XOR U19453 ( .A(n9004), .B(n9005), .Z(n8318) );
  ANDN U19454 ( .B(n9006), .A(n9007), .Z(n9004) );
  AND U19455 ( .A(b[14]), .B(a[101]), .Z(n9003) );
  XNOR U19456 ( .A(n9008), .B(n8323), .Z(n8325) );
  XOR U19457 ( .A(n9009), .B(n9010), .Z(n8323) );
  ANDN U19458 ( .B(n9011), .A(n9012), .Z(n9009) );
  AND U19459 ( .A(b[13]), .B(a[102]), .Z(n9008) );
  XNOR U19460 ( .A(n9013), .B(n8328), .Z(n8330) );
  XOR U19461 ( .A(n9014), .B(n9015), .Z(n8328) );
  ANDN U19462 ( .B(n9016), .A(n9017), .Z(n9014) );
  AND U19463 ( .A(b[12]), .B(a[103]), .Z(n9013) );
  XNOR U19464 ( .A(n9018), .B(n8333), .Z(n8335) );
  XOR U19465 ( .A(n9019), .B(n9020), .Z(n8333) );
  ANDN U19466 ( .B(n9021), .A(n9022), .Z(n9019) );
  AND U19467 ( .A(b[11]), .B(a[104]), .Z(n9018) );
  XNOR U19468 ( .A(n9023), .B(n8338), .Z(n8340) );
  XOR U19469 ( .A(n9024), .B(n9025), .Z(n8338) );
  ANDN U19470 ( .B(n9026), .A(n9027), .Z(n9024) );
  AND U19471 ( .A(b[10]), .B(a[105]), .Z(n9023) );
  XNOR U19472 ( .A(n9028), .B(n8343), .Z(n8345) );
  XOR U19473 ( .A(n9029), .B(n9030), .Z(n8343) );
  ANDN U19474 ( .B(n9031), .A(n9032), .Z(n9029) );
  AND U19475 ( .A(b[9]), .B(a[106]), .Z(n9028) );
  XNOR U19476 ( .A(n9033), .B(n8348), .Z(n8350) );
  XOR U19477 ( .A(n9034), .B(n9035), .Z(n8348) );
  ANDN U19478 ( .B(n9036), .A(n9037), .Z(n9034) );
  AND U19479 ( .A(b[8]), .B(a[107]), .Z(n9033) );
  XNOR U19480 ( .A(n9038), .B(n8353), .Z(n8355) );
  XOR U19481 ( .A(n9039), .B(n9040), .Z(n8353) );
  ANDN U19482 ( .B(n9041), .A(n9042), .Z(n9039) );
  AND U19483 ( .A(b[7]), .B(a[108]), .Z(n9038) );
  XNOR U19484 ( .A(n9043), .B(n8358), .Z(n8360) );
  XOR U19485 ( .A(n9044), .B(n9045), .Z(n8358) );
  ANDN U19486 ( .B(n9046), .A(n9047), .Z(n9044) );
  AND U19487 ( .A(b[6]), .B(a[109]), .Z(n9043) );
  XNOR U19488 ( .A(n9048), .B(n8363), .Z(n8365) );
  XOR U19489 ( .A(n9049), .B(n9050), .Z(n8363) );
  ANDN U19490 ( .B(n9051), .A(n9052), .Z(n9049) );
  AND U19491 ( .A(b[5]), .B(a[110]), .Z(n9048) );
  XNOR U19492 ( .A(n9053), .B(n8368), .Z(n8370) );
  XOR U19493 ( .A(n9054), .B(n9055), .Z(n8368) );
  ANDN U19494 ( .B(n9056), .A(n9057), .Z(n9054) );
  AND U19495 ( .A(b[4]), .B(a[111]), .Z(n9053) );
  XNOR U19496 ( .A(n9058), .B(n9059), .Z(n8382) );
  NANDN U19497 ( .A(n9060), .B(n9061), .Z(n9059) );
  XNOR U19498 ( .A(n9062), .B(n8373), .Z(n8375) );
  XNOR U19499 ( .A(n9063), .B(n9064), .Z(n8373) );
  AND U19500 ( .A(n9065), .B(n9066), .Z(n9063) );
  AND U19501 ( .A(b[3]), .B(a[112]), .Z(n9062) );
  NAND U19502 ( .A(a[115]), .B(b[0]), .Z(n7700) );
  XNOR U19503 ( .A(n8388), .B(n8389), .Z(c[114]) );
  XNOR U19504 ( .A(n9060), .B(n9061), .Z(n8389) );
  XOR U19505 ( .A(n9058), .B(n9067), .Z(n9061) );
  NAND U19506 ( .A(b[1]), .B(a[113]), .Z(n9067) );
  XOR U19507 ( .A(n9066), .B(n9068), .Z(n9060) );
  XOR U19508 ( .A(n9058), .B(n9065), .Z(n9068) );
  XNOR U19509 ( .A(n9069), .B(n9064), .Z(n9065) );
  AND U19510 ( .A(b[2]), .B(a[112]), .Z(n9069) );
  NANDN U19511 ( .A(n9070), .B(n9071), .Z(n9058) );
  XOR U19512 ( .A(n9064), .B(n9056), .Z(n9072) );
  XNOR U19513 ( .A(n9055), .B(n9051), .Z(n9073) );
  XNOR U19514 ( .A(n9050), .B(n9046), .Z(n9074) );
  XNOR U19515 ( .A(n9045), .B(n9041), .Z(n9075) );
  XNOR U19516 ( .A(n9040), .B(n9036), .Z(n9076) );
  XNOR U19517 ( .A(n9035), .B(n9031), .Z(n9077) );
  XNOR U19518 ( .A(n9030), .B(n9026), .Z(n9078) );
  XNOR U19519 ( .A(n9025), .B(n9021), .Z(n9079) );
  XNOR U19520 ( .A(n9020), .B(n9016), .Z(n9080) );
  XNOR U19521 ( .A(n9015), .B(n9011), .Z(n9081) );
  XNOR U19522 ( .A(n9010), .B(n9006), .Z(n9082) );
  XNOR U19523 ( .A(n9005), .B(n9001), .Z(n9083) );
  XNOR U19524 ( .A(n9000), .B(n8996), .Z(n9084) );
  XNOR U19525 ( .A(n8995), .B(n8991), .Z(n9085) );
  XNOR U19526 ( .A(n8990), .B(n8986), .Z(n9086) );
  XNOR U19527 ( .A(n8985), .B(n8981), .Z(n9087) );
  XNOR U19528 ( .A(n8980), .B(n8976), .Z(n9088) );
  XNOR U19529 ( .A(n8975), .B(n8971), .Z(n9089) );
  XNOR U19530 ( .A(n8970), .B(n8966), .Z(n9090) );
  XNOR U19531 ( .A(n8965), .B(n8961), .Z(n9091) );
  XNOR U19532 ( .A(n8960), .B(n8956), .Z(n9092) );
  XNOR U19533 ( .A(n8955), .B(n8951), .Z(n9093) );
  XNOR U19534 ( .A(n8950), .B(n8946), .Z(n9094) );
  XNOR U19535 ( .A(n8945), .B(n8941), .Z(n9095) );
  XNOR U19536 ( .A(n8940), .B(n8936), .Z(n9096) );
  XNOR U19537 ( .A(n8935), .B(n8931), .Z(n9097) );
  XNOR U19538 ( .A(n8930), .B(n8926), .Z(n9098) );
  XNOR U19539 ( .A(n8925), .B(n8921), .Z(n9099) );
  XNOR U19540 ( .A(n8920), .B(n8916), .Z(n9100) );
  XNOR U19541 ( .A(n8915), .B(n8911), .Z(n9101) );
  XNOR U19542 ( .A(n8910), .B(n8906), .Z(n9102) );
  XNOR U19543 ( .A(n8905), .B(n8901), .Z(n9103) );
  XNOR U19544 ( .A(n8900), .B(n8896), .Z(n9104) );
  XNOR U19545 ( .A(n8895), .B(n8891), .Z(n9105) );
  XNOR U19546 ( .A(n8890), .B(n8886), .Z(n9106) );
  XNOR U19547 ( .A(n8885), .B(n8881), .Z(n9107) );
  XNOR U19548 ( .A(n8880), .B(n8876), .Z(n9108) );
  XNOR U19549 ( .A(n8875), .B(n8871), .Z(n9109) );
  XNOR U19550 ( .A(n8870), .B(n8866), .Z(n9110) );
  XNOR U19551 ( .A(n8865), .B(n8861), .Z(n9111) );
  XNOR U19552 ( .A(n8860), .B(n8856), .Z(n9112) );
  XNOR U19553 ( .A(n8855), .B(n8851), .Z(n9113) );
  XNOR U19554 ( .A(n8850), .B(n8846), .Z(n9114) );
  XNOR U19555 ( .A(n8845), .B(n8841), .Z(n9115) );
  XNOR U19556 ( .A(n8840), .B(n8836), .Z(n9116) );
  XNOR U19557 ( .A(n8835), .B(n8831), .Z(n9117) );
  XNOR U19558 ( .A(n8830), .B(n8826), .Z(n9118) );
  XNOR U19559 ( .A(n8825), .B(n8821), .Z(n9119) );
  XNOR U19560 ( .A(n8820), .B(n8816), .Z(n9120) );
  XNOR U19561 ( .A(n8815), .B(n8811), .Z(n9121) );
  XNOR U19562 ( .A(n8810), .B(n8806), .Z(n9122) );
  XNOR U19563 ( .A(n8805), .B(n8801), .Z(n9123) );
  XNOR U19564 ( .A(n8800), .B(n8796), .Z(n9124) );
  XNOR U19565 ( .A(n8795), .B(n8791), .Z(n9125) );
  XNOR U19566 ( .A(n8790), .B(n8786), .Z(n9126) );
  XNOR U19567 ( .A(n8785), .B(n8781), .Z(n9127) );
  XNOR U19568 ( .A(n8780), .B(n8776), .Z(n9128) );
  XNOR U19569 ( .A(n8775), .B(n8771), .Z(n9129) );
  XNOR U19570 ( .A(n8770), .B(n8766), .Z(n9130) );
  XNOR U19571 ( .A(n8765), .B(n8761), .Z(n9131) );
  XNOR U19572 ( .A(n8760), .B(n8756), .Z(n9132) );
  XNOR U19573 ( .A(n8755), .B(n8751), .Z(n9133) );
  XNOR U19574 ( .A(n8750), .B(n8746), .Z(n9134) );
  XNOR U19575 ( .A(n8745), .B(n8741), .Z(n9135) );
  XNOR U19576 ( .A(n8740), .B(n8736), .Z(n9136) );
  XNOR U19577 ( .A(n8735), .B(n8731), .Z(n9137) );
  XNOR U19578 ( .A(n8730), .B(n8726), .Z(n9138) );
  XNOR U19579 ( .A(n8725), .B(n8721), .Z(n9139) );
  XNOR U19580 ( .A(n8720), .B(n8716), .Z(n9140) );
  XNOR U19581 ( .A(n8715), .B(n8711), .Z(n9141) );
  XNOR U19582 ( .A(n8710), .B(n8706), .Z(n9142) );
  XNOR U19583 ( .A(n8705), .B(n8701), .Z(n9143) );
  XNOR U19584 ( .A(n8700), .B(n8696), .Z(n9144) );
  XNOR U19585 ( .A(n8695), .B(n8691), .Z(n9145) );
  XNOR U19586 ( .A(n8690), .B(n8686), .Z(n9146) );
  XNOR U19587 ( .A(n8685), .B(n8681), .Z(n9147) );
  XNOR U19588 ( .A(n8680), .B(n8676), .Z(n9148) );
  XNOR U19589 ( .A(n8675), .B(n8671), .Z(n9149) );
  XNOR U19590 ( .A(n8670), .B(n8666), .Z(n9150) );
  XNOR U19591 ( .A(n8665), .B(n8661), .Z(n9151) );
  XNOR U19592 ( .A(n8660), .B(n8656), .Z(n9152) );
  XNOR U19593 ( .A(n8655), .B(n8651), .Z(n9153) );
  XNOR U19594 ( .A(n8650), .B(n8646), .Z(n9154) );
  XNOR U19595 ( .A(n8645), .B(n8641), .Z(n9155) );
  XNOR U19596 ( .A(n8640), .B(n8636), .Z(n9156) );
  XNOR U19597 ( .A(n8635), .B(n8631), .Z(n9157) );
  XNOR U19598 ( .A(n8630), .B(n8626), .Z(n9158) );
  XNOR U19599 ( .A(n8625), .B(n8621), .Z(n9159) );
  XNOR U19600 ( .A(n8620), .B(n8616), .Z(n9160) );
  XNOR U19601 ( .A(n8615), .B(n8611), .Z(n9161) );
  XNOR U19602 ( .A(n8610), .B(n8606), .Z(n9162) );
  XNOR U19603 ( .A(n8605), .B(n8601), .Z(n9163) );
  XNOR U19604 ( .A(n8600), .B(n8596), .Z(n9164) );
  XNOR U19605 ( .A(n8595), .B(n8591), .Z(n9165) );
  XNOR U19606 ( .A(n8590), .B(n8586), .Z(n9166) );
  XNOR U19607 ( .A(n8585), .B(n8581), .Z(n9167) );
  XNOR U19608 ( .A(n8580), .B(n8576), .Z(n9168) );
  XNOR U19609 ( .A(n8575), .B(n8571), .Z(n9169) );
  XNOR U19610 ( .A(n8570), .B(n8566), .Z(n9170) );
  XNOR U19611 ( .A(n8565), .B(n8561), .Z(n9171) );
  XNOR U19612 ( .A(n8560), .B(n8556), .Z(n9172) );
  XNOR U19613 ( .A(n8555), .B(n8551), .Z(n9173) );
  XNOR U19614 ( .A(n8550), .B(n8546), .Z(n9174) );
  XNOR U19615 ( .A(n8545), .B(n8541), .Z(n9175) );
  XNOR U19616 ( .A(n8540), .B(n8536), .Z(n9176) );
  XNOR U19617 ( .A(n8535), .B(n8531), .Z(n9177) );
  XNOR U19618 ( .A(n8530), .B(n8526), .Z(n9178) );
  XNOR U19619 ( .A(n8525), .B(n8521), .Z(n9179) );
  XNOR U19620 ( .A(n8520), .B(n8516), .Z(n9180) );
  XNOR U19621 ( .A(n8515), .B(n8511), .Z(n9181) );
  XNOR U19622 ( .A(n8510), .B(n8506), .Z(n9182) );
  XOR U19623 ( .A(n9183), .B(n8505), .Z(n8506) );
  AND U19624 ( .A(a[0]), .B(b[114]), .Z(n9183) );
  XNOR U19625 ( .A(n9184), .B(n8505), .Z(n8507) );
  XNOR U19626 ( .A(n9185), .B(n9186), .Z(n8505) );
  ANDN U19627 ( .B(n9187), .A(n9188), .Z(n9185) );
  AND U19628 ( .A(a[1]), .B(b[113]), .Z(n9184) );
  XNOR U19629 ( .A(n9189), .B(n8510), .Z(n8512) );
  XOR U19630 ( .A(n9190), .B(n9191), .Z(n8510) );
  ANDN U19631 ( .B(n9192), .A(n9193), .Z(n9190) );
  AND U19632 ( .A(a[2]), .B(b[112]), .Z(n9189) );
  XNOR U19633 ( .A(n9194), .B(n8515), .Z(n8517) );
  XOR U19634 ( .A(n9195), .B(n9196), .Z(n8515) );
  ANDN U19635 ( .B(n9197), .A(n9198), .Z(n9195) );
  AND U19636 ( .A(a[3]), .B(b[111]), .Z(n9194) );
  XNOR U19637 ( .A(n9199), .B(n8520), .Z(n8522) );
  XOR U19638 ( .A(n9200), .B(n9201), .Z(n8520) );
  ANDN U19639 ( .B(n9202), .A(n9203), .Z(n9200) );
  AND U19640 ( .A(a[4]), .B(b[110]), .Z(n9199) );
  XNOR U19641 ( .A(n9204), .B(n8525), .Z(n8527) );
  XOR U19642 ( .A(n9205), .B(n9206), .Z(n8525) );
  ANDN U19643 ( .B(n9207), .A(n9208), .Z(n9205) );
  AND U19644 ( .A(a[5]), .B(b[109]), .Z(n9204) );
  XNOR U19645 ( .A(n9209), .B(n8530), .Z(n8532) );
  XOR U19646 ( .A(n9210), .B(n9211), .Z(n8530) );
  ANDN U19647 ( .B(n9212), .A(n9213), .Z(n9210) );
  AND U19648 ( .A(a[6]), .B(b[108]), .Z(n9209) );
  XNOR U19649 ( .A(n9214), .B(n8535), .Z(n8537) );
  XOR U19650 ( .A(n9215), .B(n9216), .Z(n8535) );
  ANDN U19651 ( .B(n9217), .A(n9218), .Z(n9215) );
  AND U19652 ( .A(a[7]), .B(b[107]), .Z(n9214) );
  XNOR U19653 ( .A(n9219), .B(n8540), .Z(n8542) );
  XOR U19654 ( .A(n9220), .B(n9221), .Z(n8540) );
  ANDN U19655 ( .B(n9222), .A(n9223), .Z(n9220) );
  AND U19656 ( .A(a[8]), .B(b[106]), .Z(n9219) );
  XNOR U19657 ( .A(n9224), .B(n8545), .Z(n8547) );
  XOR U19658 ( .A(n9225), .B(n9226), .Z(n8545) );
  ANDN U19659 ( .B(n9227), .A(n9228), .Z(n9225) );
  AND U19660 ( .A(a[9]), .B(b[105]), .Z(n9224) );
  XNOR U19661 ( .A(n9229), .B(n8550), .Z(n8552) );
  XOR U19662 ( .A(n9230), .B(n9231), .Z(n8550) );
  ANDN U19663 ( .B(n9232), .A(n9233), .Z(n9230) );
  AND U19664 ( .A(a[10]), .B(b[104]), .Z(n9229) );
  XNOR U19665 ( .A(n9234), .B(n8555), .Z(n8557) );
  XOR U19666 ( .A(n9235), .B(n9236), .Z(n8555) );
  ANDN U19667 ( .B(n9237), .A(n9238), .Z(n9235) );
  AND U19668 ( .A(a[11]), .B(b[103]), .Z(n9234) );
  XNOR U19669 ( .A(n9239), .B(n8560), .Z(n8562) );
  XOR U19670 ( .A(n9240), .B(n9241), .Z(n8560) );
  ANDN U19671 ( .B(n9242), .A(n9243), .Z(n9240) );
  AND U19672 ( .A(a[12]), .B(b[102]), .Z(n9239) );
  XNOR U19673 ( .A(n9244), .B(n8565), .Z(n8567) );
  XOR U19674 ( .A(n9245), .B(n9246), .Z(n8565) );
  ANDN U19675 ( .B(n9247), .A(n9248), .Z(n9245) );
  AND U19676 ( .A(a[13]), .B(b[101]), .Z(n9244) );
  XNOR U19677 ( .A(n9249), .B(n8570), .Z(n8572) );
  XOR U19678 ( .A(n9250), .B(n9251), .Z(n8570) );
  ANDN U19679 ( .B(n9252), .A(n9253), .Z(n9250) );
  AND U19680 ( .A(a[14]), .B(b[100]), .Z(n9249) );
  XNOR U19681 ( .A(n9254), .B(n8575), .Z(n8577) );
  XOR U19682 ( .A(n9255), .B(n9256), .Z(n8575) );
  ANDN U19683 ( .B(n9257), .A(n9258), .Z(n9255) );
  AND U19684 ( .A(a[15]), .B(b[99]), .Z(n9254) );
  XNOR U19685 ( .A(n9259), .B(n8580), .Z(n8582) );
  XOR U19686 ( .A(n9260), .B(n9261), .Z(n8580) );
  ANDN U19687 ( .B(n9262), .A(n9263), .Z(n9260) );
  AND U19688 ( .A(a[16]), .B(b[98]), .Z(n9259) );
  XNOR U19689 ( .A(n9264), .B(n8585), .Z(n8587) );
  XOR U19690 ( .A(n9265), .B(n9266), .Z(n8585) );
  ANDN U19691 ( .B(n9267), .A(n9268), .Z(n9265) );
  AND U19692 ( .A(a[17]), .B(b[97]), .Z(n9264) );
  XNOR U19693 ( .A(n9269), .B(n8590), .Z(n8592) );
  XOR U19694 ( .A(n9270), .B(n9271), .Z(n8590) );
  ANDN U19695 ( .B(n9272), .A(n9273), .Z(n9270) );
  AND U19696 ( .A(a[18]), .B(b[96]), .Z(n9269) );
  XNOR U19697 ( .A(n9274), .B(n8595), .Z(n8597) );
  XOR U19698 ( .A(n9275), .B(n9276), .Z(n8595) );
  ANDN U19699 ( .B(n9277), .A(n9278), .Z(n9275) );
  AND U19700 ( .A(a[19]), .B(b[95]), .Z(n9274) );
  XNOR U19701 ( .A(n9279), .B(n8600), .Z(n8602) );
  XOR U19702 ( .A(n9280), .B(n9281), .Z(n8600) );
  ANDN U19703 ( .B(n9282), .A(n9283), .Z(n9280) );
  AND U19704 ( .A(a[20]), .B(b[94]), .Z(n9279) );
  XNOR U19705 ( .A(n9284), .B(n8605), .Z(n8607) );
  XOR U19706 ( .A(n9285), .B(n9286), .Z(n8605) );
  ANDN U19707 ( .B(n9287), .A(n9288), .Z(n9285) );
  AND U19708 ( .A(a[21]), .B(b[93]), .Z(n9284) );
  XNOR U19709 ( .A(n9289), .B(n8610), .Z(n8612) );
  XOR U19710 ( .A(n9290), .B(n9291), .Z(n8610) );
  ANDN U19711 ( .B(n9292), .A(n9293), .Z(n9290) );
  AND U19712 ( .A(a[22]), .B(b[92]), .Z(n9289) );
  XNOR U19713 ( .A(n9294), .B(n8615), .Z(n8617) );
  XOR U19714 ( .A(n9295), .B(n9296), .Z(n8615) );
  ANDN U19715 ( .B(n9297), .A(n9298), .Z(n9295) );
  AND U19716 ( .A(a[23]), .B(b[91]), .Z(n9294) );
  XNOR U19717 ( .A(n9299), .B(n8620), .Z(n8622) );
  XOR U19718 ( .A(n9300), .B(n9301), .Z(n8620) );
  ANDN U19719 ( .B(n9302), .A(n9303), .Z(n9300) );
  AND U19720 ( .A(a[24]), .B(b[90]), .Z(n9299) );
  XNOR U19721 ( .A(n9304), .B(n8625), .Z(n8627) );
  XOR U19722 ( .A(n9305), .B(n9306), .Z(n8625) );
  ANDN U19723 ( .B(n9307), .A(n9308), .Z(n9305) );
  AND U19724 ( .A(a[25]), .B(b[89]), .Z(n9304) );
  XNOR U19725 ( .A(n9309), .B(n8630), .Z(n8632) );
  XOR U19726 ( .A(n9310), .B(n9311), .Z(n8630) );
  ANDN U19727 ( .B(n9312), .A(n9313), .Z(n9310) );
  AND U19728 ( .A(a[26]), .B(b[88]), .Z(n9309) );
  XNOR U19729 ( .A(n9314), .B(n8635), .Z(n8637) );
  XOR U19730 ( .A(n9315), .B(n9316), .Z(n8635) );
  ANDN U19731 ( .B(n9317), .A(n9318), .Z(n9315) );
  AND U19732 ( .A(a[27]), .B(b[87]), .Z(n9314) );
  XNOR U19733 ( .A(n9319), .B(n8640), .Z(n8642) );
  XOR U19734 ( .A(n9320), .B(n9321), .Z(n8640) );
  ANDN U19735 ( .B(n9322), .A(n9323), .Z(n9320) );
  AND U19736 ( .A(a[28]), .B(b[86]), .Z(n9319) );
  XNOR U19737 ( .A(n9324), .B(n8645), .Z(n8647) );
  XOR U19738 ( .A(n9325), .B(n9326), .Z(n8645) );
  ANDN U19739 ( .B(n9327), .A(n9328), .Z(n9325) );
  AND U19740 ( .A(a[29]), .B(b[85]), .Z(n9324) );
  XNOR U19741 ( .A(n9329), .B(n8650), .Z(n8652) );
  XOR U19742 ( .A(n9330), .B(n9331), .Z(n8650) );
  ANDN U19743 ( .B(n9332), .A(n9333), .Z(n9330) );
  AND U19744 ( .A(a[30]), .B(b[84]), .Z(n9329) );
  XNOR U19745 ( .A(n9334), .B(n8655), .Z(n8657) );
  XOR U19746 ( .A(n9335), .B(n9336), .Z(n8655) );
  ANDN U19747 ( .B(n9337), .A(n9338), .Z(n9335) );
  AND U19748 ( .A(a[31]), .B(b[83]), .Z(n9334) );
  XNOR U19749 ( .A(n9339), .B(n8660), .Z(n8662) );
  XOR U19750 ( .A(n9340), .B(n9341), .Z(n8660) );
  ANDN U19751 ( .B(n9342), .A(n9343), .Z(n9340) );
  AND U19752 ( .A(a[32]), .B(b[82]), .Z(n9339) );
  XNOR U19753 ( .A(n9344), .B(n8665), .Z(n8667) );
  XOR U19754 ( .A(n9345), .B(n9346), .Z(n8665) );
  ANDN U19755 ( .B(n9347), .A(n9348), .Z(n9345) );
  AND U19756 ( .A(a[33]), .B(b[81]), .Z(n9344) );
  XNOR U19757 ( .A(n9349), .B(n8670), .Z(n8672) );
  XOR U19758 ( .A(n9350), .B(n9351), .Z(n8670) );
  ANDN U19759 ( .B(n9352), .A(n9353), .Z(n9350) );
  AND U19760 ( .A(a[34]), .B(b[80]), .Z(n9349) );
  XNOR U19761 ( .A(n9354), .B(n8675), .Z(n8677) );
  XOR U19762 ( .A(n9355), .B(n9356), .Z(n8675) );
  ANDN U19763 ( .B(n9357), .A(n9358), .Z(n9355) );
  AND U19764 ( .A(a[35]), .B(b[79]), .Z(n9354) );
  XNOR U19765 ( .A(n9359), .B(n8680), .Z(n8682) );
  XOR U19766 ( .A(n9360), .B(n9361), .Z(n8680) );
  ANDN U19767 ( .B(n9362), .A(n9363), .Z(n9360) );
  AND U19768 ( .A(a[36]), .B(b[78]), .Z(n9359) );
  XNOR U19769 ( .A(n9364), .B(n8685), .Z(n8687) );
  XOR U19770 ( .A(n9365), .B(n9366), .Z(n8685) );
  ANDN U19771 ( .B(n9367), .A(n9368), .Z(n9365) );
  AND U19772 ( .A(a[37]), .B(b[77]), .Z(n9364) );
  XNOR U19773 ( .A(n9369), .B(n8690), .Z(n8692) );
  XOR U19774 ( .A(n9370), .B(n9371), .Z(n8690) );
  ANDN U19775 ( .B(n9372), .A(n9373), .Z(n9370) );
  AND U19776 ( .A(a[38]), .B(b[76]), .Z(n9369) );
  XNOR U19777 ( .A(n9374), .B(n8695), .Z(n8697) );
  XOR U19778 ( .A(n9375), .B(n9376), .Z(n8695) );
  ANDN U19779 ( .B(n9377), .A(n9378), .Z(n9375) );
  AND U19780 ( .A(a[39]), .B(b[75]), .Z(n9374) );
  XNOR U19781 ( .A(n9379), .B(n8700), .Z(n8702) );
  XOR U19782 ( .A(n9380), .B(n9381), .Z(n8700) );
  ANDN U19783 ( .B(n9382), .A(n9383), .Z(n9380) );
  AND U19784 ( .A(a[40]), .B(b[74]), .Z(n9379) );
  XNOR U19785 ( .A(n9384), .B(n8705), .Z(n8707) );
  XOR U19786 ( .A(n9385), .B(n9386), .Z(n8705) );
  ANDN U19787 ( .B(n9387), .A(n9388), .Z(n9385) );
  AND U19788 ( .A(a[41]), .B(b[73]), .Z(n9384) );
  XNOR U19789 ( .A(n9389), .B(n8710), .Z(n8712) );
  XOR U19790 ( .A(n9390), .B(n9391), .Z(n8710) );
  ANDN U19791 ( .B(n9392), .A(n9393), .Z(n9390) );
  AND U19792 ( .A(a[42]), .B(b[72]), .Z(n9389) );
  XNOR U19793 ( .A(n9394), .B(n8715), .Z(n8717) );
  XOR U19794 ( .A(n9395), .B(n9396), .Z(n8715) );
  ANDN U19795 ( .B(n9397), .A(n9398), .Z(n9395) );
  AND U19796 ( .A(a[43]), .B(b[71]), .Z(n9394) );
  XNOR U19797 ( .A(n9399), .B(n8720), .Z(n8722) );
  XOR U19798 ( .A(n9400), .B(n9401), .Z(n8720) );
  ANDN U19799 ( .B(n9402), .A(n9403), .Z(n9400) );
  AND U19800 ( .A(a[44]), .B(b[70]), .Z(n9399) );
  XNOR U19801 ( .A(n9404), .B(n8725), .Z(n8727) );
  XOR U19802 ( .A(n9405), .B(n9406), .Z(n8725) );
  ANDN U19803 ( .B(n9407), .A(n9408), .Z(n9405) );
  AND U19804 ( .A(a[45]), .B(b[69]), .Z(n9404) );
  XNOR U19805 ( .A(n9409), .B(n8730), .Z(n8732) );
  XOR U19806 ( .A(n9410), .B(n9411), .Z(n8730) );
  ANDN U19807 ( .B(n9412), .A(n9413), .Z(n9410) );
  AND U19808 ( .A(a[46]), .B(b[68]), .Z(n9409) );
  XNOR U19809 ( .A(n9414), .B(n8735), .Z(n8737) );
  XOR U19810 ( .A(n9415), .B(n9416), .Z(n8735) );
  ANDN U19811 ( .B(n9417), .A(n9418), .Z(n9415) );
  AND U19812 ( .A(a[47]), .B(b[67]), .Z(n9414) );
  XNOR U19813 ( .A(n9419), .B(n8740), .Z(n8742) );
  XOR U19814 ( .A(n9420), .B(n9421), .Z(n8740) );
  ANDN U19815 ( .B(n9422), .A(n9423), .Z(n9420) );
  AND U19816 ( .A(a[48]), .B(b[66]), .Z(n9419) );
  XNOR U19817 ( .A(n9424), .B(n8745), .Z(n8747) );
  XOR U19818 ( .A(n9425), .B(n9426), .Z(n8745) );
  ANDN U19819 ( .B(n9427), .A(n9428), .Z(n9425) );
  AND U19820 ( .A(a[49]), .B(b[65]), .Z(n9424) );
  XNOR U19821 ( .A(n9429), .B(n8750), .Z(n8752) );
  XOR U19822 ( .A(n9430), .B(n9431), .Z(n8750) );
  ANDN U19823 ( .B(n9432), .A(n9433), .Z(n9430) );
  AND U19824 ( .A(a[50]), .B(b[64]), .Z(n9429) );
  XNOR U19825 ( .A(n9434), .B(n8755), .Z(n8757) );
  XOR U19826 ( .A(n9435), .B(n9436), .Z(n8755) );
  ANDN U19827 ( .B(n9437), .A(n9438), .Z(n9435) );
  AND U19828 ( .A(a[51]), .B(b[63]), .Z(n9434) );
  XNOR U19829 ( .A(n9439), .B(n8760), .Z(n8762) );
  XOR U19830 ( .A(n9440), .B(n9441), .Z(n8760) );
  ANDN U19831 ( .B(n9442), .A(n9443), .Z(n9440) );
  AND U19832 ( .A(a[52]), .B(b[62]), .Z(n9439) );
  XNOR U19833 ( .A(n9444), .B(n8765), .Z(n8767) );
  XOR U19834 ( .A(n9445), .B(n9446), .Z(n8765) );
  ANDN U19835 ( .B(n9447), .A(n9448), .Z(n9445) );
  AND U19836 ( .A(a[53]), .B(b[61]), .Z(n9444) );
  XNOR U19837 ( .A(n9449), .B(n8770), .Z(n8772) );
  XOR U19838 ( .A(n9450), .B(n9451), .Z(n8770) );
  ANDN U19839 ( .B(n9452), .A(n9453), .Z(n9450) );
  AND U19840 ( .A(a[54]), .B(b[60]), .Z(n9449) );
  XNOR U19841 ( .A(n9454), .B(n8775), .Z(n8777) );
  XOR U19842 ( .A(n9455), .B(n9456), .Z(n8775) );
  ANDN U19843 ( .B(n9457), .A(n9458), .Z(n9455) );
  AND U19844 ( .A(a[55]), .B(b[59]), .Z(n9454) );
  XNOR U19845 ( .A(n9459), .B(n8780), .Z(n8782) );
  XOR U19846 ( .A(n9460), .B(n9461), .Z(n8780) );
  ANDN U19847 ( .B(n9462), .A(n9463), .Z(n9460) );
  AND U19848 ( .A(a[56]), .B(b[58]), .Z(n9459) );
  XNOR U19849 ( .A(n9464), .B(n8785), .Z(n8787) );
  XOR U19850 ( .A(n9465), .B(n9466), .Z(n8785) );
  ANDN U19851 ( .B(n9467), .A(n9468), .Z(n9465) );
  AND U19852 ( .A(a[57]), .B(b[57]), .Z(n9464) );
  XNOR U19853 ( .A(n9469), .B(n8790), .Z(n8792) );
  XOR U19854 ( .A(n9470), .B(n9471), .Z(n8790) );
  ANDN U19855 ( .B(n9472), .A(n9473), .Z(n9470) );
  AND U19856 ( .A(a[58]), .B(b[56]), .Z(n9469) );
  XNOR U19857 ( .A(n9474), .B(n8795), .Z(n8797) );
  XOR U19858 ( .A(n9475), .B(n9476), .Z(n8795) );
  ANDN U19859 ( .B(n9477), .A(n9478), .Z(n9475) );
  AND U19860 ( .A(a[59]), .B(b[55]), .Z(n9474) );
  XNOR U19861 ( .A(n9479), .B(n8800), .Z(n8802) );
  XOR U19862 ( .A(n9480), .B(n9481), .Z(n8800) );
  ANDN U19863 ( .B(n9482), .A(n9483), .Z(n9480) );
  AND U19864 ( .A(a[60]), .B(b[54]), .Z(n9479) );
  XNOR U19865 ( .A(n9484), .B(n8805), .Z(n8807) );
  XOR U19866 ( .A(n9485), .B(n9486), .Z(n8805) );
  ANDN U19867 ( .B(n9487), .A(n9488), .Z(n9485) );
  AND U19868 ( .A(a[61]), .B(b[53]), .Z(n9484) );
  XNOR U19869 ( .A(n9489), .B(n8810), .Z(n8812) );
  XOR U19870 ( .A(n9490), .B(n9491), .Z(n8810) );
  ANDN U19871 ( .B(n9492), .A(n9493), .Z(n9490) );
  AND U19872 ( .A(a[62]), .B(b[52]), .Z(n9489) );
  XNOR U19873 ( .A(n9494), .B(n8815), .Z(n8817) );
  XOR U19874 ( .A(n9495), .B(n9496), .Z(n8815) );
  ANDN U19875 ( .B(n9497), .A(n9498), .Z(n9495) );
  AND U19876 ( .A(a[63]), .B(b[51]), .Z(n9494) );
  XNOR U19877 ( .A(n9499), .B(n8820), .Z(n8822) );
  XOR U19878 ( .A(n9500), .B(n9501), .Z(n8820) );
  ANDN U19879 ( .B(n9502), .A(n9503), .Z(n9500) );
  AND U19880 ( .A(a[64]), .B(b[50]), .Z(n9499) );
  XNOR U19881 ( .A(n9504), .B(n8825), .Z(n8827) );
  XOR U19882 ( .A(n9505), .B(n9506), .Z(n8825) );
  ANDN U19883 ( .B(n9507), .A(n9508), .Z(n9505) );
  AND U19884 ( .A(a[65]), .B(b[49]), .Z(n9504) );
  XNOR U19885 ( .A(n9509), .B(n8830), .Z(n8832) );
  XOR U19886 ( .A(n9510), .B(n9511), .Z(n8830) );
  ANDN U19887 ( .B(n9512), .A(n9513), .Z(n9510) );
  AND U19888 ( .A(a[66]), .B(b[48]), .Z(n9509) );
  XNOR U19889 ( .A(n9514), .B(n8835), .Z(n8837) );
  XOR U19890 ( .A(n9515), .B(n9516), .Z(n8835) );
  ANDN U19891 ( .B(n9517), .A(n9518), .Z(n9515) );
  AND U19892 ( .A(a[67]), .B(b[47]), .Z(n9514) );
  XNOR U19893 ( .A(n9519), .B(n8840), .Z(n8842) );
  XOR U19894 ( .A(n9520), .B(n9521), .Z(n8840) );
  ANDN U19895 ( .B(n9522), .A(n9523), .Z(n9520) );
  AND U19896 ( .A(a[68]), .B(b[46]), .Z(n9519) );
  XNOR U19897 ( .A(n9524), .B(n8845), .Z(n8847) );
  XOR U19898 ( .A(n9525), .B(n9526), .Z(n8845) );
  ANDN U19899 ( .B(n9527), .A(n9528), .Z(n9525) );
  AND U19900 ( .A(a[69]), .B(b[45]), .Z(n9524) );
  XNOR U19901 ( .A(n9529), .B(n8850), .Z(n8852) );
  XOR U19902 ( .A(n9530), .B(n9531), .Z(n8850) );
  ANDN U19903 ( .B(n9532), .A(n9533), .Z(n9530) );
  AND U19904 ( .A(a[70]), .B(b[44]), .Z(n9529) );
  XNOR U19905 ( .A(n9534), .B(n8855), .Z(n8857) );
  XOR U19906 ( .A(n9535), .B(n9536), .Z(n8855) );
  ANDN U19907 ( .B(n9537), .A(n9538), .Z(n9535) );
  AND U19908 ( .A(a[71]), .B(b[43]), .Z(n9534) );
  XNOR U19909 ( .A(n9539), .B(n8860), .Z(n8862) );
  XOR U19910 ( .A(n9540), .B(n9541), .Z(n8860) );
  ANDN U19911 ( .B(n9542), .A(n9543), .Z(n9540) );
  AND U19912 ( .A(a[72]), .B(b[42]), .Z(n9539) );
  XNOR U19913 ( .A(n9544), .B(n8865), .Z(n8867) );
  XOR U19914 ( .A(n9545), .B(n9546), .Z(n8865) );
  ANDN U19915 ( .B(n9547), .A(n9548), .Z(n9545) );
  AND U19916 ( .A(a[73]), .B(b[41]), .Z(n9544) );
  XNOR U19917 ( .A(n9549), .B(n8870), .Z(n8872) );
  XOR U19918 ( .A(n9550), .B(n9551), .Z(n8870) );
  ANDN U19919 ( .B(n9552), .A(n9553), .Z(n9550) );
  AND U19920 ( .A(a[74]), .B(b[40]), .Z(n9549) );
  XNOR U19921 ( .A(n9554), .B(n8875), .Z(n8877) );
  XOR U19922 ( .A(n9555), .B(n9556), .Z(n8875) );
  ANDN U19923 ( .B(n9557), .A(n9558), .Z(n9555) );
  AND U19924 ( .A(a[75]), .B(b[39]), .Z(n9554) );
  XNOR U19925 ( .A(n9559), .B(n8880), .Z(n8882) );
  XOR U19926 ( .A(n9560), .B(n9561), .Z(n8880) );
  ANDN U19927 ( .B(n9562), .A(n9563), .Z(n9560) );
  AND U19928 ( .A(a[76]), .B(b[38]), .Z(n9559) );
  XNOR U19929 ( .A(n9564), .B(n8885), .Z(n8887) );
  XOR U19930 ( .A(n9565), .B(n9566), .Z(n8885) );
  ANDN U19931 ( .B(n9567), .A(n9568), .Z(n9565) );
  AND U19932 ( .A(a[77]), .B(b[37]), .Z(n9564) );
  XNOR U19933 ( .A(n9569), .B(n8890), .Z(n8892) );
  XOR U19934 ( .A(n9570), .B(n9571), .Z(n8890) );
  ANDN U19935 ( .B(n9572), .A(n9573), .Z(n9570) );
  AND U19936 ( .A(a[78]), .B(b[36]), .Z(n9569) );
  XNOR U19937 ( .A(n9574), .B(n8895), .Z(n8897) );
  XOR U19938 ( .A(n9575), .B(n9576), .Z(n8895) );
  ANDN U19939 ( .B(n9577), .A(n9578), .Z(n9575) );
  AND U19940 ( .A(a[79]), .B(b[35]), .Z(n9574) );
  XNOR U19941 ( .A(n9579), .B(n8900), .Z(n8902) );
  XOR U19942 ( .A(n9580), .B(n9581), .Z(n8900) );
  ANDN U19943 ( .B(n9582), .A(n9583), .Z(n9580) );
  AND U19944 ( .A(a[80]), .B(b[34]), .Z(n9579) );
  XNOR U19945 ( .A(n9584), .B(n8905), .Z(n8907) );
  XOR U19946 ( .A(n9585), .B(n9586), .Z(n8905) );
  ANDN U19947 ( .B(n9587), .A(n9588), .Z(n9585) );
  AND U19948 ( .A(a[81]), .B(b[33]), .Z(n9584) );
  XNOR U19949 ( .A(n9589), .B(n8910), .Z(n8912) );
  XOR U19950 ( .A(n9590), .B(n9591), .Z(n8910) );
  ANDN U19951 ( .B(n9592), .A(n9593), .Z(n9590) );
  AND U19952 ( .A(a[82]), .B(b[32]), .Z(n9589) );
  XNOR U19953 ( .A(n9594), .B(n8915), .Z(n8917) );
  XOR U19954 ( .A(n9595), .B(n9596), .Z(n8915) );
  ANDN U19955 ( .B(n9597), .A(n9598), .Z(n9595) );
  AND U19956 ( .A(a[83]), .B(b[31]), .Z(n9594) );
  XNOR U19957 ( .A(n9599), .B(n8920), .Z(n8922) );
  XOR U19958 ( .A(n9600), .B(n9601), .Z(n8920) );
  ANDN U19959 ( .B(n9602), .A(n9603), .Z(n9600) );
  AND U19960 ( .A(a[84]), .B(b[30]), .Z(n9599) );
  XNOR U19961 ( .A(n9604), .B(n8925), .Z(n8927) );
  XOR U19962 ( .A(n9605), .B(n9606), .Z(n8925) );
  ANDN U19963 ( .B(n9607), .A(n9608), .Z(n9605) );
  AND U19964 ( .A(a[85]), .B(b[29]), .Z(n9604) );
  XNOR U19965 ( .A(n9609), .B(n8930), .Z(n8932) );
  XOR U19966 ( .A(n9610), .B(n9611), .Z(n8930) );
  ANDN U19967 ( .B(n9612), .A(n9613), .Z(n9610) );
  AND U19968 ( .A(a[86]), .B(b[28]), .Z(n9609) );
  XNOR U19969 ( .A(n9614), .B(n8935), .Z(n8937) );
  XOR U19970 ( .A(n9615), .B(n9616), .Z(n8935) );
  ANDN U19971 ( .B(n9617), .A(n9618), .Z(n9615) );
  AND U19972 ( .A(a[87]), .B(b[27]), .Z(n9614) );
  XNOR U19973 ( .A(n9619), .B(n8940), .Z(n8942) );
  XOR U19974 ( .A(n9620), .B(n9621), .Z(n8940) );
  ANDN U19975 ( .B(n9622), .A(n9623), .Z(n9620) );
  AND U19976 ( .A(a[88]), .B(b[26]), .Z(n9619) );
  XNOR U19977 ( .A(n9624), .B(n8945), .Z(n8947) );
  XOR U19978 ( .A(n9625), .B(n9626), .Z(n8945) );
  ANDN U19979 ( .B(n9627), .A(n9628), .Z(n9625) );
  AND U19980 ( .A(a[89]), .B(b[25]), .Z(n9624) );
  XNOR U19981 ( .A(n9629), .B(n8950), .Z(n8952) );
  XOR U19982 ( .A(n9630), .B(n9631), .Z(n8950) );
  ANDN U19983 ( .B(n9632), .A(n9633), .Z(n9630) );
  AND U19984 ( .A(a[90]), .B(b[24]), .Z(n9629) );
  XNOR U19985 ( .A(n9634), .B(n8955), .Z(n8957) );
  XOR U19986 ( .A(n9635), .B(n9636), .Z(n8955) );
  ANDN U19987 ( .B(n9637), .A(n9638), .Z(n9635) );
  AND U19988 ( .A(a[91]), .B(b[23]), .Z(n9634) );
  XNOR U19989 ( .A(n9639), .B(n8960), .Z(n8962) );
  XOR U19990 ( .A(n9640), .B(n9641), .Z(n8960) );
  ANDN U19991 ( .B(n9642), .A(n9643), .Z(n9640) );
  AND U19992 ( .A(a[92]), .B(b[22]), .Z(n9639) );
  XNOR U19993 ( .A(n9644), .B(n8965), .Z(n8967) );
  XOR U19994 ( .A(n9645), .B(n9646), .Z(n8965) );
  ANDN U19995 ( .B(n9647), .A(n9648), .Z(n9645) );
  AND U19996 ( .A(a[93]), .B(b[21]), .Z(n9644) );
  XNOR U19997 ( .A(n9649), .B(n8970), .Z(n8972) );
  XOR U19998 ( .A(n9650), .B(n9651), .Z(n8970) );
  ANDN U19999 ( .B(n9652), .A(n9653), .Z(n9650) );
  AND U20000 ( .A(a[94]), .B(b[20]), .Z(n9649) );
  XNOR U20001 ( .A(n9654), .B(n8975), .Z(n8977) );
  XOR U20002 ( .A(n9655), .B(n9656), .Z(n8975) );
  ANDN U20003 ( .B(n9657), .A(n9658), .Z(n9655) );
  AND U20004 ( .A(a[95]), .B(b[19]), .Z(n9654) );
  XNOR U20005 ( .A(n9659), .B(n8980), .Z(n8982) );
  XOR U20006 ( .A(n9660), .B(n9661), .Z(n8980) );
  ANDN U20007 ( .B(n9662), .A(n9663), .Z(n9660) );
  AND U20008 ( .A(a[96]), .B(b[18]), .Z(n9659) );
  XNOR U20009 ( .A(n9664), .B(n8985), .Z(n8987) );
  XOR U20010 ( .A(n9665), .B(n9666), .Z(n8985) );
  ANDN U20011 ( .B(n9667), .A(n9668), .Z(n9665) );
  AND U20012 ( .A(a[97]), .B(b[17]), .Z(n9664) );
  XNOR U20013 ( .A(n9669), .B(n8990), .Z(n8992) );
  XOR U20014 ( .A(n9670), .B(n9671), .Z(n8990) );
  ANDN U20015 ( .B(n9672), .A(n9673), .Z(n9670) );
  AND U20016 ( .A(a[98]), .B(b[16]), .Z(n9669) );
  XNOR U20017 ( .A(n9674), .B(n8995), .Z(n8997) );
  XOR U20018 ( .A(n9675), .B(n9676), .Z(n8995) );
  ANDN U20019 ( .B(n9677), .A(n9678), .Z(n9675) );
  AND U20020 ( .A(a[99]), .B(b[15]), .Z(n9674) );
  XNOR U20021 ( .A(n9679), .B(n9000), .Z(n9002) );
  XOR U20022 ( .A(n9680), .B(n9681), .Z(n9000) );
  ANDN U20023 ( .B(n9682), .A(n9683), .Z(n9680) );
  AND U20024 ( .A(b[14]), .B(a[100]), .Z(n9679) );
  XNOR U20025 ( .A(n9684), .B(n9005), .Z(n9007) );
  XOR U20026 ( .A(n9685), .B(n9686), .Z(n9005) );
  ANDN U20027 ( .B(n9687), .A(n9688), .Z(n9685) );
  AND U20028 ( .A(b[13]), .B(a[101]), .Z(n9684) );
  XNOR U20029 ( .A(n9689), .B(n9010), .Z(n9012) );
  XOR U20030 ( .A(n9690), .B(n9691), .Z(n9010) );
  ANDN U20031 ( .B(n9692), .A(n9693), .Z(n9690) );
  AND U20032 ( .A(b[12]), .B(a[102]), .Z(n9689) );
  XNOR U20033 ( .A(n9694), .B(n9015), .Z(n9017) );
  XOR U20034 ( .A(n9695), .B(n9696), .Z(n9015) );
  ANDN U20035 ( .B(n9697), .A(n9698), .Z(n9695) );
  AND U20036 ( .A(b[11]), .B(a[103]), .Z(n9694) );
  XNOR U20037 ( .A(n9699), .B(n9020), .Z(n9022) );
  XOR U20038 ( .A(n9700), .B(n9701), .Z(n9020) );
  ANDN U20039 ( .B(n9702), .A(n9703), .Z(n9700) );
  AND U20040 ( .A(b[10]), .B(a[104]), .Z(n9699) );
  XNOR U20041 ( .A(n9704), .B(n9025), .Z(n9027) );
  XOR U20042 ( .A(n9705), .B(n9706), .Z(n9025) );
  ANDN U20043 ( .B(n9707), .A(n9708), .Z(n9705) );
  AND U20044 ( .A(b[9]), .B(a[105]), .Z(n9704) );
  XNOR U20045 ( .A(n9709), .B(n9030), .Z(n9032) );
  XOR U20046 ( .A(n9710), .B(n9711), .Z(n9030) );
  ANDN U20047 ( .B(n9712), .A(n9713), .Z(n9710) );
  AND U20048 ( .A(b[8]), .B(a[106]), .Z(n9709) );
  XNOR U20049 ( .A(n9714), .B(n9035), .Z(n9037) );
  XOR U20050 ( .A(n9715), .B(n9716), .Z(n9035) );
  ANDN U20051 ( .B(n9717), .A(n9718), .Z(n9715) );
  AND U20052 ( .A(b[7]), .B(a[107]), .Z(n9714) );
  XNOR U20053 ( .A(n9719), .B(n9040), .Z(n9042) );
  XOR U20054 ( .A(n9720), .B(n9721), .Z(n9040) );
  ANDN U20055 ( .B(n9722), .A(n9723), .Z(n9720) );
  AND U20056 ( .A(b[6]), .B(a[108]), .Z(n9719) );
  XNOR U20057 ( .A(n9724), .B(n9045), .Z(n9047) );
  XOR U20058 ( .A(n9725), .B(n9726), .Z(n9045) );
  ANDN U20059 ( .B(n9727), .A(n9728), .Z(n9725) );
  AND U20060 ( .A(b[5]), .B(a[109]), .Z(n9724) );
  XNOR U20061 ( .A(n9729), .B(n9050), .Z(n9052) );
  XOR U20062 ( .A(n9730), .B(n9731), .Z(n9050) );
  ANDN U20063 ( .B(n9732), .A(n9733), .Z(n9730) );
  AND U20064 ( .A(b[4]), .B(a[110]), .Z(n9729) );
  XNOR U20065 ( .A(n9734), .B(n9735), .Z(n9064) );
  NANDN U20066 ( .A(n9736), .B(n9737), .Z(n9735) );
  XNOR U20067 ( .A(n9738), .B(n9055), .Z(n9057) );
  XNOR U20068 ( .A(n9739), .B(n9740), .Z(n9055) );
  AND U20069 ( .A(n9741), .B(n9742), .Z(n9739) );
  AND U20070 ( .A(b[3]), .B(a[111]), .Z(n9738) );
  NAND U20071 ( .A(a[114]), .B(b[0]), .Z(n8388) );
  XNOR U20072 ( .A(n9070), .B(n9071), .Z(c[113]) );
  XNOR U20073 ( .A(n9736), .B(n9737), .Z(n9071) );
  XOR U20074 ( .A(n9734), .B(n9743), .Z(n9737) );
  NAND U20075 ( .A(b[1]), .B(a[112]), .Z(n9743) );
  XOR U20076 ( .A(n9742), .B(n9744), .Z(n9736) );
  XOR U20077 ( .A(n9734), .B(n9741), .Z(n9744) );
  XNOR U20078 ( .A(n9745), .B(n9740), .Z(n9741) );
  AND U20079 ( .A(b[2]), .B(a[111]), .Z(n9745) );
  NANDN U20080 ( .A(n9746), .B(n9747), .Z(n9734) );
  XOR U20081 ( .A(n9740), .B(n9732), .Z(n9748) );
  XNOR U20082 ( .A(n9731), .B(n9727), .Z(n9749) );
  XNOR U20083 ( .A(n9726), .B(n9722), .Z(n9750) );
  XNOR U20084 ( .A(n9721), .B(n9717), .Z(n9751) );
  XNOR U20085 ( .A(n9716), .B(n9712), .Z(n9752) );
  XNOR U20086 ( .A(n9711), .B(n9707), .Z(n9753) );
  XNOR U20087 ( .A(n9706), .B(n9702), .Z(n9754) );
  XNOR U20088 ( .A(n9701), .B(n9697), .Z(n9755) );
  XNOR U20089 ( .A(n9696), .B(n9692), .Z(n9756) );
  XNOR U20090 ( .A(n9691), .B(n9687), .Z(n9757) );
  XNOR U20091 ( .A(n9686), .B(n9682), .Z(n9758) );
  XNOR U20092 ( .A(n9681), .B(n9677), .Z(n9759) );
  XNOR U20093 ( .A(n9676), .B(n9672), .Z(n9760) );
  XNOR U20094 ( .A(n9671), .B(n9667), .Z(n9761) );
  XNOR U20095 ( .A(n9666), .B(n9662), .Z(n9762) );
  XNOR U20096 ( .A(n9661), .B(n9657), .Z(n9763) );
  XNOR U20097 ( .A(n9656), .B(n9652), .Z(n9764) );
  XNOR U20098 ( .A(n9651), .B(n9647), .Z(n9765) );
  XNOR U20099 ( .A(n9646), .B(n9642), .Z(n9766) );
  XNOR U20100 ( .A(n9641), .B(n9637), .Z(n9767) );
  XNOR U20101 ( .A(n9636), .B(n9632), .Z(n9768) );
  XNOR U20102 ( .A(n9631), .B(n9627), .Z(n9769) );
  XNOR U20103 ( .A(n9626), .B(n9622), .Z(n9770) );
  XNOR U20104 ( .A(n9621), .B(n9617), .Z(n9771) );
  XNOR U20105 ( .A(n9616), .B(n9612), .Z(n9772) );
  XNOR U20106 ( .A(n9611), .B(n9607), .Z(n9773) );
  XNOR U20107 ( .A(n9606), .B(n9602), .Z(n9774) );
  XNOR U20108 ( .A(n9601), .B(n9597), .Z(n9775) );
  XNOR U20109 ( .A(n9596), .B(n9592), .Z(n9776) );
  XNOR U20110 ( .A(n9591), .B(n9587), .Z(n9777) );
  XNOR U20111 ( .A(n9586), .B(n9582), .Z(n9778) );
  XNOR U20112 ( .A(n9581), .B(n9577), .Z(n9779) );
  XNOR U20113 ( .A(n9576), .B(n9572), .Z(n9780) );
  XNOR U20114 ( .A(n9571), .B(n9567), .Z(n9781) );
  XNOR U20115 ( .A(n9566), .B(n9562), .Z(n9782) );
  XNOR U20116 ( .A(n9561), .B(n9557), .Z(n9783) );
  XNOR U20117 ( .A(n9556), .B(n9552), .Z(n9784) );
  XNOR U20118 ( .A(n9551), .B(n9547), .Z(n9785) );
  XNOR U20119 ( .A(n9546), .B(n9542), .Z(n9786) );
  XNOR U20120 ( .A(n9541), .B(n9537), .Z(n9787) );
  XNOR U20121 ( .A(n9536), .B(n9532), .Z(n9788) );
  XNOR U20122 ( .A(n9531), .B(n9527), .Z(n9789) );
  XNOR U20123 ( .A(n9526), .B(n9522), .Z(n9790) );
  XNOR U20124 ( .A(n9521), .B(n9517), .Z(n9791) );
  XNOR U20125 ( .A(n9516), .B(n9512), .Z(n9792) );
  XNOR U20126 ( .A(n9511), .B(n9507), .Z(n9793) );
  XNOR U20127 ( .A(n9506), .B(n9502), .Z(n9794) );
  XNOR U20128 ( .A(n9501), .B(n9497), .Z(n9795) );
  XNOR U20129 ( .A(n9496), .B(n9492), .Z(n9796) );
  XNOR U20130 ( .A(n9491), .B(n9487), .Z(n9797) );
  XNOR U20131 ( .A(n9486), .B(n9482), .Z(n9798) );
  XNOR U20132 ( .A(n9481), .B(n9477), .Z(n9799) );
  XNOR U20133 ( .A(n9476), .B(n9472), .Z(n9800) );
  XNOR U20134 ( .A(n9471), .B(n9467), .Z(n9801) );
  XNOR U20135 ( .A(n9466), .B(n9462), .Z(n9802) );
  XNOR U20136 ( .A(n9461), .B(n9457), .Z(n9803) );
  XNOR U20137 ( .A(n9456), .B(n9452), .Z(n9804) );
  XNOR U20138 ( .A(n9451), .B(n9447), .Z(n9805) );
  XNOR U20139 ( .A(n9446), .B(n9442), .Z(n9806) );
  XNOR U20140 ( .A(n9441), .B(n9437), .Z(n9807) );
  XNOR U20141 ( .A(n9436), .B(n9432), .Z(n9808) );
  XNOR U20142 ( .A(n9431), .B(n9427), .Z(n9809) );
  XNOR U20143 ( .A(n9426), .B(n9422), .Z(n9810) );
  XNOR U20144 ( .A(n9421), .B(n9417), .Z(n9811) );
  XNOR U20145 ( .A(n9416), .B(n9412), .Z(n9812) );
  XNOR U20146 ( .A(n9411), .B(n9407), .Z(n9813) );
  XNOR U20147 ( .A(n9406), .B(n9402), .Z(n9814) );
  XNOR U20148 ( .A(n9401), .B(n9397), .Z(n9815) );
  XNOR U20149 ( .A(n9396), .B(n9392), .Z(n9816) );
  XNOR U20150 ( .A(n9391), .B(n9387), .Z(n9817) );
  XNOR U20151 ( .A(n9386), .B(n9382), .Z(n9818) );
  XNOR U20152 ( .A(n9381), .B(n9377), .Z(n9819) );
  XNOR U20153 ( .A(n9376), .B(n9372), .Z(n9820) );
  XNOR U20154 ( .A(n9371), .B(n9367), .Z(n9821) );
  XNOR U20155 ( .A(n9366), .B(n9362), .Z(n9822) );
  XNOR U20156 ( .A(n9361), .B(n9357), .Z(n9823) );
  XNOR U20157 ( .A(n9356), .B(n9352), .Z(n9824) );
  XNOR U20158 ( .A(n9351), .B(n9347), .Z(n9825) );
  XNOR U20159 ( .A(n9346), .B(n9342), .Z(n9826) );
  XNOR U20160 ( .A(n9341), .B(n9337), .Z(n9827) );
  XNOR U20161 ( .A(n9336), .B(n9332), .Z(n9828) );
  XNOR U20162 ( .A(n9331), .B(n9327), .Z(n9829) );
  XNOR U20163 ( .A(n9326), .B(n9322), .Z(n9830) );
  XNOR U20164 ( .A(n9321), .B(n9317), .Z(n9831) );
  XNOR U20165 ( .A(n9316), .B(n9312), .Z(n9832) );
  XNOR U20166 ( .A(n9311), .B(n9307), .Z(n9833) );
  XNOR U20167 ( .A(n9306), .B(n9302), .Z(n9834) );
  XNOR U20168 ( .A(n9301), .B(n9297), .Z(n9835) );
  XNOR U20169 ( .A(n9296), .B(n9292), .Z(n9836) );
  XNOR U20170 ( .A(n9291), .B(n9287), .Z(n9837) );
  XNOR U20171 ( .A(n9286), .B(n9282), .Z(n9838) );
  XNOR U20172 ( .A(n9281), .B(n9277), .Z(n9839) );
  XNOR U20173 ( .A(n9276), .B(n9272), .Z(n9840) );
  XNOR U20174 ( .A(n9271), .B(n9267), .Z(n9841) );
  XNOR U20175 ( .A(n9266), .B(n9262), .Z(n9842) );
  XNOR U20176 ( .A(n9261), .B(n9257), .Z(n9843) );
  XNOR U20177 ( .A(n9256), .B(n9252), .Z(n9844) );
  XNOR U20178 ( .A(n9251), .B(n9247), .Z(n9845) );
  XNOR U20179 ( .A(n9246), .B(n9242), .Z(n9846) );
  XNOR U20180 ( .A(n9241), .B(n9237), .Z(n9847) );
  XNOR U20181 ( .A(n9236), .B(n9232), .Z(n9848) );
  XNOR U20182 ( .A(n9231), .B(n9227), .Z(n9849) );
  XNOR U20183 ( .A(n9226), .B(n9222), .Z(n9850) );
  XNOR U20184 ( .A(n9221), .B(n9217), .Z(n9851) );
  XNOR U20185 ( .A(n9216), .B(n9212), .Z(n9852) );
  XNOR U20186 ( .A(n9211), .B(n9207), .Z(n9853) );
  XNOR U20187 ( .A(n9206), .B(n9202), .Z(n9854) );
  XNOR U20188 ( .A(n9201), .B(n9197), .Z(n9855) );
  XNOR U20189 ( .A(n9196), .B(n9192), .Z(n9856) );
  XNOR U20190 ( .A(n9191), .B(n9187), .Z(n9857) );
  XNOR U20191 ( .A(n9858), .B(n9186), .Z(n9187) );
  AND U20192 ( .A(a[0]), .B(b[113]), .Z(n9858) );
  XOR U20193 ( .A(n9859), .B(n9186), .Z(n9188) );
  XNOR U20194 ( .A(n9860), .B(n9861), .Z(n9186) );
  ANDN U20195 ( .B(n9862), .A(n9863), .Z(n9860) );
  AND U20196 ( .A(a[1]), .B(b[112]), .Z(n9859) );
  XNOR U20197 ( .A(n9864), .B(n9191), .Z(n9193) );
  XOR U20198 ( .A(n9865), .B(n9866), .Z(n9191) );
  ANDN U20199 ( .B(n9867), .A(n9868), .Z(n9865) );
  AND U20200 ( .A(a[2]), .B(b[111]), .Z(n9864) );
  XNOR U20201 ( .A(n9869), .B(n9196), .Z(n9198) );
  XOR U20202 ( .A(n9870), .B(n9871), .Z(n9196) );
  ANDN U20203 ( .B(n9872), .A(n9873), .Z(n9870) );
  AND U20204 ( .A(a[3]), .B(b[110]), .Z(n9869) );
  XNOR U20205 ( .A(n9874), .B(n9201), .Z(n9203) );
  XOR U20206 ( .A(n9875), .B(n9876), .Z(n9201) );
  ANDN U20207 ( .B(n9877), .A(n9878), .Z(n9875) );
  AND U20208 ( .A(a[4]), .B(b[109]), .Z(n9874) );
  XNOR U20209 ( .A(n9879), .B(n9206), .Z(n9208) );
  XOR U20210 ( .A(n9880), .B(n9881), .Z(n9206) );
  ANDN U20211 ( .B(n9882), .A(n9883), .Z(n9880) );
  AND U20212 ( .A(a[5]), .B(b[108]), .Z(n9879) );
  XNOR U20213 ( .A(n9884), .B(n9211), .Z(n9213) );
  XOR U20214 ( .A(n9885), .B(n9886), .Z(n9211) );
  ANDN U20215 ( .B(n9887), .A(n9888), .Z(n9885) );
  AND U20216 ( .A(a[6]), .B(b[107]), .Z(n9884) );
  XNOR U20217 ( .A(n9889), .B(n9216), .Z(n9218) );
  XOR U20218 ( .A(n9890), .B(n9891), .Z(n9216) );
  ANDN U20219 ( .B(n9892), .A(n9893), .Z(n9890) );
  AND U20220 ( .A(a[7]), .B(b[106]), .Z(n9889) );
  XNOR U20221 ( .A(n9894), .B(n9221), .Z(n9223) );
  XOR U20222 ( .A(n9895), .B(n9896), .Z(n9221) );
  ANDN U20223 ( .B(n9897), .A(n9898), .Z(n9895) );
  AND U20224 ( .A(a[8]), .B(b[105]), .Z(n9894) );
  XNOR U20225 ( .A(n9899), .B(n9226), .Z(n9228) );
  XOR U20226 ( .A(n9900), .B(n9901), .Z(n9226) );
  ANDN U20227 ( .B(n9902), .A(n9903), .Z(n9900) );
  AND U20228 ( .A(a[9]), .B(b[104]), .Z(n9899) );
  XNOR U20229 ( .A(n9904), .B(n9231), .Z(n9233) );
  XOR U20230 ( .A(n9905), .B(n9906), .Z(n9231) );
  ANDN U20231 ( .B(n9907), .A(n9908), .Z(n9905) );
  AND U20232 ( .A(a[10]), .B(b[103]), .Z(n9904) );
  XNOR U20233 ( .A(n9909), .B(n9236), .Z(n9238) );
  XOR U20234 ( .A(n9910), .B(n9911), .Z(n9236) );
  ANDN U20235 ( .B(n9912), .A(n9913), .Z(n9910) );
  AND U20236 ( .A(a[11]), .B(b[102]), .Z(n9909) );
  XNOR U20237 ( .A(n9914), .B(n9241), .Z(n9243) );
  XOR U20238 ( .A(n9915), .B(n9916), .Z(n9241) );
  ANDN U20239 ( .B(n9917), .A(n9918), .Z(n9915) );
  AND U20240 ( .A(a[12]), .B(b[101]), .Z(n9914) );
  XNOR U20241 ( .A(n9919), .B(n9246), .Z(n9248) );
  XOR U20242 ( .A(n9920), .B(n9921), .Z(n9246) );
  ANDN U20243 ( .B(n9922), .A(n9923), .Z(n9920) );
  AND U20244 ( .A(a[13]), .B(b[100]), .Z(n9919) );
  XNOR U20245 ( .A(n9924), .B(n9251), .Z(n9253) );
  XOR U20246 ( .A(n9925), .B(n9926), .Z(n9251) );
  ANDN U20247 ( .B(n9927), .A(n9928), .Z(n9925) );
  AND U20248 ( .A(a[14]), .B(b[99]), .Z(n9924) );
  XNOR U20249 ( .A(n9929), .B(n9256), .Z(n9258) );
  XOR U20250 ( .A(n9930), .B(n9931), .Z(n9256) );
  ANDN U20251 ( .B(n9932), .A(n9933), .Z(n9930) );
  AND U20252 ( .A(a[15]), .B(b[98]), .Z(n9929) );
  XNOR U20253 ( .A(n9934), .B(n9261), .Z(n9263) );
  XOR U20254 ( .A(n9935), .B(n9936), .Z(n9261) );
  ANDN U20255 ( .B(n9937), .A(n9938), .Z(n9935) );
  AND U20256 ( .A(a[16]), .B(b[97]), .Z(n9934) );
  XNOR U20257 ( .A(n9939), .B(n9266), .Z(n9268) );
  XOR U20258 ( .A(n9940), .B(n9941), .Z(n9266) );
  ANDN U20259 ( .B(n9942), .A(n9943), .Z(n9940) );
  AND U20260 ( .A(a[17]), .B(b[96]), .Z(n9939) );
  XNOR U20261 ( .A(n9944), .B(n9271), .Z(n9273) );
  XOR U20262 ( .A(n9945), .B(n9946), .Z(n9271) );
  ANDN U20263 ( .B(n9947), .A(n9948), .Z(n9945) );
  AND U20264 ( .A(a[18]), .B(b[95]), .Z(n9944) );
  XNOR U20265 ( .A(n9949), .B(n9276), .Z(n9278) );
  XOR U20266 ( .A(n9950), .B(n9951), .Z(n9276) );
  ANDN U20267 ( .B(n9952), .A(n9953), .Z(n9950) );
  AND U20268 ( .A(a[19]), .B(b[94]), .Z(n9949) );
  XNOR U20269 ( .A(n9954), .B(n9281), .Z(n9283) );
  XOR U20270 ( .A(n9955), .B(n9956), .Z(n9281) );
  ANDN U20271 ( .B(n9957), .A(n9958), .Z(n9955) );
  AND U20272 ( .A(a[20]), .B(b[93]), .Z(n9954) );
  XNOR U20273 ( .A(n9959), .B(n9286), .Z(n9288) );
  XOR U20274 ( .A(n9960), .B(n9961), .Z(n9286) );
  ANDN U20275 ( .B(n9962), .A(n9963), .Z(n9960) );
  AND U20276 ( .A(a[21]), .B(b[92]), .Z(n9959) );
  XNOR U20277 ( .A(n9964), .B(n9291), .Z(n9293) );
  XOR U20278 ( .A(n9965), .B(n9966), .Z(n9291) );
  ANDN U20279 ( .B(n9967), .A(n9968), .Z(n9965) );
  AND U20280 ( .A(a[22]), .B(b[91]), .Z(n9964) );
  XNOR U20281 ( .A(n9969), .B(n9296), .Z(n9298) );
  XOR U20282 ( .A(n9970), .B(n9971), .Z(n9296) );
  ANDN U20283 ( .B(n9972), .A(n9973), .Z(n9970) );
  AND U20284 ( .A(a[23]), .B(b[90]), .Z(n9969) );
  XNOR U20285 ( .A(n9974), .B(n9301), .Z(n9303) );
  XOR U20286 ( .A(n9975), .B(n9976), .Z(n9301) );
  ANDN U20287 ( .B(n9977), .A(n9978), .Z(n9975) );
  AND U20288 ( .A(a[24]), .B(b[89]), .Z(n9974) );
  XNOR U20289 ( .A(n9979), .B(n9306), .Z(n9308) );
  XOR U20290 ( .A(n9980), .B(n9981), .Z(n9306) );
  ANDN U20291 ( .B(n9982), .A(n9983), .Z(n9980) );
  AND U20292 ( .A(a[25]), .B(b[88]), .Z(n9979) );
  XNOR U20293 ( .A(n9984), .B(n9311), .Z(n9313) );
  XOR U20294 ( .A(n9985), .B(n9986), .Z(n9311) );
  ANDN U20295 ( .B(n9987), .A(n9988), .Z(n9985) );
  AND U20296 ( .A(a[26]), .B(b[87]), .Z(n9984) );
  XNOR U20297 ( .A(n9989), .B(n9316), .Z(n9318) );
  XOR U20298 ( .A(n9990), .B(n9991), .Z(n9316) );
  ANDN U20299 ( .B(n9992), .A(n9993), .Z(n9990) );
  AND U20300 ( .A(a[27]), .B(b[86]), .Z(n9989) );
  XNOR U20301 ( .A(n9994), .B(n9321), .Z(n9323) );
  XOR U20302 ( .A(n9995), .B(n9996), .Z(n9321) );
  ANDN U20303 ( .B(n9997), .A(n9998), .Z(n9995) );
  AND U20304 ( .A(a[28]), .B(b[85]), .Z(n9994) );
  XNOR U20305 ( .A(n9999), .B(n9326), .Z(n9328) );
  XOR U20306 ( .A(n10000), .B(n10001), .Z(n9326) );
  ANDN U20307 ( .B(n10002), .A(n10003), .Z(n10000) );
  AND U20308 ( .A(a[29]), .B(b[84]), .Z(n9999) );
  XNOR U20309 ( .A(n10004), .B(n9331), .Z(n9333) );
  XOR U20310 ( .A(n10005), .B(n10006), .Z(n9331) );
  ANDN U20311 ( .B(n10007), .A(n10008), .Z(n10005) );
  AND U20312 ( .A(a[30]), .B(b[83]), .Z(n10004) );
  XNOR U20313 ( .A(n10009), .B(n9336), .Z(n9338) );
  XOR U20314 ( .A(n10010), .B(n10011), .Z(n9336) );
  ANDN U20315 ( .B(n10012), .A(n10013), .Z(n10010) );
  AND U20316 ( .A(a[31]), .B(b[82]), .Z(n10009) );
  XNOR U20317 ( .A(n10014), .B(n9341), .Z(n9343) );
  XOR U20318 ( .A(n10015), .B(n10016), .Z(n9341) );
  ANDN U20319 ( .B(n10017), .A(n10018), .Z(n10015) );
  AND U20320 ( .A(a[32]), .B(b[81]), .Z(n10014) );
  XNOR U20321 ( .A(n10019), .B(n9346), .Z(n9348) );
  XOR U20322 ( .A(n10020), .B(n10021), .Z(n9346) );
  ANDN U20323 ( .B(n10022), .A(n10023), .Z(n10020) );
  AND U20324 ( .A(a[33]), .B(b[80]), .Z(n10019) );
  XNOR U20325 ( .A(n10024), .B(n9351), .Z(n9353) );
  XOR U20326 ( .A(n10025), .B(n10026), .Z(n9351) );
  ANDN U20327 ( .B(n10027), .A(n10028), .Z(n10025) );
  AND U20328 ( .A(a[34]), .B(b[79]), .Z(n10024) );
  XNOR U20329 ( .A(n10029), .B(n9356), .Z(n9358) );
  XOR U20330 ( .A(n10030), .B(n10031), .Z(n9356) );
  ANDN U20331 ( .B(n10032), .A(n10033), .Z(n10030) );
  AND U20332 ( .A(a[35]), .B(b[78]), .Z(n10029) );
  XNOR U20333 ( .A(n10034), .B(n9361), .Z(n9363) );
  XOR U20334 ( .A(n10035), .B(n10036), .Z(n9361) );
  ANDN U20335 ( .B(n10037), .A(n10038), .Z(n10035) );
  AND U20336 ( .A(a[36]), .B(b[77]), .Z(n10034) );
  XNOR U20337 ( .A(n10039), .B(n9366), .Z(n9368) );
  XOR U20338 ( .A(n10040), .B(n10041), .Z(n9366) );
  ANDN U20339 ( .B(n10042), .A(n10043), .Z(n10040) );
  AND U20340 ( .A(a[37]), .B(b[76]), .Z(n10039) );
  XNOR U20341 ( .A(n10044), .B(n9371), .Z(n9373) );
  XOR U20342 ( .A(n10045), .B(n10046), .Z(n9371) );
  ANDN U20343 ( .B(n10047), .A(n10048), .Z(n10045) );
  AND U20344 ( .A(a[38]), .B(b[75]), .Z(n10044) );
  XNOR U20345 ( .A(n10049), .B(n9376), .Z(n9378) );
  XOR U20346 ( .A(n10050), .B(n10051), .Z(n9376) );
  ANDN U20347 ( .B(n10052), .A(n10053), .Z(n10050) );
  AND U20348 ( .A(a[39]), .B(b[74]), .Z(n10049) );
  XNOR U20349 ( .A(n10054), .B(n9381), .Z(n9383) );
  XOR U20350 ( .A(n10055), .B(n10056), .Z(n9381) );
  ANDN U20351 ( .B(n10057), .A(n10058), .Z(n10055) );
  AND U20352 ( .A(a[40]), .B(b[73]), .Z(n10054) );
  XNOR U20353 ( .A(n10059), .B(n9386), .Z(n9388) );
  XOR U20354 ( .A(n10060), .B(n10061), .Z(n9386) );
  ANDN U20355 ( .B(n10062), .A(n10063), .Z(n10060) );
  AND U20356 ( .A(a[41]), .B(b[72]), .Z(n10059) );
  XNOR U20357 ( .A(n10064), .B(n9391), .Z(n9393) );
  XOR U20358 ( .A(n10065), .B(n10066), .Z(n9391) );
  ANDN U20359 ( .B(n10067), .A(n10068), .Z(n10065) );
  AND U20360 ( .A(a[42]), .B(b[71]), .Z(n10064) );
  XNOR U20361 ( .A(n10069), .B(n9396), .Z(n9398) );
  XOR U20362 ( .A(n10070), .B(n10071), .Z(n9396) );
  ANDN U20363 ( .B(n10072), .A(n10073), .Z(n10070) );
  AND U20364 ( .A(a[43]), .B(b[70]), .Z(n10069) );
  XNOR U20365 ( .A(n10074), .B(n9401), .Z(n9403) );
  XOR U20366 ( .A(n10075), .B(n10076), .Z(n9401) );
  ANDN U20367 ( .B(n10077), .A(n10078), .Z(n10075) );
  AND U20368 ( .A(a[44]), .B(b[69]), .Z(n10074) );
  XNOR U20369 ( .A(n10079), .B(n9406), .Z(n9408) );
  XOR U20370 ( .A(n10080), .B(n10081), .Z(n9406) );
  ANDN U20371 ( .B(n10082), .A(n10083), .Z(n10080) );
  AND U20372 ( .A(a[45]), .B(b[68]), .Z(n10079) );
  XNOR U20373 ( .A(n10084), .B(n9411), .Z(n9413) );
  XOR U20374 ( .A(n10085), .B(n10086), .Z(n9411) );
  ANDN U20375 ( .B(n10087), .A(n10088), .Z(n10085) );
  AND U20376 ( .A(a[46]), .B(b[67]), .Z(n10084) );
  XNOR U20377 ( .A(n10089), .B(n9416), .Z(n9418) );
  XOR U20378 ( .A(n10090), .B(n10091), .Z(n9416) );
  ANDN U20379 ( .B(n10092), .A(n10093), .Z(n10090) );
  AND U20380 ( .A(a[47]), .B(b[66]), .Z(n10089) );
  XNOR U20381 ( .A(n10094), .B(n9421), .Z(n9423) );
  XOR U20382 ( .A(n10095), .B(n10096), .Z(n9421) );
  ANDN U20383 ( .B(n10097), .A(n10098), .Z(n10095) );
  AND U20384 ( .A(a[48]), .B(b[65]), .Z(n10094) );
  XNOR U20385 ( .A(n10099), .B(n9426), .Z(n9428) );
  XOR U20386 ( .A(n10100), .B(n10101), .Z(n9426) );
  ANDN U20387 ( .B(n10102), .A(n10103), .Z(n10100) );
  AND U20388 ( .A(a[49]), .B(b[64]), .Z(n10099) );
  XNOR U20389 ( .A(n10104), .B(n9431), .Z(n9433) );
  XOR U20390 ( .A(n10105), .B(n10106), .Z(n9431) );
  ANDN U20391 ( .B(n10107), .A(n10108), .Z(n10105) );
  AND U20392 ( .A(a[50]), .B(b[63]), .Z(n10104) );
  XNOR U20393 ( .A(n10109), .B(n9436), .Z(n9438) );
  XOR U20394 ( .A(n10110), .B(n10111), .Z(n9436) );
  ANDN U20395 ( .B(n10112), .A(n10113), .Z(n10110) );
  AND U20396 ( .A(a[51]), .B(b[62]), .Z(n10109) );
  XNOR U20397 ( .A(n10114), .B(n9441), .Z(n9443) );
  XOR U20398 ( .A(n10115), .B(n10116), .Z(n9441) );
  ANDN U20399 ( .B(n10117), .A(n10118), .Z(n10115) );
  AND U20400 ( .A(a[52]), .B(b[61]), .Z(n10114) );
  XNOR U20401 ( .A(n10119), .B(n9446), .Z(n9448) );
  XOR U20402 ( .A(n10120), .B(n10121), .Z(n9446) );
  ANDN U20403 ( .B(n10122), .A(n10123), .Z(n10120) );
  AND U20404 ( .A(a[53]), .B(b[60]), .Z(n10119) );
  XNOR U20405 ( .A(n10124), .B(n9451), .Z(n9453) );
  XOR U20406 ( .A(n10125), .B(n10126), .Z(n9451) );
  ANDN U20407 ( .B(n10127), .A(n10128), .Z(n10125) );
  AND U20408 ( .A(a[54]), .B(b[59]), .Z(n10124) );
  XNOR U20409 ( .A(n10129), .B(n9456), .Z(n9458) );
  XOR U20410 ( .A(n10130), .B(n10131), .Z(n9456) );
  ANDN U20411 ( .B(n10132), .A(n10133), .Z(n10130) );
  AND U20412 ( .A(a[55]), .B(b[58]), .Z(n10129) );
  XNOR U20413 ( .A(n10134), .B(n9461), .Z(n9463) );
  XOR U20414 ( .A(n10135), .B(n10136), .Z(n9461) );
  ANDN U20415 ( .B(n10137), .A(n10138), .Z(n10135) );
  AND U20416 ( .A(a[56]), .B(b[57]), .Z(n10134) );
  XNOR U20417 ( .A(n10139), .B(n9466), .Z(n9468) );
  XOR U20418 ( .A(n10140), .B(n10141), .Z(n9466) );
  ANDN U20419 ( .B(n10142), .A(n10143), .Z(n10140) );
  AND U20420 ( .A(a[57]), .B(b[56]), .Z(n10139) );
  XNOR U20421 ( .A(n10144), .B(n9471), .Z(n9473) );
  XOR U20422 ( .A(n10145), .B(n10146), .Z(n9471) );
  ANDN U20423 ( .B(n10147), .A(n10148), .Z(n10145) );
  AND U20424 ( .A(a[58]), .B(b[55]), .Z(n10144) );
  XNOR U20425 ( .A(n10149), .B(n9476), .Z(n9478) );
  XOR U20426 ( .A(n10150), .B(n10151), .Z(n9476) );
  ANDN U20427 ( .B(n10152), .A(n10153), .Z(n10150) );
  AND U20428 ( .A(a[59]), .B(b[54]), .Z(n10149) );
  XNOR U20429 ( .A(n10154), .B(n9481), .Z(n9483) );
  XOR U20430 ( .A(n10155), .B(n10156), .Z(n9481) );
  ANDN U20431 ( .B(n10157), .A(n10158), .Z(n10155) );
  AND U20432 ( .A(a[60]), .B(b[53]), .Z(n10154) );
  XNOR U20433 ( .A(n10159), .B(n9486), .Z(n9488) );
  XOR U20434 ( .A(n10160), .B(n10161), .Z(n9486) );
  ANDN U20435 ( .B(n10162), .A(n10163), .Z(n10160) );
  AND U20436 ( .A(a[61]), .B(b[52]), .Z(n10159) );
  XNOR U20437 ( .A(n10164), .B(n9491), .Z(n9493) );
  XOR U20438 ( .A(n10165), .B(n10166), .Z(n9491) );
  ANDN U20439 ( .B(n10167), .A(n10168), .Z(n10165) );
  AND U20440 ( .A(a[62]), .B(b[51]), .Z(n10164) );
  XNOR U20441 ( .A(n10169), .B(n9496), .Z(n9498) );
  XOR U20442 ( .A(n10170), .B(n10171), .Z(n9496) );
  ANDN U20443 ( .B(n10172), .A(n10173), .Z(n10170) );
  AND U20444 ( .A(a[63]), .B(b[50]), .Z(n10169) );
  XNOR U20445 ( .A(n10174), .B(n9501), .Z(n9503) );
  XOR U20446 ( .A(n10175), .B(n10176), .Z(n9501) );
  ANDN U20447 ( .B(n10177), .A(n10178), .Z(n10175) );
  AND U20448 ( .A(a[64]), .B(b[49]), .Z(n10174) );
  XNOR U20449 ( .A(n10179), .B(n9506), .Z(n9508) );
  XOR U20450 ( .A(n10180), .B(n10181), .Z(n9506) );
  ANDN U20451 ( .B(n10182), .A(n10183), .Z(n10180) );
  AND U20452 ( .A(a[65]), .B(b[48]), .Z(n10179) );
  XNOR U20453 ( .A(n10184), .B(n9511), .Z(n9513) );
  XOR U20454 ( .A(n10185), .B(n10186), .Z(n9511) );
  ANDN U20455 ( .B(n10187), .A(n10188), .Z(n10185) );
  AND U20456 ( .A(a[66]), .B(b[47]), .Z(n10184) );
  XNOR U20457 ( .A(n10189), .B(n9516), .Z(n9518) );
  XOR U20458 ( .A(n10190), .B(n10191), .Z(n9516) );
  ANDN U20459 ( .B(n10192), .A(n10193), .Z(n10190) );
  AND U20460 ( .A(a[67]), .B(b[46]), .Z(n10189) );
  XNOR U20461 ( .A(n10194), .B(n9521), .Z(n9523) );
  XOR U20462 ( .A(n10195), .B(n10196), .Z(n9521) );
  ANDN U20463 ( .B(n10197), .A(n10198), .Z(n10195) );
  AND U20464 ( .A(a[68]), .B(b[45]), .Z(n10194) );
  XNOR U20465 ( .A(n10199), .B(n9526), .Z(n9528) );
  XOR U20466 ( .A(n10200), .B(n10201), .Z(n9526) );
  ANDN U20467 ( .B(n10202), .A(n10203), .Z(n10200) );
  AND U20468 ( .A(a[69]), .B(b[44]), .Z(n10199) );
  XNOR U20469 ( .A(n10204), .B(n9531), .Z(n9533) );
  XOR U20470 ( .A(n10205), .B(n10206), .Z(n9531) );
  ANDN U20471 ( .B(n10207), .A(n10208), .Z(n10205) );
  AND U20472 ( .A(a[70]), .B(b[43]), .Z(n10204) );
  XNOR U20473 ( .A(n10209), .B(n9536), .Z(n9538) );
  XOR U20474 ( .A(n10210), .B(n10211), .Z(n9536) );
  ANDN U20475 ( .B(n10212), .A(n10213), .Z(n10210) );
  AND U20476 ( .A(a[71]), .B(b[42]), .Z(n10209) );
  XNOR U20477 ( .A(n10214), .B(n9541), .Z(n9543) );
  XOR U20478 ( .A(n10215), .B(n10216), .Z(n9541) );
  ANDN U20479 ( .B(n10217), .A(n10218), .Z(n10215) );
  AND U20480 ( .A(a[72]), .B(b[41]), .Z(n10214) );
  XNOR U20481 ( .A(n10219), .B(n9546), .Z(n9548) );
  XOR U20482 ( .A(n10220), .B(n10221), .Z(n9546) );
  ANDN U20483 ( .B(n10222), .A(n10223), .Z(n10220) );
  AND U20484 ( .A(a[73]), .B(b[40]), .Z(n10219) );
  XNOR U20485 ( .A(n10224), .B(n9551), .Z(n9553) );
  XOR U20486 ( .A(n10225), .B(n10226), .Z(n9551) );
  ANDN U20487 ( .B(n10227), .A(n10228), .Z(n10225) );
  AND U20488 ( .A(a[74]), .B(b[39]), .Z(n10224) );
  XNOR U20489 ( .A(n10229), .B(n9556), .Z(n9558) );
  XOR U20490 ( .A(n10230), .B(n10231), .Z(n9556) );
  ANDN U20491 ( .B(n10232), .A(n10233), .Z(n10230) );
  AND U20492 ( .A(a[75]), .B(b[38]), .Z(n10229) );
  XNOR U20493 ( .A(n10234), .B(n9561), .Z(n9563) );
  XOR U20494 ( .A(n10235), .B(n10236), .Z(n9561) );
  ANDN U20495 ( .B(n10237), .A(n10238), .Z(n10235) );
  AND U20496 ( .A(a[76]), .B(b[37]), .Z(n10234) );
  XNOR U20497 ( .A(n10239), .B(n9566), .Z(n9568) );
  XOR U20498 ( .A(n10240), .B(n10241), .Z(n9566) );
  ANDN U20499 ( .B(n10242), .A(n10243), .Z(n10240) );
  AND U20500 ( .A(a[77]), .B(b[36]), .Z(n10239) );
  XNOR U20501 ( .A(n10244), .B(n9571), .Z(n9573) );
  XOR U20502 ( .A(n10245), .B(n10246), .Z(n9571) );
  ANDN U20503 ( .B(n10247), .A(n10248), .Z(n10245) );
  AND U20504 ( .A(a[78]), .B(b[35]), .Z(n10244) );
  XNOR U20505 ( .A(n10249), .B(n9576), .Z(n9578) );
  XOR U20506 ( .A(n10250), .B(n10251), .Z(n9576) );
  ANDN U20507 ( .B(n10252), .A(n10253), .Z(n10250) );
  AND U20508 ( .A(a[79]), .B(b[34]), .Z(n10249) );
  XNOR U20509 ( .A(n10254), .B(n9581), .Z(n9583) );
  XOR U20510 ( .A(n10255), .B(n10256), .Z(n9581) );
  ANDN U20511 ( .B(n10257), .A(n10258), .Z(n10255) );
  AND U20512 ( .A(a[80]), .B(b[33]), .Z(n10254) );
  XNOR U20513 ( .A(n10259), .B(n9586), .Z(n9588) );
  XOR U20514 ( .A(n10260), .B(n10261), .Z(n9586) );
  ANDN U20515 ( .B(n10262), .A(n10263), .Z(n10260) );
  AND U20516 ( .A(a[81]), .B(b[32]), .Z(n10259) );
  XNOR U20517 ( .A(n10264), .B(n9591), .Z(n9593) );
  XOR U20518 ( .A(n10265), .B(n10266), .Z(n9591) );
  ANDN U20519 ( .B(n10267), .A(n10268), .Z(n10265) );
  AND U20520 ( .A(a[82]), .B(b[31]), .Z(n10264) );
  XNOR U20521 ( .A(n10269), .B(n9596), .Z(n9598) );
  XOR U20522 ( .A(n10270), .B(n10271), .Z(n9596) );
  ANDN U20523 ( .B(n10272), .A(n10273), .Z(n10270) );
  AND U20524 ( .A(a[83]), .B(b[30]), .Z(n10269) );
  XNOR U20525 ( .A(n10274), .B(n9601), .Z(n9603) );
  XOR U20526 ( .A(n10275), .B(n10276), .Z(n9601) );
  ANDN U20527 ( .B(n10277), .A(n10278), .Z(n10275) );
  AND U20528 ( .A(a[84]), .B(b[29]), .Z(n10274) );
  XNOR U20529 ( .A(n10279), .B(n9606), .Z(n9608) );
  XOR U20530 ( .A(n10280), .B(n10281), .Z(n9606) );
  ANDN U20531 ( .B(n10282), .A(n10283), .Z(n10280) );
  AND U20532 ( .A(a[85]), .B(b[28]), .Z(n10279) );
  XNOR U20533 ( .A(n10284), .B(n9611), .Z(n9613) );
  XOR U20534 ( .A(n10285), .B(n10286), .Z(n9611) );
  ANDN U20535 ( .B(n10287), .A(n10288), .Z(n10285) );
  AND U20536 ( .A(a[86]), .B(b[27]), .Z(n10284) );
  XNOR U20537 ( .A(n10289), .B(n9616), .Z(n9618) );
  XOR U20538 ( .A(n10290), .B(n10291), .Z(n9616) );
  ANDN U20539 ( .B(n10292), .A(n10293), .Z(n10290) );
  AND U20540 ( .A(a[87]), .B(b[26]), .Z(n10289) );
  XNOR U20541 ( .A(n10294), .B(n9621), .Z(n9623) );
  XOR U20542 ( .A(n10295), .B(n10296), .Z(n9621) );
  ANDN U20543 ( .B(n10297), .A(n10298), .Z(n10295) );
  AND U20544 ( .A(a[88]), .B(b[25]), .Z(n10294) );
  XNOR U20545 ( .A(n10299), .B(n9626), .Z(n9628) );
  XOR U20546 ( .A(n10300), .B(n10301), .Z(n9626) );
  ANDN U20547 ( .B(n10302), .A(n10303), .Z(n10300) );
  AND U20548 ( .A(a[89]), .B(b[24]), .Z(n10299) );
  XNOR U20549 ( .A(n10304), .B(n9631), .Z(n9633) );
  XOR U20550 ( .A(n10305), .B(n10306), .Z(n9631) );
  ANDN U20551 ( .B(n10307), .A(n10308), .Z(n10305) );
  AND U20552 ( .A(a[90]), .B(b[23]), .Z(n10304) );
  XNOR U20553 ( .A(n10309), .B(n9636), .Z(n9638) );
  XOR U20554 ( .A(n10310), .B(n10311), .Z(n9636) );
  ANDN U20555 ( .B(n10312), .A(n10313), .Z(n10310) );
  AND U20556 ( .A(a[91]), .B(b[22]), .Z(n10309) );
  XNOR U20557 ( .A(n10314), .B(n9641), .Z(n9643) );
  XOR U20558 ( .A(n10315), .B(n10316), .Z(n9641) );
  ANDN U20559 ( .B(n10317), .A(n10318), .Z(n10315) );
  AND U20560 ( .A(a[92]), .B(b[21]), .Z(n10314) );
  XNOR U20561 ( .A(n10319), .B(n9646), .Z(n9648) );
  XOR U20562 ( .A(n10320), .B(n10321), .Z(n9646) );
  ANDN U20563 ( .B(n10322), .A(n10323), .Z(n10320) );
  AND U20564 ( .A(a[93]), .B(b[20]), .Z(n10319) );
  XNOR U20565 ( .A(n10324), .B(n9651), .Z(n9653) );
  XOR U20566 ( .A(n10325), .B(n10326), .Z(n9651) );
  ANDN U20567 ( .B(n10327), .A(n10328), .Z(n10325) );
  AND U20568 ( .A(a[94]), .B(b[19]), .Z(n10324) );
  XNOR U20569 ( .A(n10329), .B(n9656), .Z(n9658) );
  XOR U20570 ( .A(n10330), .B(n10331), .Z(n9656) );
  ANDN U20571 ( .B(n10332), .A(n10333), .Z(n10330) );
  AND U20572 ( .A(a[95]), .B(b[18]), .Z(n10329) );
  XNOR U20573 ( .A(n10334), .B(n9661), .Z(n9663) );
  XOR U20574 ( .A(n10335), .B(n10336), .Z(n9661) );
  ANDN U20575 ( .B(n10337), .A(n10338), .Z(n10335) );
  AND U20576 ( .A(a[96]), .B(b[17]), .Z(n10334) );
  XNOR U20577 ( .A(n10339), .B(n9666), .Z(n9668) );
  XOR U20578 ( .A(n10340), .B(n10341), .Z(n9666) );
  ANDN U20579 ( .B(n10342), .A(n10343), .Z(n10340) );
  AND U20580 ( .A(a[97]), .B(b[16]), .Z(n10339) );
  XNOR U20581 ( .A(n10344), .B(n9671), .Z(n9673) );
  XOR U20582 ( .A(n10345), .B(n10346), .Z(n9671) );
  ANDN U20583 ( .B(n10347), .A(n10348), .Z(n10345) );
  AND U20584 ( .A(a[98]), .B(b[15]), .Z(n10344) );
  XNOR U20585 ( .A(n10349), .B(n9676), .Z(n9678) );
  XOR U20586 ( .A(n10350), .B(n10351), .Z(n9676) );
  ANDN U20587 ( .B(n10352), .A(n10353), .Z(n10350) );
  AND U20588 ( .A(a[99]), .B(b[14]), .Z(n10349) );
  XNOR U20589 ( .A(n10354), .B(n9681), .Z(n9683) );
  XOR U20590 ( .A(n10355), .B(n10356), .Z(n9681) );
  ANDN U20591 ( .B(n10357), .A(n10358), .Z(n10355) );
  AND U20592 ( .A(b[13]), .B(a[100]), .Z(n10354) );
  XNOR U20593 ( .A(n10359), .B(n9686), .Z(n9688) );
  XOR U20594 ( .A(n10360), .B(n10361), .Z(n9686) );
  ANDN U20595 ( .B(n10362), .A(n10363), .Z(n10360) );
  AND U20596 ( .A(b[12]), .B(a[101]), .Z(n10359) );
  XNOR U20597 ( .A(n10364), .B(n9691), .Z(n9693) );
  XOR U20598 ( .A(n10365), .B(n10366), .Z(n9691) );
  ANDN U20599 ( .B(n10367), .A(n10368), .Z(n10365) );
  AND U20600 ( .A(b[11]), .B(a[102]), .Z(n10364) );
  XNOR U20601 ( .A(n10369), .B(n9696), .Z(n9698) );
  XOR U20602 ( .A(n10370), .B(n10371), .Z(n9696) );
  ANDN U20603 ( .B(n10372), .A(n10373), .Z(n10370) );
  AND U20604 ( .A(b[10]), .B(a[103]), .Z(n10369) );
  XNOR U20605 ( .A(n10374), .B(n9701), .Z(n9703) );
  XOR U20606 ( .A(n10375), .B(n10376), .Z(n9701) );
  ANDN U20607 ( .B(n10377), .A(n10378), .Z(n10375) );
  AND U20608 ( .A(b[9]), .B(a[104]), .Z(n10374) );
  XNOR U20609 ( .A(n10379), .B(n9706), .Z(n9708) );
  XOR U20610 ( .A(n10380), .B(n10381), .Z(n9706) );
  ANDN U20611 ( .B(n10382), .A(n10383), .Z(n10380) );
  AND U20612 ( .A(b[8]), .B(a[105]), .Z(n10379) );
  XNOR U20613 ( .A(n10384), .B(n9711), .Z(n9713) );
  XOR U20614 ( .A(n10385), .B(n10386), .Z(n9711) );
  ANDN U20615 ( .B(n10387), .A(n10388), .Z(n10385) );
  AND U20616 ( .A(b[7]), .B(a[106]), .Z(n10384) );
  XNOR U20617 ( .A(n10389), .B(n9716), .Z(n9718) );
  XOR U20618 ( .A(n10390), .B(n10391), .Z(n9716) );
  ANDN U20619 ( .B(n10392), .A(n10393), .Z(n10390) );
  AND U20620 ( .A(b[6]), .B(a[107]), .Z(n10389) );
  XNOR U20621 ( .A(n10394), .B(n9721), .Z(n9723) );
  XOR U20622 ( .A(n10395), .B(n10396), .Z(n9721) );
  ANDN U20623 ( .B(n10397), .A(n10398), .Z(n10395) );
  AND U20624 ( .A(b[5]), .B(a[108]), .Z(n10394) );
  XNOR U20625 ( .A(n10399), .B(n9726), .Z(n9728) );
  XOR U20626 ( .A(n10400), .B(n10401), .Z(n9726) );
  ANDN U20627 ( .B(n10402), .A(n10403), .Z(n10400) );
  AND U20628 ( .A(b[4]), .B(a[109]), .Z(n10399) );
  XNOR U20629 ( .A(n10404), .B(n10405), .Z(n9740) );
  NANDN U20630 ( .A(n10406), .B(n10407), .Z(n10405) );
  XNOR U20631 ( .A(n10408), .B(n9731), .Z(n9733) );
  XNOR U20632 ( .A(n10409), .B(n10410), .Z(n9731) );
  AND U20633 ( .A(n10411), .B(n10412), .Z(n10409) );
  AND U20634 ( .A(b[3]), .B(a[110]), .Z(n10408) );
  NAND U20635 ( .A(a[113]), .B(b[0]), .Z(n9070) );
  XNOR U20636 ( .A(n9746), .B(n9747), .Z(c[112]) );
  XNOR U20637 ( .A(n10406), .B(n10407), .Z(n9747) );
  XOR U20638 ( .A(n10404), .B(n10413), .Z(n10407) );
  NAND U20639 ( .A(b[1]), .B(a[111]), .Z(n10413) );
  XOR U20640 ( .A(n10412), .B(n10414), .Z(n10406) );
  XOR U20641 ( .A(n10404), .B(n10411), .Z(n10414) );
  XNOR U20642 ( .A(n10415), .B(n10410), .Z(n10411) );
  AND U20643 ( .A(b[2]), .B(a[110]), .Z(n10415) );
  NANDN U20644 ( .A(n10416), .B(n10417), .Z(n10404) );
  XOR U20645 ( .A(n10410), .B(n10402), .Z(n10418) );
  XNOR U20646 ( .A(n10401), .B(n10397), .Z(n10419) );
  XNOR U20647 ( .A(n10396), .B(n10392), .Z(n10420) );
  XNOR U20648 ( .A(n10391), .B(n10387), .Z(n10421) );
  XNOR U20649 ( .A(n10386), .B(n10382), .Z(n10422) );
  XNOR U20650 ( .A(n10381), .B(n10377), .Z(n10423) );
  XNOR U20651 ( .A(n10376), .B(n10372), .Z(n10424) );
  XNOR U20652 ( .A(n10371), .B(n10367), .Z(n10425) );
  XNOR U20653 ( .A(n10366), .B(n10362), .Z(n10426) );
  XNOR U20654 ( .A(n10361), .B(n10357), .Z(n10427) );
  XNOR U20655 ( .A(n10356), .B(n10352), .Z(n10428) );
  XNOR U20656 ( .A(n10351), .B(n10347), .Z(n10429) );
  XNOR U20657 ( .A(n10346), .B(n10342), .Z(n10430) );
  XNOR U20658 ( .A(n10341), .B(n10337), .Z(n10431) );
  XNOR U20659 ( .A(n10336), .B(n10332), .Z(n10432) );
  XNOR U20660 ( .A(n10331), .B(n10327), .Z(n10433) );
  XNOR U20661 ( .A(n10326), .B(n10322), .Z(n10434) );
  XNOR U20662 ( .A(n10321), .B(n10317), .Z(n10435) );
  XNOR U20663 ( .A(n10316), .B(n10312), .Z(n10436) );
  XNOR U20664 ( .A(n10311), .B(n10307), .Z(n10437) );
  XNOR U20665 ( .A(n10306), .B(n10302), .Z(n10438) );
  XNOR U20666 ( .A(n10301), .B(n10297), .Z(n10439) );
  XNOR U20667 ( .A(n10296), .B(n10292), .Z(n10440) );
  XNOR U20668 ( .A(n10291), .B(n10287), .Z(n10441) );
  XNOR U20669 ( .A(n10286), .B(n10282), .Z(n10442) );
  XNOR U20670 ( .A(n10281), .B(n10277), .Z(n10443) );
  XNOR U20671 ( .A(n10276), .B(n10272), .Z(n10444) );
  XNOR U20672 ( .A(n10271), .B(n10267), .Z(n10445) );
  XNOR U20673 ( .A(n10266), .B(n10262), .Z(n10446) );
  XNOR U20674 ( .A(n10261), .B(n10257), .Z(n10447) );
  XNOR U20675 ( .A(n10256), .B(n10252), .Z(n10448) );
  XNOR U20676 ( .A(n10251), .B(n10247), .Z(n10449) );
  XNOR U20677 ( .A(n10246), .B(n10242), .Z(n10450) );
  XNOR U20678 ( .A(n10241), .B(n10237), .Z(n10451) );
  XNOR U20679 ( .A(n10236), .B(n10232), .Z(n10452) );
  XNOR U20680 ( .A(n10231), .B(n10227), .Z(n10453) );
  XNOR U20681 ( .A(n10226), .B(n10222), .Z(n10454) );
  XNOR U20682 ( .A(n10221), .B(n10217), .Z(n10455) );
  XNOR U20683 ( .A(n10216), .B(n10212), .Z(n10456) );
  XNOR U20684 ( .A(n10211), .B(n10207), .Z(n10457) );
  XNOR U20685 ( .A(n10206), .B(n10202), .Z(n10458) );
  XNOR U20686 ( .A(n10201), .B(n10197), .Z(n10459) );
  XNOR U20687 ( .A(n10196), .B(n10192), .Z(n10460) );
  XNOR U20688 ( .A(n10191), .B(n10187), .Z(n10461) );
  XNOR U20689 ( .A(n10186), .B(n10182), .Z(n10462) );
  XNOR U20690 ( .A(n10181), .B(n10177), .Z(n10463) );
  XNOR U20691 ( .A(n10176), .B(n10172), .Z(n10464) );
  XNOR U20692 ( .A(n10171), .B(n10167), .Z(n10465) );
  XNOR U20693 ( .A(n10166), .B(n10162), .Z(n10466) );
  XNOR U20694 ( .A(n10161), .B(n10157), .Z(n10467) );
  XNOR U20695 ( .A(n10156), .B(n10152), .Z(n10468) );
  XNOR U20696 ( .A(n10151), .B(n10147), .Z(n10469) );
  XNOR U20697 ( .A(n10146), .B(n10142), .Z(n10470) );
  XNOR U20698 ( .A(n10141), .B(n10137), .Z(n10471) );
  XNOR U20699 ( .A(n10136), .B(n10132), .Z(n10472) );
  XNOR U20700 ( .A(n10131), .B(n10127), .Z(n10473) );
  XNOR U20701 ( .A(n10126), .B(n10122), .Z(n10474) );
  XNOR U20702 ( .A(n10121), .B(n10117), .Z(n10475) );
  XNOR U20703 ( .A(n10116), .B(n10112), .Z(n10476) );
  XNOR U20704 ( .A(n10111), .B(n10107), .Z(n10477) );
  XNOR U20705 ( .A(n10106), .B(n10102), .Z(n10478) );
  XNOR U20706 ( .A(n10101), .B(n10097), .Z(n10479) );
  XNOR U20707 ( .A(n10096), .B(n10092), .Z(n10480) );
  XNOR U20708 ( .A(n10091), .B(n10087), .Z(n10481) );
  XNOR U20709 ( .A(n10086), .B(n10082), .Z(n10482) );
  XNOR U20710 ( .A(n10081), .B(n10077), .Z(n10483) );
  XNOR U20711 ( .A(n10076), .B(n10072), .Z(n10484) );
  XNOR U20712 ( .A(n10071), .B(n10067), .Z(n10485) );
  XNOR U20713 ( .A(n10066), .B(n10062), .Z(n10486) );
  XNOR U20714 ( .A(n10061), .B(n10057), .Z(n10487) );
  XNOR U20715 ( .A(n10056), .B(n10052), .Z(n10488) );
  XNOR U20716 ( .A(n10051), .B(n10047), .Z(n10489) );
  XNOR U20717 ( .A(n10046), .B(n10042), .Z(n10490) );
  XNOR U20718 ( .A(n10041), .B(n10037), .Z(n10491) );
  XNOR U20719 ( .A(n10036), .B(n10032), .Z(n10492) );
  XNOR U20720 ( .A(n10031), .B(n10027), .Z(n10493) );
  XNOR U20721 ( .A(n10026), .B(n10022), .Z(n10494) );
  XNOR U20722 ( .A(n10021), .B(n10017), .Z(n10495) );
  XNOR U20723 ( .A(n10016), .B(n10012), .Z(n10496) );
  XNOR U20724 ( .A(n10011), .B(n10007), .Z(n10497) );
  XNOR U20725 ( .A(n10006), .B(n10002), .Z(n10498) );
  XNOR U20726 ( .A(n10001), .B(n9997), .Z(n10499) );
  XNOR U20727 ( .A(n9996), .B(n9992), .Z(n10500) );
  XNOR U20728 ( .A(n9991), .B(n9987), .Z(n10501) );
  XNOR U20729 ( .A(n9986), .B(n9982), .Z(n10502) );
  XNOR U20730 ( .A(n9981), .B(n9977), .Z(n10503) );
  XNOR U20731 ( .A(n9976), .B(n9972), .Z(n10504) );
  XNOR U20732 ( .A(n9971), .B(n9967), .Z(n10505) );
  XNOR U20733 ( .A(n9966), .B(n9962), .Z(n10506) );
  XNOR U20734 ( .A(n9961), .B(n9957), .Z(n10507) );
  XNOR U20735 ( .A(n9956), .B(n9952), .Z(n10508) );
  XNOR U20736 ( .A(n9951), .B(n9947), .Z(n10509) );
  XNOR U20737 ( .A(n9946), .B(n9942), .Z(n10510) );
  XNOR U20738 ( .A(n9941), .B(n9937), .Z(n10511) );
  XNOR U20739 ( .A(n9936), .B(n9932), .Z(n10512) );
  XNOR U20740 ( .A(n9931), .B(n9927), .Z(n10513) );
  XNOR U20741 ( .A(n9926), .B(n9922), .Z(n10514) );
  XNOR U20742 ( .A(n9921), .B(n9917), .Z(n10515) );
  XNOR U20743 ( .A(n9916), .B(n9912), .Z(n10516) );
  XNOR U20744 ( .A(n9911), .B(n9907), .Z(n10517) );
  XNOR U20745 ( .A(n9906), .B(n9902), .Z(n10518) );
  XNOR U20746 ( .A(n9901), .B(n9897), .Z(n10519) );
  XNOR U20747 ( .A(n9896), .B(n9892), .Z(n10520) );
  XNOR U20748 ( .A(n9891), .B(n9887), .Z(n10521) );
  XNOR U20749 ( .A(n9886), .B(n9882), .Z(n10522) );
  XNOR U20750 ( .A(n9881), .B(n9877), .Z(n10523) );
  XNOR U20751 ( .A(n9876), .B(n9872), .Z(n10524) );
  XNOR U20752 ( .A(n9871), .B(n9867), .Z(n10525) );
  XNOR U20753 ( .A(n9866), .B(n9862), .Z(n10526) );
  XOR U20754 ( .A(n10527), .B(n9861), .Z(n9862) );
  AND U20755 ( .A(a[0]), .B(b[112]), .Z(n10527) );
  XNOR U20756 ( .A(n10528), .B(n9861), .Z(n9863) );
  XNOR U20757 ( .A(n10529), .B(n10530), .Z(n9861) );
  ANDN U20758 ( .B(n10531), .A(n10532), .Z(n10529) );
  AND U20759 ( .A(a[1]), .B(b[111]), .Z(n10528) );
  XNOR U20760 ( .A(n10533), .B(n9866), .Z(n9868) );
  XOR U20761 ( .A(n10534), .B(n10535), .Z(n9866) );
  ANDN U20762 ( .B(n10536), .A(n10537), .Z(n10534) );
  AND U20763 ( .A(a[2]), .B(b[110]), .Z(n10533) );
  XNOR U20764 ( .A(n10538), .B(n9871), .Z(n9873) );
  XOR U20765 ( .A(n10539), .B(n10540), .Z(n9871) );
  ANDN U20766 ( .B(n10541), .A(n10542), .Z(n10539) );
  AND U20767 ( .A(a[3]), .B(b[109]), .Z(n10538) );
  XNOR U20768 ( .A(n10543), .B(n9876), .Z(n9878) );
  XOR U20769 ( .A(n10544), .B(n10545), .Z(n9876) );
  ANDN U20770 ( .B(n10546), .A(n10547), .Z(n10544) );
  AND U20771 ( .A(a[4]), .B(b[108]), .Z(n10543) );
  XNOR U20772 ( .A(n10548), .B(n9881), .Z(n9883) );
  XOR U20773 ( .A(n10549), .B(n10550), .Z(n9881) );
  ANDN U20774 ( .B(n10551), .A(n10552), .Z(n10549) );
  AND U20775 ( .A(a[5]), .B(b[107]), .Z(n10548) );
  XNOR U20776 ( .A(n10553), .B(n9886), .Z(n9888) );
  XOR U20777 ( .A(n10554), .B(n10555), .Z(n9886) );
  ANDN U20778 ( .B(n10556), .A(n10557), .Z(n10554) );
  AND U20779 ( .A(a[6]), .B(b[106]), .Z(n10553) );
  XNOR U20780 ( .A(n10558), .B(n9891), .Z(n9893) );
  XOR U20781 ( .A(n10559), .B(n10560), .Z(n9891) );
  ANDN U20782 ( .B(n10561), .A(n10562), .Z(n10559) );
  AND U20783 ( .A(a[7]), .B(b[105]), .Z(n10558) );
  XNOR U20784 ( .A(n10563), .B(n9896), .Z(n9898) );
  XOR U20785 ( .A(n10564), .B(n10565), .Z(n9896) );
  ANDN U20786 ( .B(n10566), .A(n10567), .Z(n10564) );
  AND U20787 ( .A(a[8]), .B(b[104]), .Z(n10563) );
  XNOR U20788 ( .A(n10568), .B(n9901), .Z(n9903) );
  XOR U20789 ( .A(n10569), .B(n10570), .Z(n9901) );
  ANDN U20790 ( .B(n10571), .A(n10572), .Z(n10569) );
  AND U20791 ( .A(a[9]), .B(b[103]), .Z(n10568) );
  XNOR U20792 ( .A(n10573), .B(n9906), .Z(n9908) );
  XOR U20793 ( .A(n10574), .B(n10575), .Z(n9906) );
  ANDN U20794 ( .B(n10576), .A(n10577), .Z(n10574) );
  AND U20795 ( .A(a[10]), .B(b[102]), .Z(n10573) );
  XNOR U20796 ( .A(n10578), .B(n9911), .Z(n9913) );
  XOR U20797 ( .A(n10579), .B(n10580), .Z(n9911) );
  ANDN U20798 ( .B(n10581), .A(n10582), .Z(n10579) );
  AND U20799 ( .A(a[11]), .B(b[101]), .Z(n10578) );
  XNOR U20800 ( .A(n10583), .B(n9916), .Z(n9918) );
  XOR U20801 ( .A(n10584), .B(n10585), .Z(n9916) );
  ANDN U20802 ( .B(n10586), .A(n10587), .Z(n10584) );
  AND U20803 ( .A(a[12]), .B(b[100]), .Z(n10583) );
  XNOR U20804 ( .A(n10588), .B(n9921), .Z(n9923) );
  XOR U20805 ( .A(n10589), .B(n10590), .Z(n9921) );
  ANDN U20806 ( .B(n10591), .A(n10592), .Z(n10589) );
  AND U20807 ( .A(a[13]), .B(b[99]), .Z(n10588) );
  XNOR U20808 ( .A(n10593), .B(n9926), .Z(n9928) );
  XOR U20809 ( .A(n10594), .B(n10595), .Z(n9926) );
  ANDN U20810 ( .B(n10596), .A(n10597), .Z(n10594) );
  AND U20811 ( .A(a[14]), .B(b[98]), .Z(n10593) );
  XNOR U20812 ( .A(n10598), .B(n9931), .Z(n9933) );
  XOR U20813 ( .A(n10599), .B(n10600), .Z(n9931) );
  ANDN U20814 ( .B(n10601), .A(n10602), .Z(n10599) );
  AND U20815 ( .A(a[15]), .B(b[97]), .Z(n10598) );
  XNOR U20816 ( .A(n10603), .B(n9936), .Z(n9938) );
  XOR U20817 ( .A(n10604), .B(n10605), .Z(n9936) );
  ANDN U20818 ( .B(n10606), .A(n10607), .Z(n10604) );
  AND U20819 ( .A(a[16]), .B(b[96]), .Z(n10603) );
  XNOR U20820 ( .A(n10608), .B(n9941), .Z(n9943) );
  XOR U20821 ( .A(n10609), .B(n10610), .Z(n9941) );
  ANDN U20822 ( .B(n10611), .A(n10612), .Z(n10609) );
  AND U20823 ( .A(a[17]), .B(b[95]), .Z(n10608) );
  XNOR U20824 ( .A(n10613), .B(n9946), .Z(n9948) );
  XOR U20825 ( .A(n10614), .B(n10615), .Z(n9946) );
  ANDN U20826 ( .B(n10616), .A(n10617), .Z(n10614) );
  AND U20827 ( .A(a[18]), .B(b[94]), .Z(n10613) );
  XNOR U20828 ( .A(n10618), .B(n9951), .Z(n9953) );
  XOR U20829 ( .A(n10619), .B(n10620), .Z(n9951) );
  ANDN U20830 ( .B(n10621), .A(n10622), .Z(n10619) );
  AND U20831 ( .A(a[19]), .B(b[93]), .Z(n10618) );
  XNOR U20832 ( .A(n10623), .B(n9956), .Z(n9958) );
  XOR U20833 ( .A(n10624), .B(n10625), .Z(n9956) );
  ANDN U20834 ( .B(n10626), .A(n10627), .Z(n10624) );
  AND U20835 ( .A(a[20]), .B(b[92]), .Z(n10623) );
  XNOR U20836 ( .A(n10628), .B(n9961), .Z(n9963) );
  XOR U20837 ( .A(n10629), .B(n10630), .Z(n9961) );
  ANDN U20838 ( .B(n10631), .A(n10632), .Z(n10629) );
  AND U20839 ( .A(a[21]), .B(b[91]), .Z(n10628) );
  XNOR U20840 ( .A(n10633), .B(n9966), .Z(n9968) );
  XOR U20841 ( .A(n10634), .B(n10635), .Z(n9966) );
  ANDN U20842 ( .B(n10636), .A(n10637), .Z(n10634) );
  AND U20843 ( .A(a[22]), .B(b[90]), .Z(n10633) );
  XNOR U20844 ( .A(n10638), .B(n9971), .Z(n9973) );
  XOR U20845 ( .A(n10639), .B(n10640), .Z(n9971) );
  ANDN U20846 ( .B(n10641), .A(n10642), .Z(n10639) );
  AND U20847 ( .A(a[23]), .B(b[89]), .Z(n10638) );
  XNOR U20848 ( .A(n10643), .B(n9976), .Z(n9978) );
  XOR U20849 ( .A(n10644), .B(n10645), .Z(n9976) );
  ANDN U20850 ( .B(n10646), .A(n10647), .Z(n10644) );
  AND U20851 ( .A(a[24]), .B(b[88]), .Z(n10643) );
  XNOR U20852 ( .A(n10648), .B(n9981), .Z(n9983) );
  XOR U20853 ( .A(n10649), .B(n10650), .Z(n9981) );
  ANDN U20854 ( .B(n10651), .A(n10652), .Z(n10649) );
  AND U20855 ( .A(a[25]), .B(b[87]), .Z(n10648) );
  XNOR U20856 ( .A(n10653), .B(n9986), .Z(n9988) );
  XOR U20857 ( .A(n10654), .B(n10655), .Z(n9986) );
  ANDN U20858 ( .B(n10656), .A(n10657), .Z(n10654) );
  AND U20859 ( .A(a[26]), .B(b[86]), .Z(n10653) );
  XNOR U20860 ( .A(n10658), .B(n9991), .Z(n9993) );
  XOR U20861 ( .A(n10659), .B(n10660), .Z(n9991) );
  ANDN U20862 ( .B(n10661), .A(n10662), .Z(n10659) );
  AND U20863 ( .A(a[27]), .B(b[85]), .Z(n10658) );
  XNOR U20864 ( .A(n10663), .B(n9996), .Z(n9998) );
  XOR U20865 ( .A(n10664), .B(n10665), .Z(n9996) );
  ANDN U20866 ( .B(n10666), .A(n10667), .Z(n10664) );
  AND U20867 ( .A(a[28]), .B(b[84]), .Z(n10663) );
  XNOR U20868 ( .A(n10668), .B(n10001), .Z(n10003) );
  XOR U20869 ( .A(n10669), .B(n10670), .Z(n10001) );
  ANDN U20870 ( .B(n10671), .A(n10672), .Z(n10669) );
  AND U20871 ( .A(a[29]), .B(b[83]), .Z(n10668) );
  XNOR U20872 ( .A(n10673), .B(n10006), .Z(n10008) );
  XOR U20873 ( .A(n10674), .B(n10675), .Z(n10006) );
  ANDN U20874 ( .B(n10676), .A(n10677), .Z(n10674) );
  AND U20875 ( .A(a[30]), .B(b[82]), .Z(n10673) );
  XNOR U20876 ( .A(n10678), .B(n10011), .Z(n10013) );
  XOR U20877 ( .A(n10679), .B(n10680), .Z(n10011) );
  ANDN U20878 ( .B(n10681), .A(n10682), .Z(n10679) );
  AND U20879 ( .A(a[31]), .B(b[81]), .Z(n10678) );
  XNOR U20880 ( .A(n10683), .B(n10016), .Z(n10018) );
  XOR U20881 ( .A(n10684), .B(n10685), .Z(n10016) );
  ANDN U20882 ( .B(n10686), .A(n10687), .Z(n10684) );
  AND U20883 ( .A(a[32]), .B(b[80]), .Z(n10683) );
  XNOR U20884 ( .A(n10688), .B(n10021), .Z(n10023) );
  XOR U20885 ( .A(n10689), .B(n10690), .Z(n10021) );
  ANDN U20886 ( .B(n10691), .A(n10692), .Z(n10689) );
  AND U20887 ( .A(a[33]), .B(b[79]), .Z(n10688) );
  XNOR U20888 ( .A(n10693), .B(n10026), .Z(n10028) );
  XOR U20889 ( .A(n10694), .B(n10695), .Z(n10026) );
  ANDN U20890 ( .B(n10696), .A(n10697), .Z(n10694) );
  AND U20891 ( .A(a[34]), .B(b[78]), .Z(n10693) );
  XNOR U20892 ( .A(n10698), .B(n10031), .Z(n10033) );
  XOR U20893 ( .A(n10699), .B(n10700), .Z(n10031) );
  ANDN U20894 ( .B(n10701), .A(n10702), .Z(n10699) );
  AND U20895 ( .A(a[35]), .B(b[77]), .Z(n10698) );
  XNOR U20896 ( .A(n10703), .B(n10036), .Z(n10038) );
  XOR U20897 ( .A(n10704), .B(n10705), .Z(n10036) );
  ANDN U20898 ( .B(n10706), .A(n10707), .Z(n10704) );
  AND U20899 ( .A(a[36]), .B(b[76]), .Z(n10703) );
  XNOR U20900 ( .A(n10708), .B(n10041), .Z(n10043) );
  XOR U20901 ( .A(n10709), .B(n10710), .Z(n10041) );
  ANDN U20902 ( .B(n10711), .A(n10712), .Z(n10709) );
  AND U20903 ( .A(a[37]), .B(b[75]), .Z(n10708) );
  XNOR U20904 ( .A(n10713), .B(n10046), .Z(n10048) );
  XOR U20905 ( .A(n10714), .B(n10715), .Z(n10046) );
  ANDN U20906 ( .B(n10716), .A(n10717), .Z(n10714) );
  AND U20907 ( .A(a[38]), .B(b[74]), .Z(n10713) );
  XNOR U20908 ( .A(n10718), .B(n10051), .Z(n10053) );
  XOR U20909 ( .A(n10719), .B(n10720), .Z(n10051) );
  ANDN U20910 ( .B(n10721), .A(n10722), .Z(n10719) );
  AND U20911 ( .A(a[39]), .B(b[73]), .Z(n10718) );
  XNOR U20912 ( .A(n10723), .B(n10056), .Z(n10058) );
  XOR U20913 ( .A(n10724), .B(n10725), .Z(n10056) );
  ANDN U20914 ( .B(n10726), .A(n10727), .Z(n10724) );
  AND U20915 ( .A(a[40]), .B(b[72]), .Z(n10723) );
  XNOR U20916 ( .A(n10728), .B(n10061), .Z(n10063) );
  XOR U20917 ( .A(n10729), .B(n10730), .Z(n10061) );
  ANDN U20918 ( .B(n10731), .A(n10732), .Z(n10729) );
  AND U20919 ( .A(a[41]), .B(b[71]), .Z(n10728) );
  XNOR U20920 ( .A(n10733), .B(n10066), .Z(n10068) );
  XOR U20921 ( .A(n10734), .B(n10735), .Z(n10066) );
  ANDN U20922 ( .B(n10736), .A(n10737), .Z(n10734) );
  AND U20923 ( .A(a[42]), .B(b[70]), .Z(n10733) );
  XNOR U20924 ( .A(n10738), .B(n10071), .Z(n10073) );
  XOR U20925 ( .A(n10739), .B(n10740), .Z(n10071) );
  ANDN U20926 ( .B(n10741), .A(n10742), .Z(n10739) );
  AND U20927 ( .A(a[43]), .B(b[69]), .Z(n10738) );
  XNOR U20928 ( .A(n10743), .B(n10076), .Z(n10078) );
  XOR U20929 ( .A(n10744), .B(n10745), .Z(n10076) );
  ANDN U20930 ( .B(n10746), .A(n10747), .Z(n10744) );
  AND U20931 ( .A(a[44]), .B(b[68]), .Z(n10743) );
  XNOR U20932 ( .A(n10748), .B(n10081), .Z(n10083) );
  XOR U20933 ( .A(n10749), .B(n10750), .Z(n10081) );
  ANDN U20934 ( .B(n10751), .A(n10752), .Z(n10749) );
  AND U20935 ( .A(a[45]), .B(b[67]), .Z(n10748) );
  XNOR U20936 ( .A(n10753), .B(n10086), .Z(n10088) );
  XOR U20937 ( .A(n10754), .B(n10755), .Z(n10086) );
  ANDN U20938 ( .B(n10756), .A(n10757), .Z(n10754) );
  AND U20939 ( .A(a[46]), .B(b[66]), .Z(n10753) );
  XNOR U20940 ( .A(n10758), .B(n10091), .Z(n10093) );
  XOR U20941 ( .A(n10759), .B(n10760), .Z(n10091) );
  ANDN U20942 ( .B(n10761), .A(n10762), .Z(n10759) );
  AND U20943 ( .A(a[47]), .B(b[65]), .Z(n10758) );
  XNOR U20944 ( .A(n10763), .B(n10096), .Z(n10098) );
  XOR U20945 ( .A(n10764), .B(n10765), .Z(n10096) );
  ANDN U20946 ( .B(n10766), .A(n10767), .Z(n10764) );
  AND U20947 ( .A(a[48]), .B(b[64]), .Z(n10763) );
  XNOR U20948 ( .A(n10768), .B(n10101), .Z(n10103) );
  XOR U20949 ( .A(n10769), .B(n10770), .Z(n10101) );
  ANDN U20950 ( .B(n10771), .A(n10772), .Z(n10769) );
  AND U20951 ( .A(a[49]), .B(b[63]), .Z(n10768) );
  XNOR U20952 ( .A(n10773), .B(n10106), .Z(n10108) );
  XOR U20953 ( .A(n10774), .B(n10775), .Z(n10106) );
  ANDN U20954 ( .B(n10776), .A(n10777), .Z(n10774) );
  AND U20955 ( .A(a[50]), .B(b[62]), .Z(n10773) );
  XNOR U20956 ( .A(n10778), .B(n10111), .Z(n10113) );
  XOR U20957 ( .A(n10779), .B(n10780), .Z(n10111) );
  ANDN U20958 ( .B(n10781), .A(n10782), .Z(n10779) );
  AND U20959 ( .A(a[51]), .B(b[61]), .Z(n10778) );
  XNOR U20960 ( .A(n10783), .B(n10116), .Z(n10118) );
  XOR U20961 ( .A(n10784), .B(n10785), .Z(n10116) );
  ANDN U20962 ( .B(n10786), .A(n10787), .Z(n10784) );
  AND U20963 ( .A(a[52]), .B(b[60]), .Z(n10783) );
  XNOR U20964 ( .A(n10788), .B(n10121), .Z(n10123) );
  XOR U20965 ( .A(n10789), .B(n10790), .Z(n10121) );
  ANDN U20966 ( .B(n10791), .A(n10792), .Z(n10789) );
  AND U20967 ( .A(a[53]), .B(b[59]), .Z(n10788) );
  XNOR U20968 ( .A(n10793), .B(n10126), .Z(n10128) );
  XOR U20969 ( .A(n10794), .B(n10795), .Z(n10126) );
  ANDN U20970 ( .B(n10796), .A(n10797), .Z(n10794) );
  AND U20971 ( .A(a[54]), .B(b[58]), .Z(n10793) );
  XNOR U20972 ( .A(n10798), .B(n10131), .Z(n10133) );
  XOR U20973 ( .A(n10799), .B(n10800), .Z(n10131) );
  ANDN U20974 ( .B(n10801), .A(n10802), .Z(n10799) );
  AND U20975 ( .A(a[55]), .B(b[57]), .Z(n10798) );
  XNOR U20976 ( .A(n10803), .B(n10136), .Z(n10138) );
  XOR U20977 ( .A(n10804), .B(n10805), .Z(n10136) );
  ANDN U20978 ( .B(n10806), .A(n10807), .Z(n10804) );
  AND U20979 ( .A(a[56]), .B(b[56]), .Z(n10803) );
  XNOR U20980 ( .A(n10808), .B(n10141), .Z(n10143) );
  XOR U20981 ( .A(n10809), .B(n10810), .Z(n10141) );
  ANDN U20982 ( .B(n10811), .A(n10812), .Z(n10809) );
  AND U20983 ( .A(a[57]), .B(b[55]), .Z(n10808) );
  XNOR U20984 ( .A(n10813), .B(n10146), .Z(n10148) );
  XOR U20985 ( .A(n10814), .B(n10815), .Z(n10146) );
  ANDN U20986 ( .B(n10816), .A(n10817), .Z(n10814) );
  AND U20987 ( .A(a[58]), .B(b[54]), .Z(n10813) );
  XNOR U20988 ( .A(n10818), .B(n10151), .Z(n10153) );
  XOR U20989 ( .A(n10819), .B(n10820), .Z(n10151) );
  ANDN U20990 ( .B(n10821), .A(n10822), .Z(n10819) );
  AND U20991 ( .A(a[59]), .B(b[53]), .Z(n10818) );
  XNOR U20992 ( .A(n10823), .B(n10156), .Z(n10158) );
  XOR U20993 ( .A(n10824), .B(n10825), .Z(n10156) );
  ANDN U20994 ( .B(n10826), .A(n10827), .Z(n10824) );
  AND U20995 ( .A(a[60]), .B(b[52]), .Z(n10823) );
  XNOR U20996 ( .A(n10828), .B(n10161), .Z(n10163) );
  XOR U20997 ( .A(n10829), .B(n10830), .Z(n10161) );
  ANDN U20998 ( .B(n10831), .A(n10832), .Z(n10829) );
  AND U20999 ( .A(a[61]), .B(b[51]), .Z(n10828) );
  XNOR U21000 ( .A(n10833), .B(n10166), .Z(n10168) );
  XOR U21001 ( .A(n10834), .B(n10835), .Z(n10166) );
  ANDN U21002 ( .B(n10836), .A(n10837), .Z(n10834) );
  AND U21003 ( .A(a[62]), .B(b[50]), .Z(n10833) );
  XNOR U21004 ( .A(n10838), .B(n10171), .Z(n10173) );
  XOR U21005 ( .A(n10839), .B(n10840), .Z(n10171) );
  ANDN U21006 ( .B(n10841), .A(n10842), .Z(n10839) );
  AND U21007 ( .A(a[63]), .B(b[49]), .Z(n10838) );
  XNOR U21008 ( .A(n10843), .B(n10176), .Z(n10178) );
  XOR U21009 ( .A(n10844), .B(n10845), .Z(n10176) );
  ANDN U21010 ( .B(n10846), .A(n10847), .Z(n10844) );
  AND U21011 ( .A(a[64]), .B(b[48]), .Z(n10843) );
  XNOR U21012 ( .A(n10848), .B(n10181), .Z(n10183) );
  XOR U21013 ( .A(n10849), .B(n10850), .Z(n10181) );
  ANDN U21014 ( .B(n10851), .A(n10852), .Z(n10849) );
  AND U21015 ( .A(a[65]), .B(b[47]), .Z(n10848) );
  XNOR U21016 ( .A(n10853), .B(n10186), .Z(n10188) );
  XOR U21017 ( .A(n10854), .B(n10855), .Z(n10186) );
  ANDN U21018 ( .B(n10856), .A(n10857), .Z(n10854) );
  AND U21019 ( .A(a[66]), .B(b[46]), .Z(n10853) );
  XNOR U21020 ( .A(n10858), .B(n10191), .Z(n10193) );
  XOR U21021 ( .A(n10859), .B(n10860), .Z(n10191) );
  ANDN U21022 ( .B(n10861), .A(n10862), .Z(n10859) );
  AND U21023 ( .A(a[67]), .B(b[45]), .Z(n10858) );
  XNOR U21024 ( .A(n10863), .B(n10196), .Z(n10198) );
  XOR U21025 ( .A(n10864), .B(n10865), .Z(n10196) );
  ANDN U21026 ( .B(n10866), .A(n10867), .Z(n10864) );
  AND U21027 ( .A(a[68]), .B(b[44]), .Z(n10863) );
  XNOR U21028 ( .A(n10868), .B(n10201), .Z(n10203) );
  XOR U21029 ( .A(n10869), .B(n10870), .Z(n10201) );
  ANDN U21030 ( .B(n10871), .A(n10872), .Z(n10869) );
  AND U21031 ( .A(a[69]), .B(b[43]), .Z(n10868) );
  XNOR U21032 ( .A(n10873), .B(n10206), .Z(n10208) );
  XOR U21033 ( .A(n10874), .B(n10875), .Z(n10206) );
  ANDN U21034 ( .B(n10876), .A(n10877), .Z(n10874) );
  AND U21035 ( .A(a[70]), .B(b[42]), .Z(n10873) );
  XNOR U21036 ( .A(n10878), .B(n10211), .Z(n10213) );
  XOR U21037 ( .A(n10879), .B(n10880), .Z(n10211) );
  ANDN U21038 ( .B(n10881), .A(n10882), .Z(n10879) );
  AND U21039 ( .A(a[71]), .B(b[41]), .Z(n10878) );
  XNOR U21040 ( .A(n10883), .B(n10216), .Z(n10218) );
  XOR U21041 ( .A(n10884), .B(n10885), .Z(n10216) );
  ANDN U21042 ( .B(n10886), .A(n10887), .Z(n10884) );
  AND U21043 ( .A(a[72]), .B(b[40]), .Z(n10883) );
  XNOR U21044 ( .A(n10888), .B(n10221), .Z(n10223) );
  XOR U21045 ( .A(n10889), .B(n10890), .Z(n10221) );
  ANDN U21046 ( .B(n10891), .A(n10892), .Z(n10889) );
  AND U21047 ( .A(a[73]), .B(b[39]), .Z(n10888) );
  XNOR U21048 ( .A(n10893), .B(n10226), .Z(n10228) );
  XOR U21049 ( .A(n10894), .B(n10895), .Z(n10226) );
  ANDN U21050 ( .B(n10896), .A(n10897), .Z(n10894) );
  AND U21051 ( .A(a[74]), .B(b[38]), .Z(n10893) );
  XNOR U21052 ( .A(n10898), .B(n10231), .Z(n10233) );
  XOR U21053 ( .A(n10899), .B(n10900), .Z(n10231) );
  ANDN U21054 ( .B(n10901), .A(n10902), .Z(n10899) );
  AND U21055 ( .A(a[75]), .B(b[37]), .Z(n10898) );
  XNOR U21056 ( .A(n10903), .B(n10236), .Z(n10238) );
  XOR U21057 ( .A(n10904), .B(n10905), .Z(n10236) );
  ANDN U21058 ( .B(n10906), .A(n10907), .Z(n10904) );
  AND U21059 ( .A(a[76]), .B(b[36]), .Z(n10903) );
  XNOR U21060 ( .A(n10908), .B(n10241), .Z(n10243) );
  XOR U21061 ( .A(n10909), .B(n10910), .Z(n10241) );
  ANDN U21062 ( .B(n10911), .A(n10912), .Z(n10909) );
  AND U21063 ( .A(a[77]), .B(b[35]), .Z(n10908) );
  XNOR U21064 ( .A(n10913), .B(n10246), .Z(n10248) );
  XOR U21065 ( .A(n10914), .B(n10915), .Z(n10246) );
  ANDN U21066 ( .B(n10916), .A(n10917), .Z(n10914) );
  AND U21067 ( .A(a[78]), .B(b[34]), .Z(n10913) );
  XNOR U21068 ( .A(n10918), .B(n10251), .Z(n10253) );
  XOR U21069 ( .A(n10919), .B(n10920), .Z(n10251) );
  ANDN U21070 ( .B(n10921), .A(n10922), .Z(n10919) );
  AND U21071 ( .A(a[79]), .B(b[33]), .Z(n10918) );
  XNOR U21072 ( .A(n10923), .B(n10256), .Z(n10258) );
  XOR U21073 ( .A(n10924), .B(n10925), .Z(n10256) );
  ANDN U21074 ( .B(n10926), .A(n10927), .Z(n10924) );
  AND U21075 ( .A(a[80]), .B(b[32]), .Z(n10923) );
  XNOR U21076 ( .A(n10928), .B(n10261), .Z(n10263) );
  XOR U21077 ( .A(n10929), .B(n10930), .Z(n10261) );
  ANDN U21078 ( .B(n10931), .A(n10932), .Z(n10929) );
  AND U21079 ( .A(a[81]), .B(b[31]), .Z(n10928) );
  XNOR U21080 ( .A(n10933), .B(n10266), .Z(n10268) );
  XOR U21081 ( .A(n10934), .B(n10935), .Z(n10266) );
  ANDN U21082 ( .B(n10936), .A(n10937), .Z(n10934) );
  AND U21083 ( .A(a[82]), .B(b[30]), .Z(n10933) );
  XNOR U21084 ( .A(n10938), .B(n10271), .Z(n10273) );
  XOR U21085 ( .A(n10939), .B(n10940), .Z(n10271) );
  ANDN U21086 ( .B(n10941), .A(n10942), .Z(n10939) );
  AND U21087 ( .A(a[83]), .B(b[29]), .Z(n10938) );
  XNOR U21088 ( .A(n10943), .B(n10276), .Z(n10278) );
  XOR U21089 ( .A(n10944), .B(n10945), .Z(n10276) );
  ANDN U21090 ( .B(n10946), .A(n10947), .Z(n10944) );
  AND U21091 ( .A(a[84]), .B(b[28]), .Z(n10943) );
  XNOR U21092 ( .A(n10948), .B(n10281), .Z(n10283) );
  XOR U21093 ( .A(n10949), .B(n10950), .Z(n10281) );
  ANDN U21094 ( .B(n10951), .A(n10952), .Z(n10949) );
  AND U21095 ( .A(a[85]), .B(b[27]), .Z(n10948) );
  XNOR U21096 ( .A(n10953), .B(n10286), .Z(n10288) );
  XOR U21097 ( .A(n10954), .B(n10955), .Z(n10286) );
  ANDN U21098 ( .B(n10956), .A(n10957), .Z(n10954) );
  AND U21099 ( .A(a[86]), .B(b[26]), .Z(n10953) );
  XNOR U21100 ( .A(n10958), .B(n10291), .Z(n10293) );
  XOR U21101 ( .A(n10959), .B(n10960), .Z(n10291) );
  ANDN U21102 ( .B(n10961), .A(n10962), .Z(n10959) );
  AND U21103 ( .A(a[87]), .B(b[25]), .Z(n10958) );
  XNOR U21104 ( .A(n10963), .B(n10296), .Z(n10298) );
  XOR U21105 ( .A(n10964), .B(n10965), .Z(n10296) );
  ANDN U21106 ( .B(n10966), .A(n10967), .Z(n10964) );
  AND U21107 ( .A(a[88]), .B(b[24]), .Z(n10963) );
  XNOR U21108 ( .A(n10968), .B(n10301), .Z(n10303) );
  XOR U21109 ( .A(n10969), .B(n10970), .Z(n10301) );
  ANDN U21110 ( .B(n10971), .A(n10972), .Z(n10969) );
  AND U21111 ( .A(a[89]), .B(b[23]), .Z(n10968) );
  XNOR U21112 ( .A(n10973), .B(n10306), .Z(n10308) );
  XOR U21113 ( .A(n10974), .B(n10975), .Z(n10306) );
  ANDN U21114 ( .B(n10976), .A(n10977), .Z(n10974) );
  AND U21115 ( .A(a[90]), .B(b[22]), .Z(n10973) );
  XNOR U21116 ( .A(n10978), .B(n10311), .Z(n10313) );
  XOR U21117 ( .A(n10979), .B(n10980), .Z(n10311) );
  ANDN U21118 ( .B(n10981), .A(n10982), .Z(n10979) );
  AND U21119 ( .A(a[91]), .B(b[21]), .Z(n10978) );
  XNOR U21120 ( .A(n10983), .B(n10316), .Z(n10318) );
  XOR U21121 ( .A(n10984), .B(n10985), .Z(n10316) );
  ANDN U21122 ( .B(n10986), .A(n10987), .Z(n10984) );
  AND U21123 ( .A(a[92]), .B(b[20]), .Z(n10983) );
  XNOR U21124 ( .A(n10988), .B(n10321), .Z(n10323) );
  XOR U21125 ( .A(n10989), .B(n10990), .Z(n10321) );
  ANDN U21126 ( .B(n10991), .A(n10992), .Z(n10989) );
  AND U21127 ( .A(a[93]), .B(b[19]), .Z(n10988) );
  XNOR U21128 ( .A(n10993), .B(n10326), .Z(n10328) );
  XOR U21129 ( .A(n10994), .B(n10995), .Z(n10326) );
  ANDN U21130 ( .B(n10996), .A(n10997), .Z(n10994) );
  AND U21131 ( .A(a[94]), .B(b[18]), .Z(n10993) );
  XNOR U21132 ( .A(n10998), .B(n10331), .Z(n10333) );
  XOR U21133 ( .A(n10999), .B(n11000), .Z(n10331) );
  ANDN U21134 ( .B(n11001), .A(n11002), .Z(n10999) );
  AND U21135 ( .A(a[95]), .B(b[17]), .Z(n10998) );
  XNOR U21136 ( .A(n11003), .B(n10336), .Z(n10338) );
  XOR U21137 ( .A(n11004), .B(n11005), .Z(n10336) );
  ANDN U21138 ( .B(n11006), .A(n11007), .Z(n11004) );
  AND U21139 ( .A(a[96]), .B(b[16]), .Z(n11003) );
  XNOR U21140 ( .A(n11008), .B(n10341), .Z(n10343) );
  XOR U21141 ( .A(n11009), .B(n11010), .Z(n10341) );
  ANDN U21142 ( .B(n11011), .A(n11012), .Z(n11009) );
  AND U21143 ( .A(a[97]), .B(b[15]), .Z(n11008) );
  XNOR U21144 ( .A(n11013), .B(n10346), .Z(n10348) );
  XOR U21145 ( .A(n11014), .B(n11015), .Z(n10346) );
  ANDN U21146 ( .B(n11016), .A(n11017), .Z(n11014) );
  AND U21147 ( .A(a[98]), .B(b[14]), .Z(n11013) );
  XNOR U21148 ( .A(n11018), .B(n10351), .Z(n10353) );
  XOR U21149 ( .A(n11019), .B(n11020), .Z(n10351) );
  ANDN U21150 ( .B(n11021), .A(n11022), .Z(n11019) );
  AND U21151 ( .A(a[99]), .B(b[13]), .Z(n11018) );
  XNOR U21152 ( .A(n11023), .B(n10356), .Z(n10358) );
  XOR U21153 ( .A(n11024), .B(n11025), .Z(n10356) );
  ANDN U21154 ( .B(n11026), .A(n11027), .Z(n11024) );
  AND U21155 ( .A(b[12]), .B(a[100]), .Z(n11023) );
  XNOR U21156 ( .A(n11028), .B(n10361), .Z(n10363) );
  XOR U21157 ( .A(n11029), .B(n11030), .Z(n10361) );
  ANDN U21158 ( .B(n11031), .A(n11032), .Z(n11029) );
  AND U21159 ( .A(b[11]), .B(a[101]), .Z(n11028) );
  XNOR U21160 ( .A(n11033), .B(n10366), .Z(n10368) );
  XOR U21161 ( .A(n11034), .B(n11035), .Z(n10366) );
  ANDN U21162 ( .B(n11036), .A(n11037), .Z(n11034) );
  AND U21163 ( .A(b[10]), .B(a[102]), .Z(n11033) );
  XNOR U21164 ( .A(n11038), .B(n10371), .Z(n10373) );
  XOR U21165 ( .A(n11039), .B(n11040), .Z(n10371) );
  ANDN U21166 ( .B(n11041), .A(n11042), .Z(n11039) );
  AND U21167 ( .A(b[9]), .B(a[103]), .Z(n11038) );
  XNOR U21168 ( .A(n11043), .B(n10376), .Z(n10378) );
  XOR U21169 ( .A(n11044), .B(n11045), .Z(n10376) );
  ANDN U21170 ( .B(n11046), .A(n11047), .Z(n11044) );
  AND U21171 ( .A(b[8]), .B(a[104]), .Z(n11043) );
  XNOR U21172 ( .A(n11048), .B(n10381), .Z(n10383) );
  XOR U21173 ( .A(n11049), .B(n11050), .Z(n10381) );
  ANDN U21174 ( .B(n11051), .A(n11052), .Z(n11049) );
  AND U21175 ( .A(b[7]), .B(a[105]), .Z(n11048) );
  XNOR U21176 ( .A(n11053), .B(n10386), .Z(n10388) );
  XOR U21177 ( .A(n11054), .B(n11055), .Z(n10386) );
  ANDN U21178 ( .B(n11056), .A(n11057), .Z(n11054) );
  AND U21179 ( .A(b[6]), .B(a[106]), .Z(n11053) );
  XNOR U21180 ( .A(n11058), .B(n10391), .Z(n10393) );
  XOR U21181 ( .A(n11059), .B(n11060), .Z(n10391) );
  ANDN U21182 ( .B(n11061), .A(n11062), .Z(n11059) );
  AND U21183 ( .A(b[5]), .B(a[107]), .Z(n11058) );
  XNOR U21184 ( .A(n11063), .B(n10396), .Z(n10398) );
  XOR U21185 ( .A(n11064), .B(n11065), .Z(n10396) );
  ANDN U21186 ( .B(n11066), .A(n11067), .Z(n11064) );
  AND U21187 ( .A(b[4]), .B(a[108]), .Z(n11063) );
  XNOR U21188 ( .A(n11068), .B(n11069), .Z(n10410) );
  NANDN U21189 ( .A(n11070), .B(n11071), .Z(n11069) );
  XNOR U21190 ( .A(n11072), .B(n10401), .Z(n10403) );
  XNOR U21191 ( .A(n11073), .B(n11074), .Z(n10401) );
  AND U21192 ( .A(n11075), .B(n11076), .Z(n11073) );
  AND U21193 ( .A(b[3]), .B(a[109]), .Z(n11072) );
  NAND U21194 ( .A(a[112]), .B(b[0]), .Z(n9746) );
  XNOR U21195 ( .A(n10416), .B(n10417), .Z(c[111]) );
  XNOR U21196 ( .A(n11070), .B(n11071), .Z(n10417) );
  XOR U21197 ( .A(n11068), .B(n11077), .Z(n11071) );
  NAND U21198 ( .A(b[1]), .B(a[110]), .Z(n11077) );
  XOR U21199 ( .A(n11076), .B(n11078), .Z(n11070) );
  XOR U21200 ( .A(n11068), .B(n11075), .Z(n11078) );
  XNOR U21201 ( .A(n11079), .B(n11074), .Z(n11075) );
  AND U21202 ( .A(b[2]), .B(a[109]), .Z(n11079) );
  NANDN U21203 ( .A(n11080), .B(n11081), .Z(n11068) );
  XOR U21204 ( .A(n11074), .B(n11066), .Z(n11082) );
  XNOR U21205 ( .A(n11065), .B(n11061), .Z(n11083) );
  XNOR U21206 ( .A(n11060), .B(n11056), .Z(n11084) );
  XNOR U21207 ( .A(n11055), .B(n11051), .Z(n11085) );
  XNOR U21208 ( .A(n11050), .B(n11046), .Z(n11086) );
  XNOR U21209 ( .A(n11045), .B(n11041), .Z(n11087) );
  XNOR U21210 ( .A(n11040), .B(n11036), .Z(n11088) );
  XNOR U21211 ( .A(n11035), .B(n11031), .Z(n11089) );
  XNOR U21212 ( .A(n11030), .B(n11026), .Z(n11090) );
  XNOR U21213 ( .A(n11025), .B(n11021), .Z(n11091) );
  XNOR U21214 ( .A(n11020), .B(n11016), .Z(n11092) );
  XNOR U21215 ( .A(n11015), .B(n11011), .Z(n11093) );
  XNOR U21216 ( .A(n11010), .B(n11006), .Z(n11094) );
  XNOR U21217 ( .A(n11005), .B(n11001), .Z(n11095) );
  XNOR U21218 ( .A(n11000), .B(n10996), .Z(n11096) );
  XNOR U21219 ( .A(n10995), .B(n10991), .Z(n11097) );
  XNOR U21220 ( .A(n10990), .B(n10986), .Z(n11098) );
  XNOR U21221 ( .A(n10985), .B(n10981), .Z(n11099) );
  XNOR U21222 ( .A(n10980), .B(n10976), .Z(n11100) );
  XNOR U21223 ( .A(n10975), .B(n10971), .Z(n11101) );
  XNOR U21224 ( .A(n10970), .B(n10966), .Z(n11102) );
  XNOR U21225 ( .A(n10965), .B(n10961), .Z(n11103) );
  XNOR U21226 ( .A(n10960), .B(n10956), .Z(n11104) );
  XNOR U21227 ( .A(n10955), .B(n10951), .Z(n11105) );
  XNOR U21228 ( .A(n10950), .B(n10946), .Z(n11106) );
  XNOR U21229 ( .A(n10945), .B(n10941), .Z(n11107) );
  XNOR U21230 ( .A(n10940), .B(n10936), .Z(n11108) );
  XNOR U21231 ( .A(n10935), .B(n10931), .Z(n11109) );
  XNOR U21232 ( .A(n10930), .B(n10926), .Z(n11110) );
  XNOR U21233 ( .A(n10925), .B(n10921), .Z(n11111) );
  XNOR U21234 ( .A(n10920), .B(n10916), .Z(n11112) );
  XNOR U21235 ( .A(n10915), .B(n10911), .Z(n11113) );
  XNOR U21236 ( .A(n10910), .B(n10906), .Z(n11114) );
  XNOR U21237 ( .A(n10905), .B(n10901), .Z(n11115) );
  XNOR U21238 ( .A(n10900), .B(n10896), .Z(n11116) );
  XNOR U21239 ( .A(n10895), .B(n10891), .Z(n11117) );
  XNOR U21240 ( .A(n10890), .B(n10886), .Z(n11118) );
  XNOR U21241 ( .A(n10885), .B(n10881), .Z(n11119) );
  XNOR U21242 ( .A(n10880), .B(n10876), .Z(n11120) );
  XNOR U21243 ( .A(n10875), .B(n10871), .Z(n11121) );
  XNOR U21244 ( .A(n10870), .B(n10866), .Z(n11122) );
  XNOR U21245 ( .A(n10865), .B(n10861), .Z(n11123) );
  XNOR U21246 ( .A(n10860), .B(n10856), .Z(n11124) );
  XNOR U21247 ( .A(n10855), .B(n10851), .Z(n11125) );
  XNOR U21248 ( .A(n10850), .B(n10846), .Z(n11126) );
  XNOR U21249 ( .A(n10845), .B(n10841), .Z(n11127) );
  XNOR U21250 ( .A(n10840), .B(n10836), .Z(n11128) );
  XNOR U21251 ( .A(n10835), .B(n10831), .Z(n11129) );
  XNOR U21252 ( .A(n10830), .B(n10826), .Z(n11130) );
  XNOR U21253 ( .A(n10825), .B(n10821), .Z(n11131) );
  XNOR U21254 ( .A(n10820), .B(n10816), .Z(n11132) );
  XNOR U21255 ( .A(n10815), .B(n10811), .Z(n11133) );
  XNOR U21256 ( .A(n10810), .B(n10806), .Z(n11134) );
  XNOR U21257 ( .A(n10805), .B(n10801), .Z(n11135) );
  XNOR U21258 ( .A(n10800), .B(n10796), .Z(n11136) );
  XNOR U21259 ( .A(n10795), .B(n10791), .Z(n11137) );
  XNOR U21260 ( .A(n10790), .B(n10786), .Z(n11138) );
  XNOR U21261 ( .A(n10785), .B(n10781), .Z(n11139) );
  XNOR U21262 ( .A(n10780), .B(n10776), .Z(n11140) );
  XNOR U21263 ( .A(n10775), .B(n10771), .Z(n11141) );
  XNOR U21264 ( .A(n10770), .B(n10766), .Z(n11142) );
  XNOR U21265 ( .A(n10765), .B(n10761), .Z(n11143) );
  XNOR U21266 ( .A(n10760), .B(n10756), .Z(n11144) );
  XNOR U21267 ( .A(n10755), .B(n10751), .Z(n11145) );
  XNOR U21268 ( .A(n10750), .B(n10746), .Z(n11146) );
  XNOR U21269 ( .A(n10745), .B(n10741), .Z(n11147) );
  XNOR U21270 ( .A(n10740), .B(n10736), .Z(n11148) );
  XNOR U21271 ( .A(n10735), .B(n10731), .Z(n11149) );
  XNOR U21272 ( .A(n10730), .B(n10726), .Z(n11150) );
  XNOR U21273 ( .A(n10725), .B(n10721), .Z(n11151) );
  XNOR U21274 ( .A(n10720), .B(n10716), .Z(n11152) );
  XNOR U21275 ( .A(n10715), .B(n10711), .Z(n11153) );
  XNOR U21276 ( .A(n10710), .B(n10706), .Z(n11154) );
  XNOR U21277 ( .A(n10705), .B(n10701), .Z(n11155) );
  XNOR U21278 ( .A(n10700), .B(n10696), .Z(n11156) );
  XNOR U21279 ( .A(n10695), .B(n10691), .Z(n11157) );
  XNOR U21280 ( .A(n10690), .B(n10686), .Z(n11158) );
  XNOR U21281 ( .A(n10685), .B(n10681), .Z(n11159) );
  XNOR U21282 ( .A(n10680), .B(n10676), .Z(n11160) );
  XNOR U21283 ( .A(n10675), .B(n10671), .Z(n11161) );
  XNOR U21284 ( .A(n10670), .B(n10666), .Z(n11162) );
  XNOR U21285 ( .A(n10665), .B(n10661), .Z(n11163) );
  XNOR U21286 ( .A(n10660), .B(n10656), .Z(n11164) );
  XNOR U21287 ( .A(n10655), .B(n10651), .Z(n11165) );
  XNOR U21288 ( .A(n10650), .B(n10646), .Z(n11166) );
  XNOR U21289 ( .A(n10645), .B(n10641), .Z(n11167) );
  XNOR U21290 ( .A(n10640), .B(n10636), .Z(n11168) );
  XNOR U21291 ( .A(n10635), .B(n10631), .Z(n11169) );
  XNOR U21292 ( .A(n10630), .B(n10626), .Z(n11170) );
  XNOR U21293 ( .A(n10625), .B(n10621), .Z(n11171) );
  XNOR U21294 ( .A(n10620), .B(n10616), .Z(n11172) );
  XNOR U21295 ( .A(n10615), .B(n10611), .Z(n11173) );
  XNOR U21296 ( .A(n10610), .B(n10606), .Z(n11174) );
  XNOR U21297 ( .A(n10605), .B(n10601), .Z(n11175) );
  XNOR U21298 ( .A(n10600), .B(n10596), .Z(n11176) );
  XNOR U21299 ( .A(n10595), .B(n10591), .Z(n11177) );
  XNOR U21300 ( .A(n10590), .B(n10586), .Z(n11178) );
  XNOR U21301 ( .A(n10585), .B(n10581), .Z(n11179) );
  XNOR U21302 ( .A(n10580), .B(n10576), .Z(n11180) );
  XNOR U21303 ( .A(n10575), .B(n10571), .Z(n11181) );
  XNOR U21304 ( .A(n10570), .B(n10566), .Z(n11182) );
  XNOR U21305 ( .A(n10565), .B(n10561), .Z(n11183) );
  XNOR U21306 ( .A(n10560), .B(n10556), .Z(n11184) );
  XNOR U21307 ( .A(n10555), .B(n10551), .Z(n11185) );
  XNOR U21308 ( .A(n10550), .B(n10546), .Z(n11186) );
  XNOR U21309 ( .A(n10545), .B(n10541), .Z(n11187) );
  XNOR U21310 ( .A(n10540), .B(n10536), .Z(n11188) );
  XNOR U21311 ( .A(n10535), .B(n10531), .Z(n11189) );
  XNOR U21312 ( .A(n11190), .B(n10530), .Z(n10531) );
  AND U21313 ( .A(a[0]), .B(b[111]), .Z(n11190) );
  XOR U21314 ( .A(n11191), .B(n10530), .Z(n10532) );
  XNOR U21315 ( .A(n11192), .B(n11193), .Z(n10530) );
  ANDN U21316 ( .B(n11194), .A(n11195), .Z(n11192) );
  AND U21317 ( .A(a[1]), .B(b[110]), .Z(n11191) );
  XNOR U21318 ( .A(n11196), .B(n10535), .Z(n10537) );
  XOR U21319 ( .A(n11197), .B(n11198), .Z(n10535) );
  ANDN U21320 ( .B(n11199), .A(n11200), .Z(n11197) );
  AND U21321 ( .A(a[2]), .B(b[109]), .Z(n11196) );
  XNOR U21322 ( .A(n11201), .B(n10540), .Z(n10542) );
  XOR U21323 ( .A(n11202), .B(n11203), .Z(n10540) );
  ANDN U21324 ( .B(n11204), .A(n11205), .Z(n11202) );
  AND U21325 ( .A(a[3]), .B(b[108]), .Z(n11201) );
  XNOR U21326 ( .A(n11206), .B(n10545), .Z(n10547) );
  XOR U21327 ( .A(n11207), .B(n11208), .Z(n10545) );
  ANDN U21328 ( .B(n11209), .A(n11210), .Z(n11207) );
  AND U21329 ( .A(a[4]), .B(b[107]), .Z(n11206) );
  XNOR U21330 ( .A(n11211), .B(n10550), .Z(n10552) );
  XOR U21331 ( .A(n11212), .B(n11213), .Z(n10550) );
  ANDN U21332 ( .B(n11214), .A(n11215), .Z(n11212) );
  AND U21333 ( .A(a[5]), .B(b[106]), .Z(n11211) );
  XNOR U21334 ( .A(n11216), .B(n10555), .Z(n10557) );
  XOR U21335 ( .A(n11217), .B(n11218), .Z(n10555) );
  ANDN U21336 ( .B(n11219), .A(n11220), .Z(n11217) );
  AND U21337 ( .A(a[6]), .B(b[105]), .Z(n11216) );
  XNOR U21338 ( .A(n11221), .B(n10560), .Z(n10562) );
  XOR U21339 ( .A(n11222), .B(n11223), .Z(n10560) );
  ANDN U21340 ( .B(n11224), .A(n11225), .Z(n11222) );
  AND U21341 ( .A(a[7]), .B(b[104]), .Z(n11221) );
  XNOR U21342 ( .A(n11226), .B(n10565), .Z(n10567) );
  XOR U21343 ( .A(n11227), .B(n11228), .Z(n10565) );
  ANDN U21344 ( .B(n11229), .A(n11230), .Z(n11227) );
  AND U21345 ( .A(a[8]), .B(b[103]), .Z(n11226) );
  XNOR U21346 ( .A(n11231), .B(n10570), .Z(n10572) );
  XOR U21347 ( .A(n11232), .B(n11233), .Z(n10570) );
  ANDN U21348 ( .B(n11234), .A(n11235), .Z(n11232) );
  AND U21349 ( .A(a[9]), .B(b[102]), .Z(n11231) );
  XNOR U21350 ( .A(n11236), .B(n10575), .Z(n10577) );
  XOR U21351 ( .A(n11237), .B(n11238), .Z(n10575) );
  ANDN U21352 ( .B(n11239), .A(n11240), .Z(n11237) );
  AND U21353 ( .A(a[10]), .B(b[101]), .Z(n11236) );
  XNOR U21354 ( .A(n11241), .B(n10580), .Z(n10582) );
  XOR U21355 ( .A(n11242), .B(n11243), .Z(n10580) );
  ANDN U21356 ( .B(n11244), .A(n11245), .Z(n11242) );
  AND U21357 ( .A(a[11]), .B(b[100]), .Z(n11241) );
  XNOR U21358 ( .A(n11246), .B(n10585), .Z(n10587) );
  XOR U21359 ( .A(n11247), .B(n11248), .Z(n10585) );
  ANDN U21360 ( .B(n11249), .A(n11250), .Z(n11247) );
  AND U21361 ( .A(a[12]), .B(b[99]), .Z(n11246) );
  XNOR U21362 ( .A(n11251), .B(n10590), .Z(n10592) );
  XOR U21363 ( .A(n11252), .B(n11253), .Z(n10590) );
  ANDN U21364 ( .B(n11254), .A(n11255), .Z(n11252) );
  AND U21365 ( .A(a[13]), .B(b[98]), .Z(n11251) );
  XNOR U21366 ( .A(n11256), .B(n10595), .Z(n10597) );
  XOR U21367 ( .A(n11257), .B(n11258), .Z(n10595) );
  ANDN U21368 ( .B(n11259), .A(n11260), .Z(n11257) );
  AND U21369 ( .A(a[14]), .B(b[97]), .Z(n11256) );
  XNOR U21370 ( .A(n11261), .B(n10600), .Z(n10602) );
  XOR U21371 ( .A(n11262), .B(n11263), .Z(n10600) );
  ANDN U21372 ( .B(n11264), .A(n11265), .Z(n11262) );
  AND U21373 ( .A(a[15]), .B(b[96]), .Z(n11261) );
  XNOR U21374 ( .A(n11266), .B(n10605), .Z(n10607) );
  XOR U21375 ( .A(n11267), .B(n11268), .Z(n10605) );
  ANDN U21376 ( .B(n11269), .A(n11270), .Z(n11267) );
  AND U21377 ( .A(a[16]), .B(b[95]), .Z(n11266) );
  XNOR U21378 ( .A(n11271), .B(n10610), .Z(n10612) );
  XOR U21379 ( .A(n11272), .B(n11273), .Z(n10610) );
  ANDN U21380 ( .B(n11274), .A(n11275), .Z(n11272) );
  AND U21381 ( .A(a[17]), .B(b[94]), .Z(n11271) );
  XNOR U21382 ( .A(n11276), .B(n10615), .Z(n10617) );
  XOR U21383 ( .A(n11277), .B(n11278), .Z(n10615) );
  ANDN U21384 ( .B(n11279), .A(n11280), .Z(n11277) );
  AND U21385 ( .A(a[18]), .B(b[93]), .Z(n11276) );
  XNOR U21386 ( .A(n11281), .B(n10620), .Z(n10622) );
  XOR U21387 ( .A(n11282), .B(n11283), .Z(n10620) );
  ANDN U21388 ( .B(n11284), .A(n11285), .Z(n11282) );
  AND U21389 ( .A(a[19]), .B(b[92]), .Z(n11281) );
  XNOR U21390 ( .A(n11286), .B(n10625), .Z(n10627) );
  XOR U21391 ( .A(n11287), .B(n11288), .Z(n10625) );
  ANDN U21392 ( .B(n11289), .A(n11290), .Z(n11287) );
  AND U21393 ( .A(a[20]), .B(b[91]), .Z(n11286) );
  XNOR U21394 ( .A(n11291), .B(n10630), .Z(n10632) );
  XOR U21395 ( .A(n11292), .B(n11293), .Z(n10630) );
  ANDN U21396 ( .B(n11294), .A(n11295), .Z(n11292) );
  AND U21397 ( .A(a[21]), .B(b[90]), .Z(n11291) );
  XNOR U21398 ( .A(n11296), .B(n10635), .Z(n10637) );
  XOR U21399 ( .A(n11297), .B(n11298), .Z(n10635) );
  ANDN U21400 ( .B(n11299), .A(n11300), .Z(n11297) );
  AND U21401 ( .A(a[22]), .B(b[89]), .Z(n11296) );
  XNOR U21402 ( .A(n11301), .B(n10640), .Z(n10642) );
  XOR U21403 ( .A(n11302), .B(n11303), .Z(n10640) );
  ANDN U21404 ( .B(n11304), .A(n11305), .Z(n11302) );
  AND U21405 ( .A(a[23]), .B(b[88]), .Z(n11301) );
  XNOR U21406 ( .A(n11306), .B(n10645), .Z(n10647) );
  XOR U21407 ( .A(n11307), .B(n11308), .Z(n10645) );
  ANDN U21408 ( .B(n11309), .A(n11310), .Z(n11307) );
  AND U21409 ( .A(a[24]), .B(b[87]), .Z(n11306) );
  XNOR U21410 ( .A(n11311), .B(n10650), .Z(n10652) );
  XOR U21411 ( .A(n11312), .B(n11313), .Z(n10650) );
  ANDN U21412 ( .B(n11314), .A(n11315), .Z(n11312) );
  AND U21413 ( .A(a[25]), .B(b[86]), .Z(n11311) );
  XNOR U21414 ( .A(n11316), .B(n10655), .Z(n10657) );
  XOR U21415 ( .A(n11317), .B(n11318), .Z(n10655) );
  ANDN U21416 ( .B(n11319), .A(n11320), .Z(n11317) );
  AND U21417 ( .A(a[26]), .B(b[85]), .Z(n11316) );
  XNOR U21418 ( .A(n11321), .B(n10660), .Z(n10662) );
  XOR U21419 ( .A(n11322), .B(n11323), .Z(n10660) );
  ANDN U21420 ( .B(n11324), .A(n11325), .Z(n11322) );
  AND U21421 ( .A(a[27]), .B(b[84]), .Z(n11321) );
  XNOR U21422 ( .A(n11326), .B(n10665), .Z(n10667) );
  XOR U21423 ( .A(n11327), .B(n11328), .Z(n10665) );
  ANDN U21424 ( .B(n11329), .A(n11330), .Z(n11327) );
  AND U21425 ( .A(a[28]), .B(b[83]), .Z(n11326) );
  XNOR U21426 ( .A(n11331), .B(n10670), .Z(n10672) );
  XOR U21427 ( .A(n11332), .B(n11333), .Z(n10670) );
  ANDN U21428 ( .B(n11334), .A(n11335), .Z(n11332) );
  AND U21429 ( .A(a[29]), .B(b[82]), .Z(n11331) );
  XNOR U21430 ( .A(n11336), .B(n10675), .Z(n10677) );
  XOR U21431 ( .A(n11337), .B(n11338), .Z(n10675) );
  ANDN U21432 ( .B(n11339), .A(n11340), .Z(n11337) );
  AND U21433 ( .A(a[30]), .B(b[81]), .Z(n11336) );
  XNOR U21434 ( .A(n11341), .B(n10680), .Z(n10682) );
  XOR U21435 ( .A(n11342), .B(n11343), .Z(n10680) );
  ANDN U21436 ( .B(n11344), .A(n11345), .Z(n11342) );
  AND U21437 ( .A(a[31]), .B(b[80]), .Z(n11341) );
  XNOR U21438 ( .A(n11346), .B(n10685), .Z(n10687) );
  XOR U21439 ( .A(n11347), .B(n11348), .Z(n10685) );
  ANDN U21440 ( .B(n11349), .A(n11350), .Z(n11347) );
  AND U21441 ( .A(a[32]), .B(b[79]), .Z(n11346) );
  XNOR U21442 ( .A(n11351), .B(n10690), .Z(n10692) );
  XOR U21443 ( .A(n11352), .B(n11353), .Z(n10690) );
  ANDN U21444 ( .B(n11354), .A(n11355), .Z(n11352) );
  AND U21445 ( .A(a[33]), .B(b[78]), .Z(n11351) );
  XNOR U21446 ( .A(n11356), .B(n10695), .Z(n10697) );
  XOR U21447 ( .A(n11357), .B(n11358), .Z(n10695) );
  ANDN U21448 ( .B(n11359), .A(n11360), .Z(n11357) );
  AND U21449 ( .A(a[34]), .B(b[77]), .Z(n11356) );
  XNOR U21450 ( .A(n11361), .B(n10700), .Z(n10702) );
  XOR U21451 ( .A(n11362), .B(n11363), .Z(n10700) );
  ANDN U21452 ( .B(n11364), .A(n11365), .Z(n11362) );
  AND U21453 ( .A(a[35]), .B(b[76]), .Z(n11361) );
  XNOR U21454 ( .A(n11366), .B(n10705), .Z(n10707) );
  XOR U21455 ( .A(n11367), .B(n11368), .Z(n10705) );
  ANDN U21456 ( .B(n11369), .A(n11370), .Z(n11367) );
  AND U21457 ( .A(a[36]), .B(b[75]), .Z(n11366) );
  XNOR U21458 ( .A(n11371), .B(n10710), .Z(n10712) );
  XOR U21459 ( .A(n11372), .B(n11373), .Z(n10710) );
  ANDN U21460 ( .B(n11374), .A(n11375), .Z(n11372) );
  AND U21461 ( .A(a[37]), .B(b[74]), .Z(n11371) );
  XNOR U21462 ( .A(n11376), .B(n10715), .Z(n10717) );
  XOR U21463 ( .A(n11377), .B(n11378), .Z(n10715) );
  ANDN U21464 ( .B(n11379), .A(n11380), .Z(n11377) );
  AND U21465 ( .A(a[38]), .B(b[73]), .Z(n11376) );
  XNOR U21466 ( .A(n11381), .B(n10720), .Z(n10722) );
  XOR U21467 ( .A(n11382), .B(n11383), .Z(n10720) );
  ANDN U21468 ( .B(n11384), .A(n11385), .Z(n11382) );
  AND U21469 ( .A(a[39]), .B(b[72]), .Z(n11381) );
  XNOR U21470 ( .A(n11386), .B(n10725), .Z(n10727) );
  XOR U21471 ( .A(n11387), .B(n11388), .Z(n10725) );
  ANDN U21472 ( .B(n11389), .A(n11390), .Z(n11387) );
  AND U21473 ( .A(a[40]), .B(b[71]), .Z(n11386) );
  XNOR U21474 ( .A(n11391), .B(n10730), .Z(n10732) );
  XOR U21475 ( .A(n11392), .B(n11393), .Z(n10730) );
  ANDN U21476 ( .B(n11394), .A(n11395), .Z(n11392) );
  AND U21477 ( .A(a[41]), .B(b[70]), .Z(n11391) );
  XNOR U21478 ( .A(n11396), .B(n10735), .Z(n10737) );
  XOR U21479 ( .A(n11397), .B(n11398), .Z(n10735) );
  ANDN U21480 ( .B(n11399), .A(n11400), .Z(n11397) );
  AND U21481 ( .A(a[42]), .B(b[69]), .Z(n11396) );
  XNOR U21482 ( .A(n11401), .B(n10740), .Z(n10742) );
  XOR U21483 ( .A(n11402), .B(n11403), .Z(n10740) );
  ANDN U21484 ( .B(n11404), .A(n11405), .Z(n11402) );
  AND U21485 ( .A(a[43]), .B(b[68]), .Z(n11401) );
  XNOR U21486 ( .A(n11406), .B(n10745), .Z(n10747) );
  XOR U21487 ( .A(n11407), .B(n11408), .Z(n10745) );
  ANDN U21488 ( .B(n11409), .A(n11410), .Z(n11407) );
  AND U21489 ( .A(a[44]), .B(b[67]), .Z(n11406) );
  XNOR U21490 ( .A(n11411), .B(n10750), .Z(n10752) );
  XOR U21491 ( .A(n11412), .B(n11413), .Z(n10750) );
  ANDN U21492 ( .B(n11414), .A(n11415), .Z(n11412) );
  AND U21493 ( .A(a[45]), .B(b[66]), .Z(n11411) );
  XNOR U21494 ( .A(n11416), .B(n10755), .Z(n10757) );
  XOR U21495 ( .A(n11417), .B(n11418), .Z(n10755) );
  ANDN U21496 ( .B(n11419), .A(n11420), .Z(n11417) );
  AND U21497 ( .A(a[46]), .B(b[65]), .Z(n11416) );
  XNOR U21498 ( .A(n11421), .B(n10760), .Z(n10762) );
  XOR U21499 ( .A(n11422), .B(n11423), .Z(n10760) );
  ANDN U21500 ( .B(n11424), .A(n11425), .Z(n11422) );
  AND U21501 ( .A(a[47]), .B(b[64]), .Z(n11421) );
  XNOR U21502 ( .A(n11426), .B(n10765), .Z(n10767) );
  XOR U21503 ( .A(n11427), .B(n11428), .Z(n10765) );
  ANDN U21504 ( .B(n11429), .A(n11430), .Z(n11427) );
  AND U21505 ( .A(a[48]), .B(b[63]), .Z(n11426) );
  XNOR U21506 ( .A(n11431), .B(n10770), .Z(n10772) );
  XOR U21507 ( .A(n11432), .B(n11433), .Z(n10770) );
  ANDN U21508 ( .B(n11434), .A(n11435), .Z(n11432) );
  AND U21509 ( .A(a[49]), .B(b[62]), .Z(n11431) );
  XNOR U21510 ( .A(n11436), .B(n10775), .Z(n10777) );
  XOR U21511 ( .A(n11437), .B(n11438), .Z(n10775) );
  ANDN U21512 ( .B(n11439), .A(n11440), .Z(n11437) );
  AND U21513 ( .A(a[50]), .B(b[61]), .Z(n11436) );
  XNOR U21514 ( .A(n11441), .B(n10780), .Z(n10782) );
  XOR U21515 ( .A(n11442), .B(n11443), .Z(n10780) );
  ANDN U21516 ( .B(n11444), .A(n11445), .Z(n11442) );
  AND U21517 ( .A(a[51]), .B(b[60]), .Z(n11441) );
  XNOR U21518 ( .A(n11446), .B(n10785), .Z(n10787) );
  XOR U21519 ( .A(n11447), .B(n11448), .Z(n10785) );
  ANDN U21520 ( .B(n11449), .A(n11450), .Z(n11447) );
  AND U21521 ( .A(a[52]), .B(b[59]), .Z(n11446) );
  XNOR U21522 ( .A(n11451), .B(n10790), .Z(n10792) );
  XOR U21523 ( .A(n11452), .B(n11453), .Z(n10790) );
  ANDN U21524 ( .B(n11454), .A(n11455), .Z(n11452) );
  AND U21525 ( .A(a[53]), .B(b[58]), .Z(n11451) );
  XNOR U21526 ( .A(n11456), .B(n10795), .Z(n10797) );
  XOR U21527 ( .A(n11457), .B(n11458), .Z(n10795) );
  ANDN U21528 ( .B(n11459), .A(n11460), .Z(n11457) );
  AND U21529 ( .A(a[54]), .B(b[57]), .Z(n11456) );
  XNOR U21530 ( .A(n11461), .B(n10800), .Z(n10802) );
  XOR U21531 ( .A(n11462), .B(n11463), .Z(n10800) );
  ANDN U21532 ( .B(n11464), .A(n11465), .Z(n11462) );
  AND U21533 ( .A(a[55]), .B(b[56]), .Z(n11461) );
  XNOR U21534 ( .A(n11466), .B(n10805), .Z(n10807) );
  XOR U21535 ( .A(n11467), .B(n11468), .Z(n10805) );
  ANDN U21536 ( .B(n11469), .A(n11470), .Z(n11467) );
  AND U21537 ( .A(a[56]), .B(b[55]), .Z(n11466) );
  XNOR U21538 ( .A(n11471), .B(n10810), .Z(n10812) );
  XOR U21539 ( .A(n11472), .B(n11473), .Z(n10810) );
  ANDN U21540 ( .B(n11474), .A(n11475), .Z(n11472) );
  AND U21541 ( .A(a[57]), .B(b[54]), .Z(n11471) );
  XNOR U21542 ( .A(n11476), .B(n10815), .Z(n10817) );
  XOR U21543 ( .A(n11477), .B(n11478), .Z(n10815) );
  ANDN U21544 ( .B(n11479), .A(n11480), .Z(n11477) );
  AND U21545 ( .A(a[58]), .B(b[53]), .Z(n11476) );
  XNOR U21546 ( .A(n11481), .B(n10820), .Z(n10822) );
  XOR U21547 ( .A(n11482), .B(n11483), .Z(n10820) );
  ANDN U21548 ( .B(n11484), .A(n11485), .Z(n11482) );
  AND U21549 ( .A(a[59]), .B(b[52]), .Z(n11481) );
  XNOR U21550 ( .A(n11486), .B(n10825), .Z(n10827) );
  XOR U21551 ( .A(n11487), .B(n11488), .Z(n10825) );
  ANDN U21552 ( .B(n11489), .A(n11490), .Z(n11487) );
  AND U21553 ( .A(a[60]), .B(b[51]), .Z(n11486) );
  XNOR U21554 ( .A(n11491), .B(n10830), .Z(n10832) );
  XOR U21555 ( .A(n11492), .B(n11493), .Z(n10830) );
  ANDN U21556 ( .B(n11494), .A(n11495), .Z(n11492) );
  AND U21557 ( .A(a[61]), .B(b[50]), .Z(n11491) );
  XNOR U21558 ( .A(n11496), .B(n10835), .Z(n10837) );
  XOR U21559 ( .A(n11497), .B(n11498), .Z(n10835) );
  ANDN U21560 ( .B(n11499), .A(n11500), .Z(n11497) );
  AND U21561 ( .A(a[62]), .B(b[49]), .Z(n11496) );
  XNOR U21562 ( .A(n11501), .B(n10840), .Z(n10842) );
  XOR U21563 ( .A(n11502), .B(n11503), .Z(n10840) );
  ANDN U21564 ( .B(n11504), .A(n11505), .Z(n11502) );
  AND U21565 ( .A(a[63]), .B(b[48]), .Z(n11501) );
  XNOR U21566 ( .A(n11506), .B(n10845), .Z(n10847) );
  XOR U21567 ( .A(n11507), .B(n11508), .Z(n10845) );
  ANDN U21568 ( .B(n11509), .A(n11510), .Z(n11507) );
  AND U21569 ( .A(a[64]), .B(b[47]), .Z(n11506) );
  XNOR U21570 ( .A(n11511), .B(n10850), .Z(n10852) );
  XOR U21571 ( .A(n11512), .B(n11513), .Z(n10850) );
  ANDN U21572 ( .B(n11514), .A(n11515), .Z(n11512) );
  AND U21573 ( .A(a[65]), .B(b[46]), .Z(n11511) );
  XNOR U21574 ( .A(n11516), .B(n10855), .Z(n10857) );
  XOR U21575 ( .A(n11517), .B(n11518), .Z(n10855) );
  ANDN U21576 ( .B(n11519), .A(n11520), .Z(n11517) );
  AND U21577 ( .A(a[66]), .B(b[45]), .Z(n11516) );
  XNOR U21578 ( .A(n11521), .B(n10860), .Z(n10862) );
  XOR U21579 ( .A(n11522), .B(n11523), .Z(n10860) );
  ANDN U21580 ( .B(n11524), .A(n11525), .Z(n11522) );
  AND U21581 ( .A(a[67]), .B(b[44]), .Z(n11521) );
  XNOR U21582 ( .A(n11526), .B(n10865), .Z(n10867) );
  XOR U21583 ( .A(n11527), .B(n11528), .Z(n10865) );
  ANDN U21584 ( .B(n11529), .A(n11530), .Z(n11527) );
  AND U21585 ( .A(a[68]), .B(b[43]), .Z(n11526) );
  XNOR U21586 ( .A(n11531), .B(n10870), .Z(n10872) );
  XOR U21587 ( .A(n11532), .B(n11533), .Z(n10870) );
  ANDN U21588 ( .B(n11534), .A(n11535), .Z(n11532) );
  AND U21589 ( .A(a[69]), .B(b[42]), .Z(n11531) );
  XNOR U21590 ( .A(n11536), .B(n10875), .Z(n10877) );
  XOR U21591 ( .A(n11537), .B(n11538), .Z(n10875) );
  ANDN U21592 ( .B(n11539), .A(n11540), .Z(n11537) );
  AND U21593 ( .A(a[70]), .B(b[41]), .Z(n11536) );
  XNOR U21594 ( .A(n11541), .B(n10880), .Z(n10882) );
  XOR U21595 ( .A(n11542), .B(n11543), .Z(n10880) );
  ANDN U21596 ( .B(n11544), .A(n11545), .Z(n11542) );
  AND U21597 ( .A(a[71]), .B(b[40]), .Z(n11541) );
  XNOR U21598 ( .A(n11546), .B(n10885), .Z(n10887) );
  XOR U21599 ( .A(n11547), .B(n11548), .Z(n10885) );
  ANDN U21600 ( .B(n11549), .A(n11550), .Z(n11547) );
  AND U21601 ( .A(a[72]), .B(b[39]), .Z(n11546) );
  XNOR U21602 ( .A(n11551), .B(n10890), .Z(n10892) );
  XOR U21603 ( .A(n11552), .B(n11553), .Z(n10890) );
  ANDN U21604 ( .B(n11554), .A(n11555), .Z(n11552) );
  AND U21605 ( .A(a[73]), .B(b[38]), .Z(n11551) );
  XNOR U21606 ( .A(n11556), .B(n10895), .Z(n10897) );
  XOR U21607 ( .A(n11557), .B(n11558), .Z(n10895) );
  ANDN U21608 ( .B(n11559), .A(n11560), .Z(n11557) );
  AND U21609 ( .A(a[74]), .B(b[37]), .Z(n11556) );
  XNOR U21610 ( .A(n11561), .B(n10900), .Z(n10902) );
  XOR U21611 ( .A(n11562), .B(n11563), .Z(n10900) );
  ANDN U21612 ( .B(n11564), .A(n11565), .Z(n11562) );
  AND U21613 ( .A(a[75]), .B(b[36]), .Z(n11561) );
  XNOR U21614 ( .A(n11566), .B(n10905), .Z(n10907) );
  XOR U21615 ( .A(n11567), .B(n11568), .Z(n10905) );
  ANDN U21616 ( .B(n11569), .A(n11570), .Z(n11567) );
  AND U21617 ( .A(a[76]), .B(b[35]), .Z(n11566) );
  XNOR U21618 ( .A(n11571), .B(n10910), .Z(n10912) );
  XOR U21619 ( .A(n11572), .B(n11573), .Z(n10910) );
  ANDN U21620 ( .B(n11574), .A(n11575), .Z(n11572) );
  AND U21621 ( .A(a[77]), .B(b[34]), .Z(n11571) );
  XNOR U21622 ( .A(n11576), .B(n10915), .Z(n10917) );
  XOR U21623 ( .A(n11577), .B(n11578), .Z(n10915) );
  ANDN U21624 ( .B(n11579), .A(n11580), .Z(n11577) );
  AND U21625 ( .A(a[78]), .B(b[33]), .Z(n11576) );
  XNOR U21626 ( .A(n11581), .B(n10920), .Z(n10922) );
  XOR U21627 ( .A(n11582), .B(n11583), .Z(n10920) );
  ANDN U21628 ( .B(n11584), .A(n11585), .Z(n11582) );
  AND U21629 ( .A(a[79]), .B(b[32]), .Z(n11581) );
  XNOR U21630 ( .A(n11586), .B(n10925), .Z(n10927) );
  XOR U21631 ( .A(n11587), .B(n11588), .Z(n10925) );
  ANDN U21632 ( .B(n11589), .A(n11590), .Z(n11587) );
  AND U21633 ( .A(a[80]), .B(b[31]), .Z(n11586) );
  XNOR U21634 ( .A(n11591), .B(n10930), .Z(n10932) );
  XOR U21635 ( .A(n11592), .B(n11593), .Z(n10930) );
  ANDN U21636 ( .B(n11594), .A(n11595), .Z(n11592) );
  AND U21637 ( .A(a[81]), .B(b[30]), .Z(n11591) );
  XNOR U21638 ( .A(n11596), .B(n10935), .Z(n10937) );
  XOR U21639 ( .A(n11597), .B(n11598), .Z(n10935) );
  ANDN U21640 ( .B(n11599), .A(n11600), .Z(n11597) );
  AND U21641 ( .A(a[82]), .B(b[29]), .Z(n11596) );
  XNOR U21642 ( .A(n11601), .B(n10940), .Z(n10942) );
  XOR U21643 ( .A(n11602), .B(n11603), .Z(n10940) );
  ANDN U21644 ( .B(n11604), .A(n11605), .Z(n11602) );
  AND U21645 ( .A(a[83]), .B(b[28]), .Z(n11601) );
  XNOR U21646 ( .A(n11606), .B(n10945), .Z(n10947) );
  XOR U21647 ( .A(n11607), .B(n11608), .Z(n10945) );
  ANDN U21648 ( .B(n11609), .A(n11610), .Z(n11607) );
  AND U21649 ( .A(a[84]), .B(b[27]), .Z(n11606) );
  XNOR U21650 ( .A(n11611), .B(n10950), .Z(n10952) );
  XOR U21651 ( .A(n11612), .B(n11613), .Z(n10950) );
  ANDN U21652 ( .B(n11614), .A(n11615), .Z(n11612) );
  AND U21653 ( .A(a[85]), .B(b[26]), .Z(n11611) );
  XNOR U21654 ( .A(n11616), .B(n10955), .Z(n10957) );
  XOR U21655 ( .A(n11617), .B(n11618), .Z(n10955) );
  ANDN U21656 ( .B(n11619), .A(n11620), .Z(n11617) );
  AND U21657 ( .A(a[86]), .B(b[25]), .Z(n11616) );
  XNOR U21658 ( .A(n11621), .B(n10960), .Z(n10962) );
  XOR U21659 ( .A(n11622), .B(n11623), .Z(n10960) );
  ANDN U21660 ( .B(n11624), .A(n11625), .Z(n11622) );
  AND U21661 ( .A(a[87]), .B(b[24]), .Z(n11621) );
  XNOR U21662 ( .A(n11626), .B(n10965), .Z(n10967) );
  XOR U21663 ( .A(n11627), .B(n11628), .Z(n10965) );
  ANDN U21664 ( .B(n11629), .A(n11630), .Z(n11627) );
  AND U21665 ( .A(a[88]), .B(b[23]), .Z(n11626) );
  XNOR U21666 ( .A(n11631), .B(n10970), .Z(n10972) );
  XOR U21667 ( .A(n11632), .B(n11633), .Z(n10970) );
  ANDN U21668 ( .B(n11634), .A(n11635), .Z(n11632) );
  AND U21669 ( .A(a[89]), .B(b[22]), .Z(n11631) );
  XNOR U21670 ( .A(n11636), .B(n10975), .Z(n10977) );
  XOR U21671 ( .A(n11637), .B(n11638), .Z(n10975) );
  ANDN U21672 ( .B(n11639), .A(n11640), .Z(n11637) );
  AND U21673 ( .A(a[90]), .B(b[21]), .Z(n11636) );
  XNOR U21674 ( .A(n11641), .B(n10980), .Z(n10982) );
  XOR U21675 ( .A(n11642), .B(n11643), .Z(n10980) );
  ANDN U21676 ( .B(n11644), .A(n11645), .Z(n11642) );
  AND U21677 ( .A(a[91]), .B(b[20]), .Z(n11641) );
  XNOR U21678 ( .A(n11646), .B(n10985), .Z(n10987) );
  XOR U21679 ( .A(n11647), .B(n11648), .Z(n10985) );
  ANDN U21680 ( .B(n11649), .A(n11650), .Z(n11647) );
  AND U21681 ( .A(a[92]), .B(b[19]), .Z(n11646) );
  XNOR U21682 ( .A(n11651), .B(n10990), .Z(n10992) );
  XOR U21683 ( .A(n11652), .B(n11653), .Z(n10990) );
  ANDN U21684 ( .B(n11654), .A(n11655), .Z(n11652) );
  AND U21685 ( .A(a[93]), .B(b[18]), .Z(n11651) );
  XNOR U21686 ( .A(n11656), .B(n10995), .Z(n10997) );
  XOR U21687 ( .A(n11657), .B(n11658), .Z(n10995) );
  ANDN U21688 ( .B(n11659), .A(n11660), .Z(n11657) );
  AND U21689 ( .A(a[94]), .B(b[17]), .Z(n11656) );
  XNOR U21690 ( .A(n11661), .B(n11000), .Z(n11002) );
  XOR U21691 ( .A(n11662), .B(n11663), .Z(n11000) );
  ANDN U21692 ( .B(n11664), .A(n11665), .Z(n11662) );
  AND U21693 ( .A(a[95]), .B(b[16]), .Z(n11661) );
  XNOR U21694 ( .A(n11666), .B(n11005), .Z(n11007) );
  XOR U21695 ( .A(n11667), .B(n11668), .Z(n11005) );
  ANDN U21696 ( .B(n11669), .A(n11670), .Z(n11667) );
  AND U21697 ( .A(a[96]), .B(b[15]), .Z(n11666) );
  XNOR U21698 ( .A(n11671), .B(n11010), .Z(n11012) );
  XOR U21699 ( .A(n11672), .B(n11673), .Z(n11010) );
  ANDN U21700 ( .B(n11674), .A(n11675), .Z(n11672) );
  AND U21701 ( .A(a[97]), .B(b[14]), .Z(n11671) );
  XNOR U21702 ( .A(n11676), .B(n11015), .Z(n11017) );
  XOR U21703 ( .A(n11677), .B(n11678), .Z(n11015) );
  ANDN U21704 ( .B(n11679), .A(n11680), .Z(n11677) );
  AND U21705 ( .A(a[98]), .B(b[13]), .Z(n11676) );
  XNOR U21706 ( .A(n11681), .B(n11020), .Z(n11022) );
  XOR U21707 ( .A(n11682), .B(n11683), .Z(n11020) );
  ANDN U21708 ( .B(n11684), .A(n11685), .Z(n11682) );
  AND U21709 ( .A(a[99]), .B(b[12]), .Z(n11681) );
  XNOR U21710 ( .A(n11686), .B(n11025), .Z(n11027) );
  XOR U21711 ( .A(n11687), .B(n11688), .Z(n11025) );
  ANDN U21712 ( .B(n11689), .A(n11690), .Z(n11687) );
  AND U21713 ( .A(b[11]), .B(a[100]), .Z(n11686) );
  XNOR U21714 ( .A(n11691), .B(n11030), .Z(n11032) );
  XOR U21715 ( .A(n11692), .B(n11693), .Z(n11030) );
  ANDN U21716 ( .B(n11694), .A(n11695), .Z(n11692) );
  AND U21717 ( .A(b[10]), .B(a[101]), .Z(n11691) );
  XNOR U21718 ( .A(n11696), .B(n11035), .Z(n11037) );
  XOR U21719 ( .A(n11697), .B(n11698), .Z(n11035) );
  ANDN U21720 ( .B(n11699), .A(n11700), .Z(n11697) );
  AND U21721 ( .A(b[9]), .B(a[102]), .Z(n11696) );
  XNOR U21722 ( .A(n11701), .B(n11040), .Z(n11042) );
  XOR U21723 ( .A(n11702), .B(n11703), .Z(n11040) );
  ANDN U21724 ( .B(n11704), .A(n11705), .Z(n11702) );
  AND U21725 ( .A(b[8]), .B(a[103]), .Z(n11701) );
  XNOR U21726 ( .A(n11706), .B(n11045), .Z(n11047) );
  XOR U21727 ( .A(n11707), .B(n11708), .Z(n11045) );
  ANDN U21728 ( .B(n11709), .A(n11710), .Z(n11707) );
  AND U21729 ( .A(b[7]), .B(a[104]), .Z(n11706) );
  XNOR U21730 ( .A(n11711), .B(n11050), .Z(n11052) );
  XOR U21731 ( .A(n11712), .B(n11713), .Z(n11050) );
  ANDN U21732 ( .B(n11714), .A(n11715), .Z(n11712) );
  AND U21733 ( .A(b[6]), .B(a[105]), .Z(n11711) );
  XNOR U21734 ( .A(n11716), .B(n11055), .Z(n11057) );
  XOR U21735 ( .A(n11717), .B(n11718), .Z(n11055) );
  ANDN U21736 ( .B(n11719), .A(n11720), .Z(n11717) );
  AND U21737 ( .A(b[5]), .B(a[106]), .Z(n11716) );
  XNOR U21738 ( .A(n11721), .B(n11060), .Z(n11062) );
  XOR U21739 ( .A(n11722), .B(n11723), .Z(n11060) );
  ANDN U21740 ( .B(n11724), .A(n11725), .Z(n11722) );
  AND U21741 ( .A(b[4]), .B(a[107]), .Z(n11721) );
  XNOR U21742 ( .A(n11726), .B(n11727), .Z(n11074) );
  NANDN U21743 ( .A(n11728), .B(n11729), .Z(n11727) );
  XNOR U21744 ( .A(n11730), .B(n11065), .Z(n11067) );
  XNOR U21745 ( .A(n11731), .B(n11732), .Z(n11065) );
  AND U21746 ( .A(n11733), .B(n11734), .Z(n11731) );
  AND U21747 ( .A(b[3]), .B(a[108]), .Z(n11730) );
  NAND U21748 ( .A(a[111]), .B(b[0]), .Z(n10416) );
  XNOR U21749 ( .A(n11080), .B(n11081), .Z(c[110]) );
  XNOR U21750 ( .A(n11728), .B(n11729), .Z(n11081) );
  XOR U21751 ( .A(n11726), .B(n11735), .Z(n11729) );
  NAND U21752 ( .A(b[1]), .B(a[109]), .Z(n11735) );
  XOR U21753 ( .A(n11734), .B(n11736), .Z(n11728) );
  XOR U21754 ( .A(n11726), .B(n11733), .Z(n11736) );
  XNOR U21755 ( .A(n11737), .B(n11732), .Z(n11733) );
  AND U21756 ( .A(b[2]), .B(a[108]), .Z(n11737) );
  NANDN U21757 ( .A(n11738), .B(n11739), .Z(n11726) );
  XOR U21758 ( .A(n11732), .B(n11724), .Z(n11740) );
  XNOR U21759 ( .A(n11723), .B(n11719), .Z(n11741) );
  XNOR U21760 ( .A(n11718), .B(n11714), .Z(n11742) );
  XNOR U21761 ( .A(n11713), .B(n11709), .Z(n11743) );
  XNOR U21762 ( .A(n11708), .B(n11704), .Z(n11744) );
  XNOR U21763 ( .A(n11703), .B(n11699), .Z(n11745) );
  XNOR U21764 ( .A(n11698), .B(n11694), .Z(n11746) );
  XNOR U21765 ( .A(n11693), .B(n11689), .Z(n11747) );
  XNOR U21766 ( .A(n11688), .B(n11684), .Z(n11748) );
  XNOR U21767 ( .A(n11683), .B(n11679), .Z(n11749) );
  XNOR U21768 ( .A(n11678), .B(n11674), .Z(n11750) );
  XNOR U21769 ( .A(n11673), .B(n11669), .Z(n11751) );
  XNOR U21770 ( .A(n11668), .B(n11664), .Z(n11752) );
  XNOR U21771 ( .A(n11663), .B(n11659), .Z(n11753) );
  XNOR U21772 ( .A(n11658), .B(n11654), .Z(n11754) );
  XNOR U21773 ( .A(n11653), .B(n11649), .Z(n11755) );
  XNOR U21774 ( .A(n11648), .B(n11644), .Z(n11756) );
  XNOR U21775 ( .A(n11643), .B(n11639), .Z(n11757) );
  XNOR U21776 ( .A(n11638), .B(n11634), .Z(n11758) );
  XNOR U21777 ( .A(n11633), .B(n11629), .Z(n11759) );
  XNOR U21778 ( .A(n11628), .B(n11624), .Z(n11760) );
  XNOR U21779 ( .A(n11623), .B(n11619), .Z(n11761) );
  XNOR U21780 ( .A(n11618), .B(n11614), .Z(n11762) );
  XNOR U21781 ( .A(n11613), .B(n11609), .Z(n11763) );
  XNOR U21782 ( .A(n11608), .B(n11604), .Z(n11764) );
  XNOR U21783 ( .A(n11603), .B(n11599), .Z(n11765) );
  XNOR U21784 ( .A(n11598), .B(n11594), .Z(n11766) );
  XNOR U21785 ( .A(n11593), .B(n11589), .Z(n11767) );
  XNOR U21786 ( .A(n11588), .B(n11584), .Z(n11768) );
  XNOR U21787 ( .A(n11583), .B(n11579), .Z(n11769) );
  XNOR U21788 ( .A(n11578), .B(n11574), .Z(n11770) );
  XNOR U21789 ( .A(n11573), .B(n11569), .Z(n11771) );
  XNOR U21790 ( .A(n11568), .B(n11564), .Z(n11772) );
  XNOR U21791 ( .A(n11563), .B(n11559), .Z(n11773) );
  XNOR U21792 ( .A(n11558), .B(n11554), .Z(n11774) );
  XNOR U21793 ( .A(n11553), .B(n11549), .Z(n11775) );
  XNOR U21794 ( .A(n11548), .B(n11544), .Z(n11776) );
  XNOR U21795 ( .A(n11543), .B(n11539), .Z(n11777) );
  XNOR U21796 ( .A(n11538), .B(n11534), .Z(n11778) );
  XNOR U21797 ( .A(n11533), .B(n11529), .Z(n11779) );
  XNOR U21798 ( .A(n11528), .B(n11524), .Z(n11780) );
  XNOR U21799 ( .A(n11523), .B(n11519), .Z(n11781) );
  XNOR U21800 ( .A(n11518), .B(n11514), .Z(n11782) );
  XNOR U21801 ( .A(n11513), .B(n11509), .Z(n11783) );
  XNOR U21802 ( .A(n11508), .B(n11504), .Z(n11784) );
  XNOR U21803 ( .A(n11503), .B(n11499), .Z(n11785) );
  XNOR U21804 ( .A(n11498), .B(n11494), .Z(n11786) );
  XNOR U21805 ( .A(n11493), .B(n11489), .Z(n11787) );
  XNOR U21806 ( .A(n11488), .B(n11484), .Z(n11788) );
  XNOR U21807 ( .A(n11483), .B(n11479), .Z(n11789) );
  XNOR U21808 ( .A(n11478), .B(n11474), .Z(n11790) );
  XNOR U21809 ( .A(n11473), .B(n11469), .Z(n11791) );
  XNOR U21810 ( .A(n11468), .B(n11464), .Z(n11792) );
  XNOR U21811 ( .A(n11463), .B(n11459), .Z(n11793) );
  XNOR U21812 ( .A(n11458), .B(n11454), .Z(n11794) );
  XNOR U21813 ( .A(n11453), .B(n11449), .Z(n11795) );
  XNOR U21814 ( .A(n11448), .B(n11444), .Z(n11796) );
  XNOR U21815 ( .A(n11443), .B(n11439), .Z(n11797) );
  XNOR U21816 ( .A(n11438), .B(n11434), .Z(n11798) );
  XNOR U21817 ( .A(n11433), .B(n11429), .Z(n11799) );
  XNOR U21818 ( .A(n11428), .B(n11424), .Z(n11800) );
  XNOR U21819 ( .A(n11423), .B(n11419), .Z(n11801) );
  XNOR U21820 ( .A(n11418), .B(n11414), .Z(n11802) );
  XNOR U21821 ( .A(n11413), .B(n11409), .Z(n11803) );
  XNOR U21822 ( .A(n11408), .B(n11404), .Z(n11804) );
  XNOR U21823 ( .A(n11403), .B(n11399), .Z(n11805) );
  XNOR U21824 ( .A(n11398), .B(n11394), .Z(n11806) );
  XNOR U21825 ( .A(n11393), .B(n11389), .Z(n11807) );
  XNOR U21826 ( .A(n11388), .B(n11384), .Z(n11808) );
  XNOR U21827 ( .A(n11383), .B(n11379), .Z(n11809) );
  XNOR U21828 ( .A(n11378), .B(n11374), .Z(n11810) );
  XNOR U21829 ( .A(n11373), .B(n11369), .Z(n11811) );
  XNOR U21830 ( .A(n11368), .B(n11364), .Z(n11812) );
  XNOR U21831 ( .A(n11363), .B(n11359), .Z(n11813) );
  XNOR U21832 ( .A(n11358), .B(n11354), .Z(n11814) );
  XNOR U21833 ( .A(n11353), .B(n11349), .Z(n11815) );
  XNOR U21834 ( .A(n11348), .B(n11344), .Z(n11816) );
  XNOR U21835 ( .A(n11343), .B(n11339), .Z(n11817) );
  XNOR U21836 ( .A(n11338), .B(n11334), .Z(n11818) );
  XNOR U21837 ( .A(n11333), .B(n11329), .Z(n11819) );
  XNOR U21838 ( .A(n11328), .B(n11324), .Z(n11820) );
  XNOR U21839 ( .A(n11323), .B(n11319), .Z(n11821) );
  XNOR U21840 ( .A(n11318), .B(n11314), .Z(n11822) );
  XNOR U21841 ( .A(n11313), .B(n11309), .Z(n11823) );
  XNOR U21842 ( .A(n11308), .B(n11304), .Z(n11824) );
  XNOR U21843 ( .A(n11303), .B(n11299), .Z(n11825) );
  XNOR U21844 ( .A(n11298), .B(n11294), .Z(n11826) );
  XNOR U21845 ( .A(n11293), .B(n11289), .Z(n11827) );
  XNOR U21846 ( .A(n11288), .B(n11284), .Z(n11828) );
  XNOR U21847 ( .A(n11283), .B(n11279), .Z(n11829) );
  XNOR U21848 ( .A(n11278), .B(n11274), .Z(n11830) );
  XNOR U21849 ( .A(n11273), .B(n11269), .Z(n11831) );
  XNOR U21850 ( .A(n11268), .B(n11264), .Z(n11832) );
  XNOR U21851 ( .A(n11263), .B(n11259), .Z(n11833) );
  XNOR U21852 ( .A(n11258), .B(n11254), .Z(n11834) );
  XNOR U21853 ( .A(n11253), .B(n11249), .Z(n11835) );
  XNOR U21854 ( .A(n11248), .B(n11244), .Z(n11836) );
  XNOR U21855 ( .A(n11243), .B(n11239), .Z(n11837) );
  XNOR U21856 ( .A(n11238), .B(n11234), .Z(n11838) );
  XNOR U21857 ( .A(n11233), .B(n11229), .Z(n11839) );
  XNOR U21858 ( .A(n11228), .B(n11224), .Z(n11840) );
  XNOR U21859 ( .A(n11223), .B(n11219), .Z(n11841) );
  XNOR U21860 ( .A(n11218), .B(n11214), .Z(n11842) );
  XNOR U21861 ( .A(n11213), .B(n11209), .Z(n11843) );
  XNOR U21862 ( .A(n11208), .B(n11204), .Z(n11844) );
  XNOR U21863 ( .A(n11203), .B(n11199), .Z(n11845) );
  XNOR U21864 ( .A(n11198), .B(n11194), .Z(n11846) );
  XOR U21865 ( .A(n11847), .B(n11193), .Z(n11194) );
  AND U21866 ( .A(a[0]), .B(b[110]), .Z(n11847) );
  XNOR U21867 ( .A(n11848), .B(n11193), .Z(n11195) );
  XNOR U21868 ( .A(n11849), .B(n11850), .Z(n11193) );
  ANDN U21869 ( .B(n11851), .A(n11852), .Z(n11849) );
  AND U21870 ( .A(a[1]), .B(b[109]), .Z(n11848) );
  XNOR U21871 ( .A(n11853), .B(n11198), .Z(n11200) );
  XOR U21872 ( .A(n11854), .B(n11855), .Z(n11198) );
  ANDN U21873 ( .B(n11856), .A(n11857), .Z(n11854) );
  AND U21874 ( .A(a[2]), .B(b[108]), .Z(n11853) );
  XNOR U21875 ( .A(n11858), .B(n11203), .Z(n11205) );
  XOR U21876 ( .A(n11859), .B(n11860), .Z(n11203) );
  ANDN U21877 ( .B(n11861), .A(n11862), .Z(n11859) );
  AND U21878 ( .A(a[3]), .B(b[107]), .Z(n11858) );
  XNOR U21879 ( .A(n11863), .B(n11208), .Z(n11210) );
  XOR U21880 ( .A(n11864), .B(n11865), .Z(n11208) );
  ANDN U21881 ( .B(n11866), .A(n11867), .Z(n11864) );
  AND U21882 ( .A(a[4]), .B(b[106]), .Z(n11863) );
  XNOR U21883 ( .A(n11868), .B(n11213), .Z(n11215) );
  XOR U21884 ( .A(n11869), .B(n11870), .Z(n11213) );
  ANDN U21885 ( .B(n11871), .A(n11872), .Z(n11869) );
  AND U21886 ( .A(a[5]), .B(b[105]), .Z(n11868) );
  XNOR U21887 ( .A(n11873), .B(n11218), .Z(n11220) );
  XOR U21888 ( .A(n11874), .B(n11875), .Z(n11218) );
  ANDN U21889 ( .B(n11876), .A(n11877), .Z(n11874) );
  AND U21890 ( .A(a[6]), .B(b[104]), .Z(n11873) );
  XNOR U21891 ( .A(n11878), .B(n11223), .Z(n11225) );
  XOR U21892 ( .A(n11879), .B(n11880), .Z(n11223) );
  ANDN U21893 ( .B(n11881), .A(n11882), .Z(n11879) );
  AND U21894 ( .A(a[7]), .B(b[103]), .Z(n11878) );
  XNOR U21895 ( .A(n11883), .B(n11228), .Z(n11230) );
  XOR U21896 ( .A(n11884), .B(n11885), .Z(n11228) );
  ANDN U21897 ( .B(n11886), .A(n11887), .Z(n11884) );
  AND U21898 ( .A(a[8]), .B(b[102]), .Z(n11883) );
  XNOR U21899 ( .A(n11888), .B(n11233), .Z(n11235) );
  XOR U21900 ( .A(n11889), .B(n11890), .Z(n11233) );
  ANDN U21901 ( .B(n11891), .A(n11892), .Z(n11889) );
  AND U21902 ( .A(a[9]), .B(b[101]), .Z(n11888) );
  XNOR U21903 ( .A(n11893), .B(n11238), .Z(n11240) );
  XOR U21904 ( .A(n11894), .B(n11895), .Z(n11238) );
  ANDN U21905 ( .B(n11896), .A(n11897), .Z(n11894) );
  AND U21906 ( .A(a[10]), .B(b[100]), .Z(n11893) );
  XNOR U21907 ( .A(n11898), .B(n11243), .Z(n11245) );
  XOR U21908 ( .A(n11899), .B(n11900), .Z(n11243) );
  ANDN U21909 ( .B(n11901), .A(n11902), .Z(n11899) );
  AND U21910 ( .A(a[11]), .B(b[99]), .Z(n11898) );
  XNOR U21911 ( .A(n11903), .B(n11248), .Z(n11250) );
  XOR U21912 ( .A(n11904), .B(n11905), .Z(n11248) );
  ANDN U21913 ( .B(n11906), .A(n11907), .Z(n11904) );
  AND U21914 ( .A(a[12]), .B(b[98]), .Z(n11903) );
  XNOR U21915 ( .A(n11908), .B(n11253), .Z(n11255) );
  XOR U21916 ( .A(n11909), .B(n11910), .Z(n11253) );
  ANDN U21917 ( .B(n11911), .A(n11912), .Z(n11909) );
  AND U21918 ( .A(a[13]), .B(b[97]), .Z(n11908) );
  XNOR U21919 ( .A(n11913), .B(n11258), .Z(n11260) );
  XOR U21920 ( .A(n11914), .B(n11915), .Z(n11258) );
  ANDN U21921 ( .B(n11916), .A(n11917), .Z(n11914) );
  AND U21922 ( .A(a[14]), .B(b[96]), .Z(n11913) );
  XNOR U21923 ( .A(n11918), .B(n11263), .Z(n11265) );
  XOR U21924 ( .A(n11919), .B(n11920), .Z(n11263) );
  ANDN U21925 ( .B(n11921), .A(n11922), .Z(n11919) );
  AND U21926 ( .A(a[15]), .B(b[95]), .Z(n11918) );
  XNOR U21927 ( .A(n11923), .B(n11268), .Z(n11270) );
  XOR U21928 ( .A(n11924), .B(n11925), .Z(n11268) );
  ANDN U21929 ( .B(n11926), .A(n11927), .Z(n11924) );
  AND U21930 ( .A(a[16]), .B(b[94]), .Z(n11923) );
  XNOR U21931 ( .A(n11928), .B(n11273), .Z(n11275) );
  XOR U21932 ( .A(n11929), .B(n11930), .Z(n11273) );
  ANDN U21933 ( .B(n11931), .A(n11932), .Z(n11929) );
  AND U21934 ( .A(a[17]), .B(b[93]), .Z(n11928) );
  XNOR U21935 ( .A(n11933), .B(n11278), .Z(n11280) );
  XOR U21936 ( .A(n11934), .B(n11935), .Z(n11278) );
  ANDN U21937 ( .B(n11936), .A(n11937), .Z(n11934) );
  AND U21938 ( .A(a[18]), .B(b[92]), .Z(n11933) );
  XNOR U21939 ( .A(n11938), .B(n11283), .Z(n11285) );
  XOR U21940 ( .A(n11939), .B(n11940), .Z(n11283) );
  ANDN U21941 ( .B(n11941), .A(n11942), .Z(n11939) );
  AND U21942 ( .A(a[19]), .B(b[91]), .Z(n11938) );
  XNOR U21943 ( .A(n11943), .B(n11288), .Z(n11290) );
  XOR U21944 ( .A(n11944), .B(n11945), .Z(n11288) );
  ANDN U21945 ( .B(n11946), .A(n11947), .Z(n11944) );
  AND U21946 ( .A(a[20]), .B(b[90]), .Z(n11943) );
  XNOR U21947 ( .A(n11948), .B(n11293), .Z(n11295) );
  XOR U21948 ( .A(n11949), .B(n11950), .Z(n11293) );
  ANDN U21949 ( .B(n11951), .A(n11952), .Z(n11949) );
  AND U21950 ( .A(a[21]), .B(b[89]), .Z(n11948) );
  XNOR U21951 ( .A(n11953), .B(n11298), .Z(n11300) );
  XOR U21952 ( .A(n11954), .B(n11955), .Z(n11298) );
  ANDN U21953 ( .B(n11956), .A(n11957), .Z(n11954) );
  AND U21954 ( .A(a[22]), .B(b[88]), .Z(n11953) );
  XNOR U21955 ( .A(n11958), .B(n11303), .Z(n11305) );
  XOR U21956 ( .A(n11959), .B(n11960), .Z(n11303) );
  ANDN U21957 ( .B(n11961), .A(n11962), .Z(n11959) );
  AND U21958 ( .A(a[23]), .B(b[87]), .Z(n11958) );
  XNOR U21959 ( .A(n11963), .B(n11308), .Z(n11310) );
  XOR U21960 ( .A(n11964), .B(n11965), .Z(n11308) );
  ANDN U21961 ( .B(n11966), .A(n11967), .Z(n11964) );
  AND U21962 ( .A(a[24]), .B(b[86]), .Z(n11963) );
  XNOR U21963 ( .A(n11968), .B(n11313), .Z(n11315) );
  XOR U21964 ( .A(n11969), .B(n11970), .Z(n11313) );
  ANDN U21965 ( .B(n11971), .A(n11972), .Z(n11969) );
  AND U21966 ( .A(a[25]), .B(b[85]), .Z(n11968) );
  XNOR U21967 ( .A(n11973), .B(n11318), .Z(n11320) );
  XOR U21968 ( .A(n11974), .B(n11975), .Z(n11318) );
  ANDN U21969 ( .B(n11976), .A(n11977), .Z(n11974) );
  AND U21970 ( .A(a[26]), .B(b[84]), .Z(n11973) );
  XNOR U21971 ( .A(n11978), .B(n11323), .Z(n11325) );
  XOR U21972 ( .A(n11979), .B(n11980), .Z(n11323) );
  ANDN U21973 ( .B(n11981), .A(n11982), .Z(n11979) );
  AND U21974 ( .A(a[27]), .B(b[83]), .Z(n11978) );
  XNOR U21975 ( .A(n11983), .B(n11328), .Z(n11330) );
  XOR U21976 ( .A(n11984), .B(n11985), .Z(n11328) );
  ANDN U21977 ( .B(n11986), .A(n11987), .Z(n11984) );
  AND U21978 ( .A(a[28]), .B(b[82]), .Z(n11983) );
  XNOR U21979 ( .A(n11988), .B(n11333), .Z(n11335) );
  XOR U21980 ( .A(n11989), .B(n11990), .Z(n11333) );
  ANDN U21981 ( .B(n11991), .A(n11992), .Z(n11989) );
  AND U21982 ( .A(a[29]), .B(b[81]), .Z(n11988) );
  XNOR U21983 ( .A(n11993), .B(n11338), .Z(n11340) );
  XOR U21984 ( .A(n11994), .B(n11995), .Z(n11338) );
  ANDN U21985 ( .B(n11996), .A(n11997), .Z(n11994) );
  AND U21986 ( .A(a[30]), .B(b[80]), .Z(n11993) );
  XNOR U21987 ( .A(n11998), .B(n11343), .Z(n11345) );
  XOR U21988 ( .A(n11999), .B(n12000), .Z(n11343) );
  ANDN U21989 ( .B(n12001), .A(n12002), .Z(n11999) );
  AND U21990 ( .A(a[31]), .B(b[79]), .Z(n11998) );
  XNOR U21991 ( .A(n12003), .B(n11348), .Z(n11350) );
  XOR U21992 ( .A(n12004), .B(n12005), .Z(n11348) );
  ANDN U21993 ( .B(n12006), .A(n12007), .Z(n12004) );
  AND U21994 ( .A(a[32]), .B(b[78]), .Z(n12003) );
  XNOR U21995 ( .A(n12008), .B(n11353), .Z(n11355) );
  XOR U21996 ( .A(n12009), .B(n12010), .Z(n11353) );
  ANDN U21997 ( .B(n12011), .A(n12012), .Z(n12009) );
  AND U21998 ( .A(a[33]), .B(b[77]), .Z(n12008) );
  XNOR U21999 ( .A(n12013), .B(n11358), .Z(n11360) );
  XOR U22000 ( .A(n12014), .B(n12015), .Z(n11358) );
  ANDN U22001 ( .B(n12016), .A(n12017), .Z(n12014) );
  AND U22002 ( .A(a[34]), .B(b[76]), .Z(n12013) );
  XNOR U22003 ( .A(n12018), .B(n11363), .Z(n11365) );
  XOR U22004 ( .A(n12019), .B(n12020), .Z(n11363) );
  ANDN U22005 ( .B(n12021), .A(n12022), .Z(n12019) );
  AND U22006 ( .A(a[35]), .B(b[75]), .Z(n12018) );
  XNOR U22007 ( .A(n12023), .B(n11368), .Z(n11370) );
  XOR U22008 ( .A(n12024), .B(n12025), .Z(n11368) );
  ANDN U22009 ( .B(n12026), .A(n12027), .Z(n12024) );
  AND U22010 ( .A(a[36]), .B(b[74]), .Z(n12023) );
  XNOR U22011 ( .A(n12028), .B(n11373), .Z(n11375) );
  XOR U22012 ( .A(n12029), .B(n12030), .Z(n11373) );
  ANDN U22013 ( .B(n12031), .A(n12032), .Z(n12029) );
  AND U22014 ( .A(a[37]), .B(b[73]), .Z(n12028) );
  XNOR U22015 ( .A(n12033), .B(n11378), .Z(n11380) );
  XOR U22016 ( .A(n12034), .B(n12035), .Z(n11378) );
  ANDN U22017 ( .B(n12036), .A(n12037), .Z(n12034) );
  AND U22018 ( .A(a[38]), .B(b[72]), .Z(n12033) );
  XNOR U22019 ( .A(n12038), .B(n11383), .Z(n11385) );
  XOR U22020 ( .A(n12039), .B(n12040), .Z(n11383) );
  ANDN U22021 ( .B(n12041), .A(n12042), .Z(n12039) );
  AND U22022 ( .A(a[39]), .B(b[71]), .Z(n12038) );
  XNOR U22023 ( .A(n12043), .B(n11388), .Z(n11390) );
  XOR U22024 ( .A(n12044), .B(n12045), .Z(n11388) );
  ANDN U22025 ( .B(n12046), .A(n12047), .Z(n12044) );
  AND U22026 ( .A(a[40]), .B(b[70]), .Z(n12043) );
  XNOR U22027 ( .A(n12048), .B(n11393), .Z(n11395) );
  XOR U22028 ( .A(n12049), .B(n12050), .Z(n11393) );
  ANDN U22029 ( .B(n12051), .A(n12052), .Z(n12049) );
  AND U22030 ( .A(a[41]), .B(b[69]), .Z(n12048) );
  XNOR U22031 ( .A(n12053), .B(n11398), .Z(n11400) );
  XOR U22032 ( .A(n12054), .B(n12055), .Z(n11398) );
  ANDN U22033 ( .B(n12056), .A(n12057), .Z(n12054) );
  AND U22034 ( .A(a[42]), .B(b[68]), .Z(n12053) );
  XNOR U22035 ( .A(n12058), .B(n11403), .Z(n11405) );
  XOR U22036 ( .A(n12059), .B(n12060), .Z(n11403) );
  ANDN U22037 ( .B(n12061), .A(n12062), .Z(n12059) );
  AND U22038 ( .A(a[43]), .B(b[67]), .Z(n12058) );
  XNOR U22039 ( .A(n12063), .B(n11408), .Z(n11410) );
  XOR U22040 ( .A(n12064), .B(n12065), .Z(n11408) );
  ANDN U22041 ( .B(n12066), .A(n12067), .Z(n12064) );
  AND U22042 ( .A(a[44]), .B(b[66]), .Z(n12063) );
  XNOR U22043 ( .A(n12068), .B(n11413), .Z(n11415) );
  XOR U22044 ( .A(n12069), .B(n12070), .Z(n11413) );
  ANDN U22045 ( .B(n12071), .A(n12072), .Z(n12069) );
  AND U22046 ( .A(a[45]), .B(b[65]), .Z(n12068) );
  XNOR U22047 ( .A(n12073), .B(n11418), .Z(n11420) );
  XOR U22048 ( .A(n12074), .B(n12075), .Z(n11418) );
  ANDN U22049 ( .B(n12076), .A(n12077), .Z(n12074) );
  AND U22050 ( .A(a[46]), .B(b[64]), .Z(n12073) );
  XNOR U22051 ( .A(n12078), .B(n11423), .Z(n11425) );
  XOR U22052 ( .A(n12079), .B(n12080), .Z(n11423) );
  ANDN U22053 ( .B(n12081), .A(n12082), .Z(n12079) );
  AND U22054 ( .A(a[47]), .B(b[63]), .Z(n12078) );
  XNOR U22055 ( .A(n12083), .B(n11428), .Z(n11430) );
  XOR U22056 ( .A(n12084), .B(n12085), .Z(n11428) );
  ANDN U22057 ( .B(n12086), .A(n12087), .Z(n12084) );
  AND U22058 ( .A(a[48]), .B(b[62]), .Z(n12083) );
  XNOR U22059 ( .A(n12088), .B(n11433), .Z(n11435) );
  XOR U22060 ( .A(n12089), .B(n12090), .Z(n11433) );
  ANDN U22061 ( .B(n12091), .A(n12092), .Z(n12089) );
  AND U22062 ( .A(a[49]), .B(b[61]), .Z(n12088) );
  XNOR U22063 ( .A(n12093), .B(n11438), .Z(n11440) );
  XOR U22064 ( .A(n12094), .B(n12095), .Z(n11438) );
  ANDN U22065 ( .B(n12096), .A(n12097), .Z(n12094) );
  AND U22066 ( .A(a[50]), .B(b[60]), .Z(n12093) );
  XNOR U22067 ( .A(n12098), .B(n11443), .Z(n11445) );
  XOR U22068 ( .A(n12099), .B(n12100), .Z(n11443) );
  ANDN U22069 ( .B(n12101), .A(n12102), .Z(n12099) );
  AND U22070 ( .A(a[51]), .B(b[59]), .Z(n12098) );
  XNOR U22071 ( .A(n12103), .B(n11448), .Z(n11450) );
  XOR U22072 ( .A(n12104), .B(n12105), .Z(n11448) );
  ANDN U22073 ( .B(n12106), .A(n12107), .Z(n12104) );
  AND U22074 ( .A(a[52]), .B(b[58]), .Z(n12103) );
  XNOR U22075 ( .A(n12108), .B(n11453), .Z(n11455) );
  XOR U22076 ( .A(n12109), .B(n12110), .Z(n11453) );
  ANDN U22077 ( .B(n12111), .A(n12112), .Z(n12109) );
  AND U22078 ( .A(a[53]), .B(b[57]), .Z(n12108) );
  XNOR U22079 ( .A(n12113), .B(n11458), .Z(n11460) );
  XOR U22080 ( .A(n12114), .B(n12115), .Z(n11458) );
  ANDN U22081 ( .B(n12116), .A(n12117), .Z(n12114) );
  AND U22082 ( .A(a[54]), .B(b[56]), .Z(n12113) );
  XNOR U22083 ( .A(n12118), .B(n11463), .Z(n11465) );
  XOR U22084 ( .A(n12119), .B(n12120), .Z(n11463) );
  ANDN U22085 ( .B(n12121), .A(n12122), .Z(n12119) );
  AND U22086 ( .A(a[55]), .B(b[55]), .Z(n12118) );
  XNOR U22087 ( .A(n12123), .B(n11468), .Z(n11470) );
  XOR U22088 ( .A(n12124), .B(n12125), .Z(n11468) );
  ANDN U22089 ( .B(n12126), .A(n12127), .Z(n12124) );
  AND U22090 ( .A(a[56]), .B(b[54]), .Z(n12123) );
  XNOR U22091 ( .A(n12128), .B(n11473), .Z(n11475) );
  XOR U22092 ( .A(n12129), .B(n12130), .Z(n11473) );
  ANDN U22093 ( .B(n12131), .A(n12132), .Z(n12129) );
  AND U22094 ( .A(a[57]), .B(b[53]), .Z(n12128) );
  XNOR U22095 ( .A(n12133), .B(n11478), .Z(n11480) );
  XOR U22096 ( .A(n12134), .B(n12135), .Z(n11478) );
  ANDN U22097 ( .B(n12136), .A(n12137), .Z(n12134) );
  AND U22098 ( .A(a[58]), .B(b[52]), .Z(n12133) );
  XNOR U22099 ( .A(n12138), .B(n11483), .Z(n11485) );
  XOR U22100 ( .A(n12139), .B(n12140), .Z(n11483) );
  ANDN U22101 ( .B(n12141), .A(n12142), .Z(n12139) );
  AND U22102 ( .A(a[59]), .B(b[51]), .Z(n12138) );
  XNOR U22103 ( .A(n12143), .B(n11488), .Z(n11490) );
  XOR U22104 ( .A(n12144), .B(n12145), .Z(n11488) );
  ANDN U22105 ( .B(n12146), .A(n12147), .Z(n12144) );
  AND U22106 ( .A(a[60]), .B(b[50]), .Z(n12143) );
  XNOR U22107 ( .A(n12148), .B(n11493), .Z(n11495) );
  XOR U22108 ( .A(n12149), .B(n12150), .Z(n11493) );
  ANDN U22109 ( .B(n12151), .A(n12152), .Z(n12149) );
  AND U22110 ( .A(a[61]), .B(b[49]), .Z(n12148) );
  XNOR U22111 ( .A(n12153), .B(n11498), .Z(n11500) );
  XOR U22112 ( .A(n12154), .B(n12155), .Z(n11498) );
  ANDN U22113 ( .B(n12156), .A(n12157), .Z(n12154) );
  AND U22114 ( .A(a[62]), .B(b[48]), .Z(n12153) );
  XNOR U22115 ( .A(n12158), .B(n11503), .Z(n11505) );
  XOR U22116 ( .A(n12159), .B(n12160), .Z(n11503) );
  ANDN U22117 ( .B(n12161), .A(n12162), .Z(n12159) );
  AND U22118 ( .A(a[63]), .B(b[47]), .Z(n12158) );
  XNOR U22119 ( .A(n12163), .B(n11508), .Z(n11510) );
  XOR U22120 ( .A(n12164), .B(n12165), .Z(n11508) );
  ANDN U22121 ( .B(n12166), .A(n12167), .Z(n12164) );
  AND U22122 ( .A(a[64]), .B(b[46]), .Z(n12163) );
  XNOR U22123 ( .A(n12168), .B(n11513), .Z(n11515) );
  XOR U22124 ( .A(n12169), .B(n12170), .Z(n11513) );
  ANDN U22125 ( .B(n12171), .A(n12172), .Z(n12169) );
  AND U22126 ( .A(a[65]), .B(b[45]), .Z(n12168) );
  XNOR U22127 ( .A(n12173), .B(n11518), .Z(n11520) );
  XOR U22128 ( .A(n12174), .B(n12175), .Z(n11518) );
  ANDN U22129 ( .B(n12176), .A(n12177), .Z(n12174) );
  AND U22130 ( .A(a[66]), .B(b[44]), .Z(n12173) );
  XNOR U22131 ( .A(n12178), .B(n11523), .Z(n11525) );
  XOR U22132 ( .A(n12179), .B(n12180), .Z(n11523) );
  ANDN U22133 ( .B(n12181), .A(n12182), .Z(n12179) );
  AND U22134 ( .A(a[67]), .B(b[43]), .Z(n12178) );
  XNOR U22135 ( .A(n12183), .B(n11528), .Z(n11530) );
  XOR U22136 ( .A(n12184), .B(n12185), .Z(n11528) );
  ANDN U22137 ( .B(n12186), .A(n12187), .Z(n12184) );
  AND U22138 ( .A(a[68]), .B(b[42]), .Z(n12183) );
  XNOR U22139 ( .A(n12188), .B(n11533), .Z(n11535) );
  XOR U22140 ( .A(n12189), .B(n12190), .Z(n11533) );
  ANDN U22141 ( .B(n12191), .A(n12192), .Z(n12189) );
  AND U22142 ( .A(a[69]), .B(b[41]), .Z(n12188) );
  XNOR U22143 ( .A(n12193), .B(n11538), .Z(n11540) );
  XOR U22144 ( .A(n12194), .B(n12195), .Z(n11538) );
  ANDN U22145 ( .B(n12196), .A(n12197), .Z(n12194) );
  AND U22146 ( .A(a[70]), .B(b[40]), .Z(n12193) );
  XNOR U22147 ( .A(n12198), .B(n11543), .Z(n11545) );
  XOR U22148 ( .A(n12199), .B(n12200), .Z(n11543) );
  ANDN U22149 ( .B(n12201), .A(n12202), .Z(n12199) );
  AND U22150 ( .A(a[71]), .B(b[39]), .Z(n12198) );
  XNOR U22151 ( .A(n12203), .B(n11548), .Z(n11550) );
  XOR U22152 ( .A(n12204), .B(n12205), .Z(n11548) );
  ANDN U22153 ( .B(n12206), .A(n12207), .Z(n12204) );
  AND U22154 ( .A(a[72]), .B(b[38]), .Z(n12203) );
  XNOR U22155 ( .A(n12208), .B(n11553), .Z(n11555) );
  XOR U22156 ( .A(n12209), .B(n12210), .Z(n11553) );
  ANDN U22157 ( .B(n12211), .A(n12212), .Z(n12209) );
  AND U22158 ( .A(a[73]), .B(b[37]), .Z(n12208) );
  XNOR U22159 ( .A(n12213), .B(n11558), .Z(n11560) );
  XOR U22160 ( .A(n12214), .B(n12215), .Z(n11558) );
  ANDN U22161 ( .B(n12216), .A(n12217), .Z(n12214) );
  AND U22162 ( .A(a[74]), .B(b[36]), .Z(n12213) );
  XNOR U22163 ( .A(n12218), .B(n11563), .Z(n11565) );
  XOR U22164 ( .A(n12219), .B(n12220), .Z(n11563) );
  ANDN U22165 ( .B(n12221), .A(n12222), .Z(n12219) );
  AND U22166 ( .A(a[75]), .B(b[35]), .Z(n12218) );
  XNOR U22167 ( .A(n12223), .B(n11568), .Z(n11570) );
  XOR U22168 ( .A(n12224), .B(n12225), .Z(n11568) );
  ANDN U22169 ( .B(n12226), .A(n12227), .Z(n12224) );
  AND U22170 ( .A(a[76]), .B(b[34]), .Z(n12223) );
  XNOR U22171 ( .A(n12228), .B(n11573), .Z(n11575) );
  XOR U22172 ( .A(n12229), .B(n12230), .Z(n11573) );
  ANDN U22173 ( .B(n12231), .A(n12232), .Z(n12229) );
  AND U22174 ( .A(a[77]), .B(b[33]), .Z(n12228) );
  XNOR U22175 ( .A(n12233), .B(n11578), .Z(n11580) );
  XOR U22176 ( .A(n12234), .B(n12235), .Z(n11578) );
  ANDN U22177 ( .B(n12236), .A(n12237), .Z(n12234) );
  AND U22178 ( .A(a[78]), .B(b[32]), .Z(n12233) );
  XNOR U22179 ( .A(n12238), .B(n11583), .Z(n11585) );
  XOR U22180 ( .A(n12239), .B(n12240), .Z(n11583) );
  ANDN U22181 ( .B(n12241), .A(n12242), .Z(n12239) );
  AND U22182 ( .A(a[79]), .B(b[31]), .Z(n12238) );
  XNOR U22183 ( .A(n12243), .B(n11588), .Z(n11590) );
  XOR U22184 ( .A(n12244), .B(n12245), .Z(n11588) );
  ANDN U22185 ( .B(n12246), .A(n12247), .Z(n12244) );
  AND U22186 ( .A(a[80]), .B(b[30]), .Z(n12243) );
  XNOR U22187 ( .A(n12248), .B(n11593), .Z(n11595) );
  XOR U22188 ( .A(n12249), .B(n12250), .Z(n11593) );
  ANDN U22189 ( .B(n12251), .A(n12252), .Z(n12249) );
  AND U22190 ( .A(a[81]), .B(b[29]), .Z(n12248) );
  XNOR U22191 ( .A(n12253), .B(n11598), .Z(n11600) );
  XOR U22192 ( .A(n12254), .B(n12255), .Z(n11598) );
  ANDN U22193 ( .B(n12256), .A(n12257), .Z(n12254) );
  AND U22194 ( .A(a[82]), .B(b[28]), .Z(n12253) );
  XNOR U22195 ( .A(n12258), .B(n11603), .Z(n11605) );
  XOR U22196 ( .A(n12259), .B(n12260), .Z(n11603) );
  ANDN U22197 ( .B(n12261), .A(n12262), .Z(n12259) );
  AND U22198 ( .A(a[83]), .B(b[27]), .Z(n12258) );
  XNOR U22199 ( .A(n12263), .B(n11608), .Z(n11610) );
  XOR U22200 ( .A(n12264), .B(n12265), .Z(n11608) );
  ANDN U22201 ( .B(n12266), .A(n12267), .Z(n12264) );
  AND U22202 ( .A(a[84]), .B(b[26]), .Z(n12263) );
  XNOR U22203 ( .A(n12268), .B(n11613), .Z(n11615) );
  XOR U22204 ( .A(n12269), .B(n12270), .Z(n11613) );
  ANDN U22205 ( .B(n12271), .A(n12272), .Z(n12269) );
  AND U22206 ( .A(a[85]), .B(b[25]), .Z(n12268) );
  XNOR U22207 ( .A(n12273), .B(n11618), .Z(n11620) );
  XOR U22208 ( .A(n12274), .B(n12275), .Z(n11618) );
  ANDN U22209 ( .B(n12276), .A(n12277), .Z(n12274) );
  AND U22210 ( .A(a[86]), .B(b[24]), .Z(n12273) );
  XNOR U22211 ( .A(n12278), .B(n11623), .Z(n11625) );
  XOR U22212 ( .A(n12279), .B(n12280), .Z(n11623) );
  ANDN U22213 ( .B(n12281), .A(n12282), .Z(n12279) );
  AND U22214 ( .A(a[87]), .B(b[23]), .Z(n12278) );
  XNOR U22215 ( .A(n12283), .B(n11628), .Z(n11630) );
  XOR U22216 ( .A(n12284), .B(n12285), .Z(n11628) );
  ANDN U22217 ( .B(n12286), .A(n12287), .Z(n12284) );
  AND U22218 ( .A(a[88]), .B(b[22]), .Z(n12283) );
  XNOR U22219 ( .A(n12288), .B(n11633), .Z(n11635) );
  XOR U22220 ( .A(n12289), .B(n12290), .Z(n11633) );
  ANDN U22221 ( .B(n12291), .A(n12292), .Z(n12289) );
  AND U22222 ( .A(a[89]), .B(b[21]), .Z(n12288) );
  XNOR U22223 ( .A(n12293), .B(n11638), .Z(n11640) );
  XOR U22224 ( .A(n12294), .B(n12295), .Z(n11638) );
  ANDN U22225 ( .B(n12296), .A(n12297), .Z(n12294) );
  AND U22226 ( .A(a[90]), .B(b[20]), .Z(n12293) );
  XNOR U22227 ( .A(n12298), .B(n11643), .Z(n11645) );
  XOR U22228 ( .A(n12299), .B(n12300), .Z(n11643) );
  ANDN U22229 ( .B(n12301), .A(n12302), .Z(n12299) );
  AND U22230 ( .A(a[91]), .B(b[19]), .Z(n12298) );
  XNOR U22231 ( .A(n12303), .B(n11648), .Z(n11650) );
  XOR U22232 ( .A(n12304), .B(n12305), .Z(n11648) );
  ANDN U22233 ( .B(n12306), .A(n12307), .Z(n12304) );
  AND U22234 ( .A(a[92]), .B(b[18]), .Z(n12303) );
  XNOR U22235 ( .A(n12308), .B(n11653), .Z(n11655) );
  XOR U22236 ( .A(n12309), .B(n12310), .Z(n11653) );
  ANDN U22237 ( .B(n12311), .A(n12312), .Z(n12309) );
  AND U22238 ( .A(a[93]), .B(b[17]), .Z(n12308) );
  XNOR U22239 ( .A(n12313), .B(n11658), .Z(n11660) );
  XOR U22240 ( .A(n12314), .B(n12315), .Z(n11658) );
  ANDN U22241 ( .B(n12316), .A(n12317), .Z(n12314) );
  AND U22242 ( .A(a[94]), .B(b[16]), .Z(n12313) );
  XNOR U22243 ( .A(n12318), .B(n11663), .Z(n11665) );
  XOR U22244 ( .A(n12319), .B(n12320), .Z(n11663) );
  ANDN U22245 ( .B(n12321), .A(n12322), .Z(n12319) );
  AND U22246 ( .A(a[95]), .B(b[15]), .Z(n12318) );
  XNOR U22247 ( .A(n12323), .B(n11668), .Z(n11670) );
  XOR U22248 ( .A(n12324), .B(n12325), .Z(n11668) );
  ANDN U22249 ( .B(n12326), .A(n12327), .Z(n12324) );
  AND U22250 ( .A(a[96]), .B(b[14]), .Z(n12323) );
  XNOR U22251 ( .A(n12328), .B(n11673), .Z(n11675) );
  XOR U22252 ( .A(n12329), .B(n12330), .Z(n11673) );
  ANDN U22253 ( .B(n12331), .A(n12332), .Z(n12329) );
  AND U22254 ( .A(a[97]), .B(b[13]), .Z(n12328) );
  XNOR U22255 ( .A(n12333), .B(n11678), .Z(n11680) );
  XOR U22256 ( .A(n12334), .B(n12335), .Z(n11678) );
  ANDN U22257 ( .B(n12336), .A(n12337), .Z(n12334) );
  AND U22258 ( .A(a[98]), .B(b[12]), .Z(n12333) );
  XNOR U22259 ( .A(n12338), .B(n11683), .Z(n11685) );
  XOR U22260 ( .A(n12339), .B(n12340), .Z(n11683) );
  ANDN U22261 ( .B(n12341), .A(n12342), .Z(n12339) );
  AND U22262 ( .A(a[99]), .B(b[11]), .Z(n12338) );
  XNOR U22263 ( .A(n12343), .B(n11688), .Z(n11690) );
  XOR U22264 ( .A(n12344), .B(n12345), .Z(n11688) );
  ANDN U22265 ( .B(n12346), .A(n12347), .Z(n12344) );
  AND U22266 ( .A(b[10]), .B(a[100]), .Z(n12343) );
  XNOR U22267 ( .A(n12348), .B(n11693), .Z(n11695) );
  XOR U22268 ( .A(n12349), .B(n12350), .Z(n11693) );
  ANDN U22269 ( .B(n12351), .A(n12352), .Z(n12349) );
  AND U22270 ( .A(b[9]), .B(a[101]), .Z(n12348) );
  XNOR U22271 ( .A(n12353), .B(n11698), .Z(n11700) );
  XOR U22272 ( .A(n12354), .B(n12355), .Z(n11698) );
  ANDN U22273 ( .B(n12356), .A(n12357), .Z(n12354) );
  AND U22274 ( .A(b[8]), .B(a[102]), .Z(n12353) );
  XNOR U22275 ( .A(n12358), .B(n11703), .Z(n11705) );
  XOR U22276 ( .A(n12359), .B(n12360), .Z(n11703) );
  ANDN U22277 ( .B(n12361), .A(n12362), .Z(n12359) );
  AND U22278 ( .A(b[7]), .B(a[103]), .Z(n12358) );
  XNOR U22279 ( .A(n12363), .B(n11708), .Z(n11710) );
  XOR U22280 ( .A(n12364), .B(n12365), .Z(n11708) );
  ANDN U22281 ( .B(n12366), .A(n12367), .Z(n12364) );
  AND U22282 ( .A(b[6]), .B(a[104]), .Z(n12363) );
  XNOR U22283 ( .A(n12368), .B(n11713), .Z(n11715) );
  XOR U22284 ( .A(n12369), .B(n12370), .Z(n11713) );
  ANDN U22285 ( .B(n12371), .A(n12372), .Z(n12369) );
  AND U22286 ( .A(b[5]), .B(a[105]), .Z(n12368) );
  XNOR U22287 ( .A(n12373), .B(n11718), .Z(n11720) );
  XOR U22288 ( .A(n12374), .B(n12375), .Z(n11718) );
  ANDN U22289 ( .B(n12376), .A(n12377), .Z(n12374) );
  AND U22290 ( .A(b[4]), .B(a[106]), .Z(n12373) );
  XNOR U22291 ( .A(n12378), .B(n12379), .Z(n11732) );
  NANDN U22292 ( .A(n12380), .B(n12381), .Z(n12379) );
  XNOR U22293 ( .A(n12382), .B(n11723), .Z(n11725) );
  XNOR U22294 ( .A(n12383), .B(n12384), .Z(n11723) );
  AND U22295 ( .A(n12385), .B(n12386), .Z(n12383) );
  AND U22296 ( .A(b[3]), .B(a[107]), .Z(n12382) );
  NAND U22297 ( .A(a[110]), .B(b[0]), .Z(n11080) );
  XNOR U22298 ( .A(n12387), .B(n12388), .Z(c[10]) );
  XNOR U22299 ( .A(n11738), .B(n11739), .Z(c[109]) );
  XNOR U22300 ( .A(n12380), .B(n12381), .Z(n11739) );
  XOR U22301 ( .A(n12378), .B(n12389), .Z(n12381) );
  NAND U22302 ( .A(b[1]), .B(a[108]), .Z(n12389) );
  XOR U22303 ( .A(n12386), .B(n12390), .Z(n12380) );
  XOR U22304 ( .A(n12378), .B(n12385), .Z(n12390) );
  XNOR U22305 ( .A(n12391), .B(n12384), .Z(n12385) );
  AND U22306 ( .A(b[2]), .B(a[107]), .Z(n12391) );
  NANDN U22307 ( .A(n12392), .B(n12393), .Z(n12378) );
  XOR U22308 ( .A(n12384), .B(n12376), .Z(n12394) );
  XNOR U22309 ( .A(n12375), .B(n12371), .Z(n12395) );
  XNOR U22310 ( .A(n12370), .B(n12366), .Z(n12396) );
  XNOR U22311 ( .A(n12365), .B(n12361), .Z(n12397) );
  XNOR U22312 ( .A(n12360), .B(n12356), .Z(n12398) );
  XNOR U22313 ( .A(n12355), .B(n12351), .Z(n12399) );
  XNOR U22314 ( .A(n12350), .B(n12346), .Z(n12400) );
  XNOR U22315 ( .A(n12345), .B(n12341), .Z(n12401) );
  XNOR U22316 ( .A(n12340), .B(n12336), .Z(n12402) );
  XNOR U22317 ( .A(n12335), .B(n12331), .Z(n12403) );
  XNOR U22318 ( .A(n12330), .B(n12326), .Z(n12404) );
  XNOR U22319 ( .A(n12325), .B(n12321), .Z(n12405) );
  XNOR U22320 ( .A(n12320), .B(n12316), .Z(n12406) );
  XNOR U22321 ( .A(n12315), .B(n12311), .Z(n12407) );
  XNOR U22322 ( .A(n12310), .B(n12306), .Z(n12408) );
  XNOR U22323 ( .A(n12305), .B(n12301), .Z(n12409) );
  XNOR U22324 ( .A(n12300), .B(n12296), .Z(n12410) );
  XNOR U22325 ( .A(n12295), .B(n12291), .Z(n12411) );
  XNOR U22326 ( .A(n12290), .B(n12286), .Z(n12412) );
  XNOR U22327 ( .A(n12285), .B(n12281), .Z(n12413) );
  XNOR U22328 ( .A(n12280), .B(n12276), .Z(n12414) );
  XNOR U22329 ( .A(n12275), .B(n12271), .Z(n12415) );
  XNOR U22330 ( .A(n12270), .B(n12266), .Z(n12416) );
  XNOR U22331 ( .A(n12265), .B(n12261), .Z(n12417) );
  XNOR U22332 ( .A(n12260), .B(n12256), .Z(n12418) );
  XNOR U22333 ( .A(n12255), .B(n12251), .Z(n12419) );
  XNOR U22334 ( .A(n12250), .B(n12246), .Z(n12420) );
  XNOR U22335 ( .A(n12245), .B(n12241), .Z(n12421) );
  XNOR U22336 ( .A(n12240), .B(n12236), .Z(n12422) );
  XNOR U22337 ( .A(n12235), .B(n12231), .Z(n12423) );
  XNOR U22338 ( .A(n12230), .B(n12226), .Z(n12424) );
  XNOR U22339 ( .A(n12225), .B(n12221), .Z(n12425) );
  XNOR U22340 ( .A(n12220), .B(n12216), .Z(n12426) );
  XNOR U22341 ( .A(n12215), .B(n12211), .Z(n12427) );
  XNOR U22342 ( .A(n12210), .B(n12206), .Z(n12428) );
  XNOR U22343 ( .A(n12205), .B(n12201), .Z(n12429) );
  XNOR U22344 ( .A(n12200), .B(n12196), .Z(n12430) );
  XNOR U22345 ( .A(n12195), .B(n12191), .Z(n12431) );
  XNOR U22346 ( .A(n12190), .B(n12186), .Z(n12432) );
  XNOR U22347 ( .A(n12185), .B(n12181), .Z(n12433) );
  XNOR U22348 ( .A(n12180), .B(n12176), .Z(n12434) );
  XNOR U22349 ( .A(n12175), .B(n12171), .Z(n12435) );
  XNOR U22350 ( .A(n12170), .B(n12166), .Z(n12436) );
  XNOR U22351 ( .A(n12165), .B(n12161), .Z(n12437) );
  XNOR U22352 ( .A(n12160), .B(n12156), .Z(n12438) );
  XNOR U22353 ( .A(n12155), .B(n12151), .Z(n12439) );
  XNOR U22354 ( .A(n12150), .B(n12146), .Z(n12440) );
  XNOR U22355 ( .A(n12145), .B(n12141), .Z(n12441) );
  XNOR U22356 ( .A(n12140), .B(n12136), .Z(n12442) );
  XNOR U22357 ( .A(n12135), .B(n12131), .Z(n12443) );
  XNOR U22358 ( .A(n12130), .B(n12126), .Z(n12444) );
  XNOR U22359 ( .A(n12125), .B(n12121), .Z(n12445) );
  XNOR U22360 ( .A(n12120), .B(n12116), .Z(n12446) );
  XNOR U22361 ( .A(n12115), .B(n12111), .Z(n12447) );
  XNOR U22362 ( .A(n12110), .B(n12106), .Z(n12448) );
  XNOR U22363 ( .A(n12105), .B(n12101), .Z(n12449) );
  XNOR U22364 ( .A(n12100), .B(n12096), .Z(n12450) );
  XNOR U22365 ( .A(n12095), .B(n12091), .Z(n12451) );
  XNOR U22366 ( .A(n12090), .B(n12086), .Z(n12452) );
  XNOR U22367 ( .A(n12085), .B(n12081), .Z(n12453) );
  XNOR U22368 ( .A(n12080), .B(n12076), .Z(n12454) );
  XNOR U22369 ( .A(n12075), .B(n12071), .Z(n12455) );
  XNOR U22370 ( .A(n12070), .B(n12066), .Z(n12456) );
  XNOR U22371 ( .A(n12065), .B(n12061), .Z(n12457) );
  XNOR U22372 ( .A(n12060), .B(n12056), .Z(n12458) );
  XNOR U22373 ( .A(n12055), .B(n12051), .Z(n12459) );
  XNOR U22374 ( .A(n12050), .B(n12046), .Z(n12460) );
  XNOR U22375 ( .A(n12045), .B(n12041), .Z(n12461) );
  XNOR U22376 ( .A(n12040), .B(n12036), .Z(n12462) );
  XNOR U22377 ( .A(n12035), .B(n12031), .Z(n12463) );
  XNOR U22378 ( .A(n12030), .B(n12026), .Z(n12464) );
  XNOR U22379 ( .A(n12025), .B(n12021), .Z(n12465) );
  XNOR U22380 ( .A(n12020), .B(n12016), .Z(n12466) );
  XNOR U22381 ( .A(n12015), .B(n12011), .Z(n12467) );
  XNOR U22382 ( .A(n12010), .B(n12006), .Z(n12468) );
  XNOR U22383 ( .A(n12005), .B(n12001), .Z(n12469) );
  XNOR U22384 ( .A(n12000), .B(n11996), .Z(n12470) );
  XNOR U22385 ( .A(n11995), .B(n11991), .Z(n12471) );
  XNOR U22386 ( .A(n11990), .B(n11986), .Z(n12472) );
  XNOR U22387 ( .A(n11985), .B(n11981), .Z(n12473) );
  XNOR U22388 ( .A(n11980), .B(n11976), .Z(n12474) );
  XNOR U22389 ( .A(n11975), .B(n11971), .Z(n12475) );
  XNOR U22390 ( .A(n11970), .B(n11966), .Z(n12476) );
  XNOR U22391 ( .A(n11965), .B(n11961), .Z(n12477) );
  XNOR U22392 ( .A(n11960), .B(n11956), .Z(n12478) );
  XNOR U22393 ( .A(n11955), .B(n11951), .Z(n12479) );
  XNOR U22394 ( .A(n11950), .B(n11946), .Z(n12480) );
  XNOR U22395 ( .A(n11945), .B(n11941), .Z(n12481) );
  XNOR U22396 ( .A(n11940), .B(n11936), .Z(n12482) );
  XNOR U22397 ( .A(n11935), .B(n11931), .Z(n12483) );
  XNOR U22398 ( .A(n11930), .B(n11926), .Z(n12484) );
  XNOR U22399 ( .A(n11925), .B(n11921), .Z(n12485) );
  XNOR U22400 ( .A(n11920), .B(n11916), .Z(n12486) );
  XNOR U22401 ( .A(n11915), .B(n11911), .Z(n12487) );
  XNOR U22402 ( .A(n11910), .B(n11906), .Z(n12488) );
  XNOR U22403 ( .A(n11905), .B(n11901), .Z(n12489) );
  XNOR U22404 ( .A(n11900), .B(n11896), .Z(n12490) );
  XNOR U22405 ( .A(n11895), .B(n11891), .Z(n12491) );
  XNOR U22406 ( .A(n11890), .B(n11886), .Z(n12492) );
  XNOR U22407 ( .A(n11885), .B(n11881), .Z(n12493) );
  XNOR U22408 ( .A(n11880), .B(n11876), .Z(n12494) );
  XNOR U22409 ( .A(n11875), .B(n11871), .Z(n12495) );
  XNOR U22410 ( .A(n11870), .B(n11866), .Z(n12496) );
  XNOR U22411 ( .A(n11865), .B(n11861), .Z(n12497) );
  XNOR U22412 ( .A(n11860), .B(n11856), .Z(n12498) );
  XNOR U22413 ( .A(n11855), .B(n11851), .Z(n12499) );
  XNOR U22414 ( .A(n12500), .B(n11850), .Z(n11851) );
  AND U22415 ( .A(a[0]), .B(b[109]), .Z(n12500) );
  XOR U22416 ( .A(n12501), .B(n11850), .Z(n11852) );
  XNOR U22417 ( .A(n12502), .B(n12503), .Z(n11850) );
  ANDN U22418 ( .B(n12504), .A(n12505), .Z(n12502) );
  AND U22419 ( .A(a[1]), .B(b[108]), .Z(n12501) );
  XNOR U22420 ( .A(n12506), .B(n11855), .Z(n11857) );
  XOR U22421 ( .A(n12507), .B(n12508), .Z(n11855) );
  ANDN U22422 ( .B(n12509), .A(n12510), .Z(n12507) );
  AND U22423 ( .A(a[2]), .B(b[107]), .Z(n12506) );
  XNOR U22424 ( .A(n12511), .B(n11860), .Z(n11862) );
  XOR U22425 ( .A(n12512), .B(n12513), .Z(n11860) );
  ANDN U22426 ( .B(n12514), .A(n12515), .Z(n12512) );
  AND U22427 ( .A(a[3]), .B(b[106]), .Z(n12511) );
  XNOR U22428 ( .A(n12516), .B(n11865), .Z(n11867) );
  XOR U22429 ( .A(n12517), .B(n12518), .Z(n11865) );
  ANDN U22430 ( .B(n12519), .A(n12520), .Z(n12517) );
  AND U22431 ( .A(a[4]), .B(b[105]), .Z(n12516) );
  XNOR U22432 ( .A(n12521), .B(n11870), .Z(n11872) );
  XOR U22433 ( .A(n12522), .B(n12523), .Z(n11870) );
  ANDN U22434 ( .B(n12524), .A(n12525), .Z(n12522) );
  AND U22435 ( .A(a[5]), .B(b[104]), .Z(n12521) );
  XNOR U22436 ( .A(n12526), .B(n11875), .Z(n11877) );
  XOR U22437 ( .A(n12527), .B(n12528), .Z(n11875) );
  ANDN U22438 ( .B(n12529), .A(n12530), .Z(n12527) );
  AND U22439 ( .A(a[6]), .B(b[103]), .Z(n12526) );
  XNOR U22440 ( .A(n12531), .B(n11880), .Z(n11882) );
  XOR U22441 ( .A(n12532), .B(n12533), .Z(n11880) );
  ANDN U22442 ( .B(n12534), .A(n12535), .Z(n12532) );
  AND U22443 ( .A(a[7]), .B(b[102]), .Z(n12531) );
  XNOR U22444 ( .A(n12536), .B(n11885), .Z(n11887) );
  XOR U22445 ( .A(n12537), .B(n12538), .Z(n11885) );
  ANDN U22446 ( .B(n12539), .A(n12540), .Z(n12537) );
  AND U22447 ( .A(a[8]), .B(b[101]), .Z(n12536) );
  XNOR U22448 ( .A(n12541), .B(n11890), .Z(n11892) );
  XOR U22449 ( .A(n12542), .B(n12543), .Z(n11890) );
  ANDN U22450 ( .B(n12544), .A(n12545), .Z(n12542) );
  AND U22451 ( .A(a[9]), .B(b[100]), .Z(n12541) );
  XNOR U22452 ( .A(n12546), .B(n11895), .Z(n11897) );
  XOR U22453 ( .A(n12547), .B(n12548), .Z(n11895) );
  ANDN U22454 ( .B(n12549), .A(n12550), .Z(n12547) );
  AND U22455 ( .A(a[10]), .B(b[99]), .Z(n12546) );
  XNOR U22456 ( .A(n12551), .B(n11900), .Z(n11902) );
  XOR U22457 ( .A(n12552), .B(n12553), .Z(n11900) );
  ANDN U22458 ( .B(n12554), .A(n12555), .Z(n12552) );
  AND U22459 ( .A(a[11]), .B(b[98]), .Z(n12551) );
  XNOR U22460 ( .A(n12556), .B(n11905), .Z(n11907) );
  XOR U22461 ( .A(n12557), .B(n12558), .Z(n11905) );
  ANDN U22462 ( .B(n12559), .A(n12560), .Z(n12557) );
  AND U22463 ( .A(a[12]), .B(b[97]), .Z(n12556) );
  XNOR U22464 ( .A(n12561), .B(n11910), .Z(n11912) );
  XOR U22465 ( .A(n12562), .B(n12563), .Z(n11910) );
  ANDN U22466 ( .B(n12564), .A(n12565), .Z(n12562) );
  AND U22467 ( .A(a[13]), .B(b[96]), .Z(n12561) );
  XNOR U22468 ( .A(n12566), .B(n11915), .Z(n11917) );
  XOR U22469 ( .A(n12567), .B(n12568), .Z(n11915) );
  ANDN U22470 ( .B(n12569), .A(n12570), .Z(n12567) );
  AND U22471 ( .A(a[14]), .B(b[95]), .Z(n12566) );
  XNOR U22472 ( .A(n12571), .B(n11920), .Z(n11922) );
  XOR U22473 ( .A(n12572), .B(n12573), .Z(n11920) );
  ANDN U22474 ( .B(n12574), .A(n12575), .Z(n12572) );
  AND U22475 ( .A(a[15]), .B(b[94]), .Z(n12571) );
  XNOR U22476 ( .A(n12576), .B(n11925), .Z(n11927) );
  XOR U22477 ( .A(n12577), .B(n12578), .Z(n11925) );
  ANDN U22478 ( .B(n12579), .A(n12580), .Z(n12577) );
  AND U22479 ( .A(a[16]), .B(b[93]), .Z(n12576) );
  XNOR U22480 ( .A(n12581), .B(n11930), .Z(n11932) );
  XOR U22481 ( .A(n12582), .B(n12583), .Z(n11930) );
  ANDN U22482 ( .B(n12584), .A(n12585), .Z(n12582) );
  AND U22483 ( .A(a[17]), .B(b[92]), .Z(n12581) );
  XNOR U22484 ( .A(n12586), .B(n11935), .Z(n11937) );
  XOR U22485 ( .A(n12587), .B(n12588), .Z(n11935) );
  ANDN U22486 ( .B(n12589), .A(n12590), .Z(n12587) );
  AND U22487 ( .A(a[18]), .B(b[91]), .Z(n12586) );
  XNOR U22488 ( .A(n12591), .B(n11940), .Z(n11942) );
  XOR U22489 ( .A(n12592), .B(n12593), .Z(n11940) );
  ANDN U22490 ( .B(n12594), .A(n12595), .Z(n12592) );
  AND U22491 ( .A(a[19]), .B(b[90]), .Z(n12591) );
  XNOR U22492 ( .A(n12596), .B(n11945), .Z(n11947) );
  XOR U22493 ( .A(n12597), .B(n12598), .Z(n11945) );
  ANDN U22494 ( .B(n12599), .A(n12600), .Z(n12597) );
  AND U22495 ( .A(a[20]), .B(b[89]), .Z(n12596) );
  XNOR U22496 ( .A(n12601), .B(n11950), .Z(n11952) );
  XOR U22497 ( .A(n12602), .B(n12603), .Z(n11950) );
  ANDN U22498 ( .B(n12604), .A(n12605), .Z(n12602) );
  AND U22499 ( .A(a[21]), .B(b[88]), .Z(n12601) );
  XNOR U22500 ( .A(n12606), .B(n11955), .Z(n11957) );
  XOR U22501 ( .A(n12607), .B(n12608), .Z(n11955) );
  ANDN U22502 ( .B(n12609), .A(n12610), .Z(n12607) );
  AND U22503 ( .A(a[22]), .B(b[87]), .Z(n12606) );
  XNOR U22504 ( .A(n12611), .B(n11960), .Z(n11962) );
  XOR U22505 ( .A(n12612), .B(n12613), .Z(n11960) );
  ANDN U22506 ( .B(n12614), .A(n12615), .Z(n12612) );
  AND U22507 ( .A(a[23]), .B(b[86]), .Z(n12611) );
  XNOR U22508 ( .A(n12616), .B(n11965), .Z(n11967) );
  XOR U22509 ( .A(n12617), .B(n12618), .Z(n11965) );
  ANDN U22510 ( .B(n12619), .A(n12620), .Z(n12617) );
  AND U22511 ( .A(a[24]), .B(b[85]), .Z(n12616) );
  XNOR U22512 ( .A(n12621), .B(n11970), .Z(n11972) );
  XOR U22513 ( .A(n12622), .B(n12623), .Z(n11970) );
  ANDN U22514 ( .B(n12624), .A(n12625), .Z(n12622) );
  AND U22515 ( .A(a[25]), .B(b[84]), .Z(n12621) );
  XNOR U22516 ( .A(n12626), .B(n11975), .Z(n11977) );
  XOR U22517 ( .A(n12627), .B(n12628), .Z(n11975) );
  ANDN U22518 ( .B(n12629), .A(n12630), .Z(n12627) );
  AND U22519 ( .A(a[26]), .B(b[83]), .Z(n12626) );
  XNOR U22520 ( .A(n12631), .B(n11980), .Z(n11982) );
  XOR U22521 ( .A(n12632), .B(n12633), .Z(n11980) );
  ANDN U22522 ( .B(n12634), .A(n12635), .Z(n12632) );
  AND U22523 ( .A(a[27]), .B(b[82]), .Z(n12631) );
  XNOR U22524 ( .A(n12636), .B(n11985), .Z(n11987) );
  XOR U22525 ( .A(n12637), .B(n12638), .Z(n11985) );
  ANDN U22526 ( .B(n12639), .A(n12640), .Z(n12637) );
  AND U22527 ( .A(a[28]), .B(b[81]), .Z(n12636) );
  XNOR U22528 ( .A(n12641), .B(n11990), .Z(n11992) );
  XOR U22529 ( .A(n12642), .B(n12643), .Z(n11990) );
  ANDN U22530 ( .B(n12644), .A(n12645), .Z(n12642) );
  AND U22531 ( .A(a[29]), .B(b[80]), .Z(n12641) );
  XNOR U22532 ( .A(n12646), .B(n11995), .Z(n11997) );
  XOR U22533 ( .A(n12647), .B(n12648), .Z(n11995) );
  ANDN U22534 ( .B(n12649), .A(n12650), .Z(n12647) );
  AND U22535 ( .A(a[30]), .B(b[79]), .Z(n12646) );
  XNOR U22536 ( .A(n12651), .B(n12000), .Z(n12002) );
  XOR U22537 ( .A(n12652), .B(n12653), .Z(n12000) );
  ANDN U22538 ( .B(n12654), .A(n12655), .Z(n12652) );
  AND U22539 ( .A(a[31]), .B(b[78]), .Z(n12651) );
  XNOR U22540 ( .A(n12656), .B(n12005), .Z(n12007) );
  XOR U22541 ( .A(n12657), .B(n12658), .Z(n12005) );
  ANDN U22542 ( .B(n12659), .A(n12660), .Z(n12657) );
  AND U22543 ( .A(a[32]), .B(b[77]), .Z(n12656) );
  XNOR U22544 ( .A(n12661), .B(n12010), .Z(n12012) );
  XOR U22545 ( .A(n12662), .B(n12663), .Z(n12010) );
  ANDN U22546 ( .B(n12664), .A(n12665), .Z(n12662) );
  AND U22547 ( .A(a[33]), .B(b[76]), .Z(n12661) );
  XNOR U22548 ( .A(n12666), .B(n12015), .Z(n12017) );
  XOR U22549 ( .A(n12667), .B(n12668), .Z(n12015) );
  ANDN U22550 ( .B(n12669), .A(n12670), .Z(n12667) );
  AND U22551 ( .A(a[34]), .B(b[75]), .Z(n12666) );
  XNOR U22552 ( .A(n12671), .B(n12020), .Z(n12022) );
  XOR U22553 ( .A(n12672), .B(n12673), .Z(n12020) );
  ANDN U22554 ( .B(n12674), .A(n12675), .Z(n12672) );
  AND U22555 ( .A(a[35]), .B(b[74]), .Z(n12671) );
  XNOR U22556 ( .A(n12676), .B(n12025), .Z(n12027) );
  XOR U22557 ( .A(n12677), .B(n12678), .Z(n12025) );
  ANDN U22558 ( .B(n12679), .A(n12680), .Z(n12677) );
  AND U22559 ( .A(a[36]), .B(b[73]), .Z(n12676) );
  XNOR U22560 ( .A(n12681), .B(n12030), .Z(n12032) );
  XOR U22561 ( .A(n12682), .B(n12683), .Z(n12030) );
  ANDN U22562 ( .B(n12684), .A(n12685), .Z(n12682) );
  AND U22563 ( .A(a[37]), .B(b[72]), .Z(n12681) );
  XNOR U22564 ( .A(n12686), .B(n12035), .Z(n12037) );
  XOR U22565 ( .A(n12687), .B(n12688), .Z(n12035) );
  ANDN U22566 ( .B(n12689), .A(n12690), .Z(n12687) );
  AND U22567 ( .A(a[38]), .B(b[71]), .Z(n12686) );
  XNOR U22568 ( .A(n12691), .B(n12040), .Z(n12042) );
  XOR U22569 ( .A(n12692), .B(n12693), .Z(n12040) );
  ANDN U22570 ( .B(n12694), .A(n12695), .Z(n12692) );
  AND U22571 ( .A(a[39]), .B(b[70]), .Z(n12691) );
  XNOR U22572 ( .A(n12696), .B(n12045), .Z(n12047) );
  XOR U22573 ( .A(n12697), .B(n12698), .Z(n12045) );
  ANDN U22574 ( .B(n12699), .A(n12700), .Z(n12697) );
  AND U22575 ( .A(a[40]), .B(b[69]), .Z(n12696) );
  XNOR U22576 ( .A(n12701), .B(n12050), .Z(n12052) );
  XOR U22577 ( .A(n12702), .B(n12703), .Z(n12050) );
  ANDN U22578 ( .B(n12704), .A(n12705), .Z(n12702) );
  AND U22579 ( .A(a[41]), .B(b[68]), .Z(n12701) );
  XNOR U22580 ( .A(n12706), .B(n12055), .Z(n12057) );
  XOR U22581 ( .A(n12707), .B(n12708), .Z(n12055) );
  ANDN U22582 ( .B(n12709), .A(n12710), .Z(n12707) );
  AND U22583 ( .A(a[42]), .B(b[67]), .Z(n12706) );
  XNOR U22584 ( .A(n12711), .B(n12060), .Z(n12062) );
  XOR U22585 ( .A(n12712), .B(n12713), .Z(n12060) );
  ANDN U22586 ( .B(n12714), .A(n12715), .Z(n12712) );
  AND U22587 ( .A(a[43]), .B(b[66]), .Z(n12711) );
  XNOR U22588 ( .A(n12716), .B(n12065), .Z(n12067) );
  XOR U22589 ( .A(n12717), .B(n12718), .Z(n12065) );
  ANDN U22590 ( .B(n12719), .A(n12720), .Z(n12717) );
  AND U22591 ( .A(a[44]), .B(b[65]), .Z(n12716) );
  XNOR U22592 ( .A(n12721), .B(n12070), .Z(n12072) );
  XOR U22593 ( .A(n12722), .B(n12723), .Z(n12070) );
  ANDN U22594 ( .B(n12724), .A(n12725), .Z(n12722) );
  AND U22595 ( .A(a[45]), .B(b[64]), .Z(n12721) );
  XNOR U22596 ( .A(n12726), .B(n12075), .Z(n12077) );
  XOR U22597 ( .A(n12727), .B(n12728), .Z(n12075) );
  ANDN U22598 ( .B(n12729), .A(n12730), .Z(n12727) );
  AND U22599 ( .A(a[46]), .B(b[63]), .Z(n12726) );
  XNOR U22600 ( .A(n12731), .B(n12080), .Z(n12082) );
  XOR U22601 ( .A(n12732), .B(n12733), .Z(n12080) );
  ANDN U22602 ( .B(n12734), .A(n12735), .Z(n12732) );
  AND U22603 ( .A(a[47]), .B(b[62]), .Z(n12731) );
  XNOR U22604 ( .A(n12736), .B(n12085), .Z(n12087) );
  XOR U22605 ( .A(n12737), .B(n12738), .Z(n12085) );
  ANDN U22606 ( .B(n12739), .A(n12740), .Z(n12737) );
  AND U22607 ( .A(a[48]), .B(b[61]), .Z(n12736) );
  XNOR U22608 ( .A(n12741), .B(n12090), .Z(n12092) );
  XOR U22609 ( .A(n12742), .B(n12743), .Z(n12090) );
  ANDN U22610 ( .B(n12744), .A(n12745), .Z(n12742) );
  AND U22611 ( .A(a[49]), .B(b[60]), .Z(n12741) );
  XNOR U22612 ( .A(n12746), .B(n12095), .Z(n12097) );
  XOR U22613 ( .A(n12747), .B(n12748), .Z(n12095) );
  ANDN U22614 ( .B(n12749), .A(n12750), .Z(n12747) );
  AND U22615 ( .A(a[50]), .B(b[59]), .Z(n12746) );
  XNOR U22616 ( .A(n12751), .B(n12100), .Z(n12102) );
  XOR U22617 ( .A(n12752), .B(n12753), .Z(n12100) );
  ANDN U22618 ( .B(n12754), .A(n12755), .Z(n12752) );
  AND U22619 ( .A(a[51]), .B(b[58]), .Z(n12751) );
  XNOR U22620 ( .A(n12756), .B(n12105), .Z(n12107) );
  XOR U22621 ( .A(n12757), .B(n12758), .Z(n12105) );
  ANDN U22622 ( .B(n12759), .A(n12760), .Z(n12757) );
  AND U22623 ( .A(a[52]), .B(b[57]), .Z(n12756) );
  XNOR U22624 ( .A(n12761), .B(n12110), .Z(n12112) );
  XOR U22625 ( .A(n12762), .B(n12763), .Z(n12110) );
  ANDN U22626 ( .B(n12764), .A(n12765), .Z(n12762) );
  AND U22627 ( .A(a[53]), .B(b[56]), .Z(n12761) );
  XNOR U22628 ( .A(n12766), .B(n12115), .Z(n12117) );
  XOR U22629 ( .A(n12767), .B(n12768), .Z(n12115) );
  ANDN U22630 ( .B(n12769), .A(n12770), .Z(n12767) );
  AND U22631 ( .A(a[54]), .B(b[55]), .Z(n12766) );
  XNOR U22632 ( .A(n12771), .B(n12120), .Z(n12122) );
  XOR U22633 ( .A(n12772), .B(n12773), .Z(n12120) );
  ANDN U22634 ( .B(n12774), .A(n12775), .Z(n12772) );
  AND U22635 ( .A(a[55]), .B(b[54]), .Z(n12771) );
  XNOR U22636 ( .A(n12776), .B(n12125), .Z(n12127) );
  XOR U22637 ( .A(n12777), .B(n12778), .Z(n12125) );
  ANDN U22638 ( .B(n12779), .A(n12780), .Z(n12777) );
  AND U22639 ( .A(a[56]), .B(b[53]), .Z(n12776) );
  XNOR U22640 ( .A(n12781), .B(n12130), .Z(n12132) );
  XOR U22641 ( .A(n12782), .B(n12783), .Z(n12130) );
  ANDN U22642 ( .B(n12784), .A(n12785), .Z(n12782) );
  AND U22643 ( .A(a[57]), .B(b[52]), .Z(n12781) );
  XNOR U22644 ( .A(n12786), .B(n12135), .Z(n12137) );
  XOR U22645 ( .A(n12787), .B(n12788), .Z(n12135) );
  ANDN U22646 ( .B(n12789), .A(n12790), .Z(n12787) );
  AND U22647 ( .A(a[58]), .B(b[51]), .Z(n12786) );
  XNOR U22648 ( .A(n12791), .B(n12140), .Z(n12142) );
  XOR U22649 ( .A(n12792), .B(n12793), .Z(n12140) );
  ANDN U22650 ( .B(n12794), .A(n12795), .Z(n12792) );
  AND U22651 ( .A(a[59]), .B(b[50]), .Z(n12791) );
  XNOR U22652 ( .A(n12796), .B(n12145), .Z(n12147) );
  XOR U22653 ( .A(n12797), .B(n12798), .Z(n12145) );
  ANDN U22654 ( .B(n12799), .A(n12800), .Z(n12797) );
  AND U22655 ( .A(a[60]), .B(b[49]), .Z(n12796) );
  XNOR U22656 ( .A(n12801), .B(n12150), .Z(n12152) );
  XOR U22657 ( .A(n12802), .B(n12803), .Z(n12150) );
  ANDN U22658 ( .B(n12804), .A(n12805), .Z(n12802) );
  AND U22659 ( .A(a[61]), .B(b[48]), .Z(n12801) );
  XNOR U22660 ( .A(n12806), .B(n12155), .Z(n12157) );
  XOR U22661 ( .A(n12807), .B(n12808), .Z(n12155) );
  ANDN U22662 ( .B(n12809), .A(n12810), .Z(n12807) );
  AND U22663 ( .A(a[62]), .B(b[47]), .Z(n12806) );
  XNOR U22664 ( .A(n12811), .B(n12160), .Z(n12162) );
  XOR U22665 ( .A(n12812), .B(n12813), .Z(n12160) );
  ANDN U22666 ( .B(n12814), .A(n12815), .Z(n12812) );
  AND U22667 ( .A(a[63]), .B(b[46]), .Z(n12811) );
  XNOR U22668 ( .A(n12816), .B(n12165), .Z(n12167) );
  XOR U22669 ( .A(n12817), .B(n12818), .Z(n12165) );
  ANDN U22670 ( .B(n12819), .A(n12820), .Z(n12817) );
  AND U22671 ( .A(a[64]), .B(b[45]), .Z(n12816) );
  XNOR U22672 ( .A(n12821), .B(n12170), .Z(n12172) );
  XOR U22673 ( .A(n12822), .B(n12823), .Z(n12170) );
  ANDN U22674 ( .B(n12824), .A(n12825), .Z(n12822) );
  AND U22675 ( .A(a[65]), .B(b[44]), .Z(n12821) );
  XNOR U22676 ( .A(n12826), .B(n12175), .Z(n12177) );
  XOR U22677 ( .A(n12827), .B(n12828), .Z(n12175) );
  ANDN U22678 ( .B(n12829), .A(n12830), .Z(n12827) );
  AND U22679 ( .A(a[66]), .B(b[43]), .Z(n12826) );
  XNOR U22680 ( .A(n12831), .B(n12180), .Z(n12182) );
  XOR U22681 ( .A(n12832), .B(n12833), .Z(n12180) );
  ANDN U22682 ( .B(n12834), .A(n12835), .Z(n12832) );
  AND U22683 ( .A(a[67]), .B(b[42]), .Z(n12831) );
  XNOR U22684 ( .A(n12836), .B(n12185), .Z(n12187) );
  XOR U22685 ( .A(n12837), .B(n12838), .Z(n12185) );
  ANDN U22686 ( .B(n12839), .A(n12840), .Z(n12837) );
  AND U22687 ( .A(a[68]), .B(b[41]), .Z(n12836) );
  XNOR U22688 ( .A(n12841), .B(n12190), .Z(n12192) );
  XOR U22689 ( .A(n12842), .B(n12843), .Z(n12190) );
  ANDN U22690 ( .B(n12844), .A(n12845), .Z(n12842) );
  AND U22691 ( .A(a[69]), .B(b[40]), .Z(n12841) );
  XNOR U22692 ( .A(n12846), .B(n12195), .Z(n12197) );
  XOR U22693 ( .A(n12847), .B(n12848), .Z(n12195) );
  ANDN U22694 ( .B(n12849), .A(n12850), .Z(n12847) );
  AND U22695 ( .A(a[70]), .B(b[39]), .Z(n12846) );
  XNOR U22696 ( .A(n12851), .B(n12200), .Z(n12202) );
  XOR U22697 ( .A(n12852), .B(n12853), .Z(n12200) );
  ANDN U22698 ( .B(n12854), .A(n12855), .Z(n12852) );
  AND U22699 ( .A(a[71]), .B(b[38]), .Z(n12851) );
  XNOR U22700 ( .A(n12856), .B(n12205), .Z(n12207) );
  XOR U22701 ( .A(n12857), .B(n12858), .Z(n12205) );
  ANDN U22702 ( .B(n12859), .A(n12860), .Z(n12857) );
  AND U22703 ( .A(a[72]), .B(b[37]), .Z(n12856) );
  XNOR U22704 ( .A(n12861), .B(n12210), .Z(n12212) );
  XOR U22705 ( .A(n12862), .B(n12863), .Z(n12210) );
  ANDN U22706 ( .B(n12864), .A(n12865), .Z(n12862) );
  AND U22707 ( .A(a[73]), .B(b[36]), .Z(n12861) );
  XNOR U22708 ( .A(n12866), .B(n12215), .Z(n12217) );
  XOR U22709 ( .A(n12867), .B(n12868), .Z(n12215) );
  ANDN U22710 ( .B(n12869), .A(n12870), .Z(n12867) );
  AND U22711 ( .A(a[74]), .B(b[35]), .Z(n12866) );
  XNOR U22712 ( .A(n12871), .B(n12220), .Z(n12222) );
  XOR U22713 ( .A(n12872), .B(n12873), .Z(n12220) );
  ANDN U22714 ( .B(n12874), .A(n12875), .Z(n12872) );
  AND U22715 ( .A(a[75]), .B(b[34]), .Z(n12871) );
  XNOR U22716 ( .A(n12876), .B(n12225), .Z(n12227) );
  XOR U22717 ( .A(n12877), .B(n12878), .Z(n12225) );
  ANDN U22718 ( .B(n12879), .A(n12880), .Z(n12877) );
  AND U22719 ( .A(a[76]), .B(b[33]), .Z(n12876) );
  XNOR U22720 ( .A(n12881), .B(n12230), .Z(n12232) );
  XOR U22721 ( .A(n12882), .B(n12883), .Z(n12230) );
  ANDN U22722 ( .B(n12884), .A(n12885), .Z(n12882) );
  AND U22723 ( .A(a[77]), .B(b[32]), .Z(n12881) );
  XNOR U22724 ( .A(n12886), .B(n12235), .Z(n12237) );
  XOR U22725 ( .A(n12887), .B(n12888), .Z(n12235) );
  ANDN U22726 ( .B(n12889), .A(n12890), .Z(n12887) );
  AND U22727 ( .A(a[78]), .B(b[31]), .Z(n12886) );
  XNOR U22728 ( .A(n12891), .B(n12240), .Z(n12242) );
  XOR U22729 ( .A(n12892), .B(n12893), .Z(n12240) );
  ANDN U22730 ( .B(n12894), .A(n12895), .Z(n12892) );
  AND U22731 ( .A(a[79]), .B(b[30]), .Z(n12891) );
  XNOR U22732 ( .A(n12896), .B(n12245), .Z(n12247) );
  XOR U22733 ( .A(n12897), .B(n12898), .Z(n12245) );
  ANDN U22734 ( .B(n12899), .A(n12900), .Z(n12897) );
  AND U22735 ( .A(a[80]), .B(b[29]), .Z(n12896) );
  XNOR U22736 ( .A(n12901), .B(n12250), .Z(n12252) );
  XOR U22737 ( .A(n12902), .B(n12903), .Z(n12250) );
  ANDN U22738 ( .B(n12904), .A(n12905), .Z(n12902) );
  AND U22739 ( .A(a[81]), .B(b[28]), .Z(n12901) );
  XNOR U22740 ( .A(n12906), .B(n12255), .Z(n12257) );
  XOR U22741 ( .A(n12907), .B(n12908), .Z(n12255) );
  ANDN U22742 ( .B(n12909), .A(n12910), .Z(n12907) );
  AND U22743 ( .A(a[82]), .B(b[27]), .Z(n12906) );
  XNOR U22744 ( .A(n12911), .B(n12260), .Z(n12262) );
  XOR U22745 ( .A(n12912), .B(n12913), .Z(n12260) );
  ANDN U22746 ( .B(n12914), .A(n12915), .Z(n12912) );
  AND U22747 ( .A(a[83]), .B(b[26]), .Z(n12911) );
  XNOR U22748 ( .A(n12916), .B(n12265), .Z(n12267) );
  XOR U22749 ( .A(n12917), .B(n12918), .Z(n12265) );
  ANDN U22750 ( .B(n12919), .A(n12920), .Z(n12917) );
  AND U22751 ( .A(a[84]), .B(b[25]), .Z(n12916) );
  XNOR U22752 ( .A(n12921), .B(n12270), .Z(n12272) );
  XOR U22753 ( .A(n12922), .B(n12923), .Z(n12270) );
  ANDN U22754 ( .B(n12924), .A(n12925), .Z(n12922) );
  AND U22755 ( .A(a[85]), .B(b[24]), .Z(n12921) );
  XNOR U22756 ( .A(n12926), .B(n12275), .Z(n12277) );
  XOR U22757 ( .A(n12927), .B(n12928), .Z(n12275) );
  ANDN U22758 ( .B(n12929), .A(n12930), .Z(n12927) );
  AND U22759 ( .A(a[86]), .B(b[23]), .Z(n12926) );
  XNOR U22760 ( .A(n12931), .B(n12280), .Z(n12282) );
  XOR U22761 ( .A(n12932), .B(n12933), .Z(n12280) );
  ANDN U22762 ( .B(n12934), .A(n12935), .Z(n12932) );
  AND U22763 ( .A(a[87]), .B(b[22]), .Z(n12931) );
  XNOR U22764 ( .A(n12936), .B(n12285), .Z(n12287) );
  XOR U22765 ( .A(n12937), .B(n12938), .Z(n12285) );
  ANDN U22766 ( .B(n12939), .A(n12940), .Z(n12937) );
  AND U22767 ( .A(a[88]), .B(b[21]), .Z(n12936) );
  XNOR U22768 ( .A(n12941), .B(n12290), .Z(n12292) );
  XOR U22769 ( .A(n12942), .B(n12943), .Z(n12290) );
  ANDN U22770 ( .B(n12944), .A(n12945), .Z(n12942) );
  AND U22771 ( .A(a[89]), .B(b[20]), .Z(n12941) );
  XNOR U22772 ( .A(n12946), .B(n12295), .Z(n12297) );
  XOR U22773 ( .A(n12947), .B(n12948), .Z(n12295) );
  ANDN U22774 ( .B(n12949), .A(n12950), .Z(n12947) );
  AND U22775 ( .A(a[90]), .B(b[19]), .Z(n12946) );
  XNOR U22776 ( .A(n12951), .B(n12300), .Z(n12302) );
  XOR U22777 ( .A(n12952), .B(n12953), .Z(n12300) );
  ANDN U22778 ( .B(n12954), .A(n12955), .Z(n12952) );
  AND U22779 ( .A(a[91]), .B(b[18]), .Z(n12951) );
  XNOR U22780 ( .A(n12956), .B(n12305), .Z(n12307) );
  XOR U22781 ( .A(n12957), .B(n12958), .Z(n12305) );
  ANDN U22782 ( .B(n12959), .A(n12960), .Z(n12957) );
  AND U22783 ( .A(a[92]), .B(b[17]), .Z(n12956) );
  XNOR U22784 ( .A(n12961), .B(n12310), .Z(n12312) );
  XOR U22785 ( .A(n12962), .B(n12963), .Z(n12310) );
  ANDN U22786 ( .B(n12964), .A(n12965), .Z(n12962) );
  AND U22787 ( .A(a[93]), .B(b[16]), .Z(n12961) );
  XNOR U22788 ( .A(n12966), .B(n12315), .Z(n12317) );
  XOR U22789 ( .A(n12967), .B(n12968), .Z(n12315) );
  ANDN U22790 ( .B(n12969), .A(n12970), .Z(n12967) );
  AND U22791 ( .A(a[94]), .B(b[15]), .Z(n12966) );
  XNOR U22792 ( .A(n12971), .B(n12320), .Z(n12322) );
  XOR U22793 ( .A(n12972), .B(n12973), .Z(n12320) );
  ANDN U22794 ( .B(n12974), .A(n12975), .Z(n12972) );
  AND U22795 ( .A(a[95]), .B(b[14]), .Z(n12971) );
  XNOR U22796 ( .A(n12976), .B(n12325), .Z(n12327) );
  XOR U22797 ( .A(n12977), .B(n12978), .Z(n12325) );
  ANDN U22798 ( .B(n12979), .A(n12980), .Z(n12977) );
  AND U22799 ( .A(a[96]), .B(b[13]), .Z(n12976) );
  XNOR U22800 ( .A(n12981), .B(n12330), .Z(n12332) );
  XOR U22801 ( .A(n12982), .B(n12983), .Z(n12330) );
  ANDN U22802 ( .B(n12984), .A(n12985), .Z(n12982) );
  AND U22803 ( .A(a[97]), .B(b[12]), .Z(n12981) );
  XNOR U22804 ( .A(n12986), .B(n12335), .Z(n12337) );
  XOR U22805 ( .A(n12987), .B(n12988), .Z(n12335) );
  ANDN U22806 ( .B(n12989), .A(n12990), .Z(n12987) );
  AND U22807 ( .A(a[98]), .B(b[11]), .Z(n12986) );
  XNOR U22808 ( .A(n12991), .B(n12340), .Z(n12342) );
  XOR U22809 ( .A(n12992), .B(n12993), .Z(n12340) );
  ANDN U22810 ( .B(n12994), .A(n12995), .Z(n12992) );
  AND U22811 ( .A(a[99]), .B(b[10]), .Z(n12991) );
  XNOR U22812 ( .A(n12996), .B(n12345), .Z(n12347) );
  XOR U22813 ( .A(n12997), .B(n12998), .Z(n12345) );
  ANDN U22814 ( .B(n12999), .A(n13000), .Z(n12997) );
  AND U22815 ( .A(b[9]), .B(a[100]), .Z(n12996) );
  XNOR U22816 ( .A(n13001), .B(n12350), .Z(n12352) );
  XOR U22817 ( .A(n13002), .B(n13003), .Z(n12350) );
  ANDN U22818 ( .B(n13004), .A(n13005), .Z(n13002) );
  AND U22819 ( .A(b[8]), .B(a[101]), .Z(n13001) );
  XNOR U22820 ( .A(n13006), .B(n12355), .Z(n12357) );
  XOR U22821 ( .A(n13007), .B(n13008), .Z(n12355) );
  ANDN U22822 ( .B(n13009), .A(n13010), .Z(n13007) );
  AND U22823 ( .A(b[7]), .B(a[102]), .Z(n13006) );
  XNOR U22824 ( .A(n13011), .B(n12360), .Z(n12362) );
  XOR U22825 ( .A(n13012), .B(n13013), .Z(n12360) );
  ANDN U22826 ( .B(n13014), .A(n13015), .Z(n13012) );
  AND U22827 ( .A(b[6]), .B(a[103]), .Z(n13011) );
  XNOR U22828 ( .A(n13016), .B(n12365), .Z(n12367) );
  XOR U22829 ( .A(n13017), .B(n13018), .Z(n12365) );
  ANDN U22830 ( .B(n13019), .A(n13020), .Z(n13017) );
  AND U22831 ( .A(b[5]), .B(a[104]), .Z(n13016) );
  XNOR U22832 ( .A(n13021), .B(n12370), .Z(n12372) );
  XOR U22833 ( .A(n13022), .B(n13023), .Z(n12370) );
  ANDN U22834 ( .B(n13024), .A(n13025), .Z(n13022) );
  AND U22835 ( .A(b[4]), .B(a[105]), .Z(n13021) );
  XNOR U22836 ( .A(n13026), .B(n13027), .Z(n12384) );
  NANDN U22837 ( .A(n13028), .B(n13029), .Z(n13027) );
  XNOR U22838 ( .A(n13030), .B(n12375), .Z(n12377) );
  XNOR U22839 ( .A(n13031), .B(n13032), .Z(n12375) );
  AND U22840 ( .A(n13033), .B(n13034), .Z(n13031) );
  AND U22841 ( .A(b[3]), .B(a[106]), .Z(n13030) );
  NAND U22842 ( .A(a[109]), .B(b[0]), .Z(n11738) );
  XNOR U22843 ( .A(n12392), .B(n12393), .Z(c[108]) );
  XNOR U22844 ( .A(n13028), .B(n13029), .Z(n12393) );
  XOR U22845 ( .A(n13026), .B(n13035), .Z(n13029) );
  NAND U22846 ( .A(b[1]), .B(a[107]), .Z(n13035) );
  XOR U22847 ( .A(n13034), .B(n13036), .Z(n13028) );
  XOR U22848 ( .A(n13026), .B(n13033), .Z(n13036) );
  XNOR U22849 ( .A(n13037), .B(n13032), .Z(n13033) );
  AND U22850 ( .A(b[2]), .B(a[106]), .Z(n13037) );
  NANDN U22851 ( .A(n13038), .B(n13039), .Z(n13026) );
  XOR U22852 ( .A(n13032), .B(n13024), .Z(n13040) );
  XNOR U22853 ( .A(n13023), .B(n13019), .Z(n13041) );
  XNOR U22854 ( .A(n13018), .B(n13014), .Z(n13042) );
  XNOR U22855 ( .A(n13013), .B(n13009), .Z(n13043) );
  XNOR U22856 ( .A(n13008), .B(n13004), .Z(n13044) );
  XNOR U22857 ( .A(n13003), .B(n12999), .Z(n13045) );
  XNOR U22858 ( .A(n12998), .B(n12994), .Z(n13046) );
  XNOR U22859 ( .A(n12993), .B(n12989), .Z(n13047) );
  XNOR U22860 ( .A(n12988), .B(n12984), .Z(n13048) );
  XNOR U22861 ( .A(n12983), .B(n12979), .Z(n13049) );
  XNOR U22862 ( .A(n12978), .B(n12974), .Z(n13050) );
  XNOR U22863 ( .A(n12973), .B(n12969), .Z(n13051) );
  XNOR U22864 ( .A(n12968), .B(n12964), .Z(n13052) );
  XNOR U22865 ( .A(n12963), .B(n12959), .Z(n13053) );
  XNOR U22866 ( .A(n12958), .B(n12954), .Z(n13054) );
  XNOR U22867 ( .A(n12953), .B(n12949), .Z(n13055) );
  XNOR U22868 ( .A(n12948), .B(n12944), .Z(n13056) );
  XNOR U22869 ( .A(n12943), .B(n12939), .Z(n13057) );
  XNOR U22870 ( .A(n12938), .B(n12934), .Z(n13058) );
  XNOR U22871 ( .A(n12933), .B(n12929), .Z(n13059) );
  XNOR U22872 ( .A(n12928), .B(n12924), .Z(n13060) );
  XNOR U22873 ( .A(n12923), .B(n12919), .Z(n13061) );
  XNOR U22874 ( .A(n12918), .B(n12914), .Z(n13062) );
  XNOR U22875 ( .A(n12913), .B(n12909), .Z(n13063) );
  XNOR U22876 ( .A(n12908), .B(n12904), .Z(n13064) );
  XNOR U22877 ( .A(n12903), .B(n12899), .Z(n13065) );
  XNOR U22878 ( .A(n12898), .B(n12894), .Z(n13066) );
  XNOR U22879 ( .A(n12893), .B(n12889), .Z(n13067) );
  XNOR U22880 ( .A(n12888), .B(n12884), .Z(n13068) );
  XNOR U22881 ( .A(n12883), .B(n12879), .Z(n13069) );
  XNOR U22882 ( .A(n12878), .B(n12874), .Z(n13070) );
  XNOR U22883 ( .A(n12873), .B(n12869), .Z(n13071) );
  XNOR U22884 ( .A(n12868), .B(n12864), .Z(n13072) );
  XNOR U22885 ( .A(n12863), .B(n12859), .Z(n13073) );
  XNOR U22886 ( .A(n12858), .B(n12854), .Z(n13074) );
  XNOR U22887 ( .A(n12853), .B(n12849), .Z(n13075) );
  XNOR U22888 ( .A(n12848), .B(n12844), .Z(n13076) );
  XNOR U22889 ( .A(n12843), .B(n12839), .Z(n13077) );
  XNOR U22890 ( .A(n12838), .B(n12834), .Z(n13078) );
  XNOR U22891 ( .A(n12833), .B(n12829), .Z(n13079) );
  XNOR U22892 ( .A(n12828), .B(n12824), .Z(n13080) );
  XNOR U22893 ( .A(n12823), .B(n12819), .Z(n13081) );
  XNOR U22894 ( .A(n12818), .B(n12814), .Z(n13082) );
  XNOR U22895 ( .A(n12813), .B(n12809), .Z(n13083) );
  XNOR U22896 ( .A(n12808), .B(n12804), .Z(n13084) );
  XNOR U22897 ( .A(n12803), .B(n12799), .Z(n13085) );
  XNOR U22898 ( .A(n12798), .B(n12794), .Z(n13086) );
  XNOR U22899 ( .A(n12793), .B(n12789), .Z(n13087) );
  XNOR U22900 ( .A(n12788), .B(n12784), .Z(n13088) );
  XNOR U22901 ( .A(n12783), .B(n12779), .Z(n13089) );
  XNOR U22902 ( .A(n12778), .B(n12774), .Z(n13090) );
  XNOR U22903 ( .A(n12773), .B(n12769), .Z(n13091) );
  XNOR U22904 ( .A(n12768), .B(n12764), .Z(n13092) );
  XNOR U22905 ( .A(n12763), .B(n12759), .Z(n13093) );
  XNOR U22906 ( .A(n12758), .B(n12754), .Z(n13094) );
  XNOR U22907 ( .A(n12753), .B(n12749), .Z(n13095) );
  XNOR U22908 ( .A(n12748), .B(n12744), .Z(n13096) );
  XNOR U22909 ( .A(n12743), .B(n12739), .Z(n13097) );
  XNOR U22910 ( .A(n12738), .B(n12734), .Z(n13098) );
  XNOR U22911 ( .A(n12733), .B(n12729), .Z(n13099) );
  XNOR U22912 ( .A(n12728), .B(n12724), .Z(n13100) );
  XNOR U22913 ( .A(n12723), .B(n12719), .Z(n13101) );
  XNOR U22914 ( .A(n12718), .B(n12714), .Z(n13102) );
  XNOR U22915 ( .A(n12713), .B(n12709), .Z(n13103) );
  XNOR U22916 ( .A(n12708), .B(n12704), .Z(n13104) );
  XNOR U22917 ( .A(n12703), .B(n12699), .Z(n13105) );
  XNOR U22918 ( .A(n12698), .B(n12694), .Z(n13106) );
  XNOR U22919 ( .A(n12693), .B(n12689), .Z(n13107) );
  XNOR U22920 ( .A(n12688), .B(n12684), .Z(n13108) );
  XNOR U22921 ( .A(n12683), .B(n12679), .Z(n13109) );
  XNOR U22922 ( .A(n12678), .B(n12674), .Z(n13110) );
  XNOR U22923 ( .A(n12673), .B(n12669), .Z(n13111) );
  XNOR U22924 ( .A(n12668), .B(n12664), .Z(n13112) );
  XNOR U22925 ( .A(n12663), .B(n12659), .Z(n13113) );
  XNOR U22926 ( .A(n12658), .B(n12654), .Z(n13114) );
  XNOR U22927 ( .A(n12653), .B(n12649), .Z(n13115) );
  XNOR U22928 ( .A(n12648), .B(n12644), .Z(n13116) );
  XNOR U22929 ( .A(n12643), .B(n12639), .Z(n13117) );
  XNOR U22930 ( .A(n12638), .B(n12634), .Z(n13118) );
  XNOR U22931 ( .A(n12633), .B(n12629), .Z(n13119) );
  XNOR U22932 ( .A(n12628), .B(n12624), .Z(n13120) );
  XNOR U22933 ( .A(n12623), .B(n12619), .Z(n13121) );
  XNOR U22934 ( .A(n12618), .B(n12614), .Z(n13122) );
  XNOR U22935 ( .A(n12613), .B(n12609), .Z(n13123) );
  XNOR U22936 ( .A(n12608), .B(n12604), .Z(n13124) );
  XNOR U22937 ( .A(n12603), .B(n12599), .Z(n13125) );
  XNOR U22938 ( .A(n12598), .B(n12594), .Z(n13126) );
  XNOR U22939 ( .A(n12593), .B(n12589), .Z(n13127) );
  XNOR U22940 ( .A(n12588), .B(n12584), .Z(n13128) );
  XNOR U22941 ( .A(n12583), .B(n12579), .Z(n13129) );
  XNOR U22942 ( .A(n12578), .B(n12574), .Z(n13130) );
  XNOR U22943 ( .A(n12573), .B(n12569), .Z(n13131) );
  XNOR U22944 ( .A(n12568), .B(n12564), .Z(n13132) );
  XNOR U22945 ( .A(n12563), .B(n12559), .Z(n13133) );
  XNOR U22946 ( .A(n12558), .B(n12554), .Z(n13134) );
  XNOR U22947 ( .A(n12553), .B(n12549), .Z(n13135) );
  XNOR U22948 ( .A(n12548), .B(n12544), .Z(n13136) );
  XNOR U22949 ( .A(n12543), .B(n12539), .Z(n13137) );
  XNOR U22950 ( .A(n12538), .B(n12534), .Z(n13138) );
  XNOR U22951 ( .A(n12533), .B(n12529), .Z(n13139) );
  XNOR U22952 ( .A(n12528), .B(n12524), .Z(n13140) );
  XNOR U22953 ( .A(n12523), .B(n12519), .Z(n13141) );
  XNOR U22954 ( .A(n12518), .B(n12514), .Z(n13142) );
  XNOR U22955 ( .A(n12513), .B(n12509), .Z(n13143) );
  XNOR U22956 ( .A(n12508), .B(n12504), .Z(n13144) );
  XOR U22957 ( .A(n13145), .B(n12503), .Z(n12504) );
  AND U22958 ( .A(a[0]), .B(b[108]), .Z(n13145) );
  XNOR U22959 ( .A(n13146), .B(n12503), .Z(n12505) );
  XNOR U22960 ( .A(n13147), .B(n13148), .Z(n12503) );
  ANDN U22961 ( .B(n13149), .A(n13150), .Z(n13147) );
  AND U22962 ( .A(a[1]), .B(b[107]), .Z(n13146) );
  XNOR U22963 ( .A(n13151), .B(n12508), .Z(n12510) );
  XOR U22964 ( .A(n13152), .B(n13153), .Z(n12508) );
  ANDN U22965 ( .B(n13154), .A(n13155), .Z(n13152) );
  AND U22966 ( .A(a[2]), .B(b[106]), .Z(n13151) );
  XNOR U22967 ( .A(n13156), .B(n12513), .Z(n12515) );
  XOR U22968 ( .A(n13157), .B(n13158), .Z(n12513) );
  ANDN U22969 ( .B(n13159), .A(n13160), .Z(n13157) );
  AND U22970 ( .A(a[3]), .B(b[105]), .Z(n13156) );
  XNOR U22971 ( .A(n13161), .B(n12518), .Z(n12520) );
  XOR U22972 ( .A(n13162), .B(n13163), .Z(n12518) );
  ANDN U22973 ( .B(n13164), .A(n13165), .Z(n13162) );
  AND U22974 ( .A(a[4]), .B(b[104]), .Z(n13161) );
  XNOR U22975 ( .A(n13166), .B(n12523), .Z(n12525) );
  XOR U22976 ( .A(n13167), .B(n13168), .Z(n12523) );
  ANDN U22977 ( .B(n13169), .A(n13170), .Z(n13167) );
  AND U22978 ( .A(a[5]), .B(b[103]), .Z(n13166) );
  XNOR U22979 ( .A(n13171), .B(n12528), .Z(n12530) );
  XOR U22980 ( .A(n13172), .B(n13173), .Z(n12528) );
  ANDN U22981 ( .B(n13174), .A(n13175), .Z(n13172) );
  AND U22982 ( .A(a[6]), .B(b[102]), .Z(n13171) );
  XNOR U22983 ( .A(n13176), .B(n12533), .Z(n12535) );
  XOR U22984 ( .A(n13177), .B(n13178), .Z(n12533) );
  ANDN U22985 ( .B(n13179), .A(n13180), .Z(n13177) );
  AND U22986 ( .A(a[7]), .B(b[101]), .Z(n13176) );
  XNOR U22987 ( .A(n13181), .B(n12538), .Z(n12540) );
  XOR U22988 ( .A(n13182), .B(n13183), .Z(n12538) );
  ANDN U22989 ( .B(n13184), .A(n13185), .Z(n13182) );
  AND U22990 ( .A(a[8]), .B(b[100]), .Z(n13181) );
  XNOR U22991 ( .A(n13186), .B(n12543), .Z(n12545) );
  XOR U22992 ( .A(n13187), .B(n13188), .Z(n12543) );
  ANDN U22993 ( .B(n13189), .A(n13190), .Z(n13187) );
  AND U22994 ( .A(a[9]), .B(b[99]), .Z(n13186) );
  XNOR U22995 ( .A(n13191), .B(n12548), .Z(n12550) );
  XOR U22996 ( .A(n13192), .B(n13193), .Z(n12548) );
  ANDN U22997 ( .B(n13194), .A(n13195), .Z(n13192) );
  AND U22998 ( .A(a[10]), .B(b[98]), .Z(n13191) );
  XNOR U22999 ( .A(n13196), .B(n12553), .Z(n12555) );
  XOR U23000 ( .A(n13197), .B(n13198), .Z(n12553) );
  ANDN U23001 ( .B(n13199), .A(n13200), .Z(n13197) );
  AND U23002 ( .A(a[11]), .B(b[97]), .Z(n13196) );
  XNOR U23003 ( .A(n13201), .B(n12558), .Z(n12560) );
  XOR U23004 ( .A(n13202), .B(n13203), .Z(n12558) );
  ANDN U23005 ( .B(n13204), .A(n13205), .Z(n13202) );
  AND U23006 ( .A(a[12]), .B(b[96]), .Z(n13201) );
  XNOR U23007 ( .A(n13206), .B(n12563), .Z(n12565) );
  XOR U23008 ( .A(n13207), .B(n13208), .Z(n12563) );
  ANDN U23009 ( .B(n13209), .A(n13210), .Z(n13207) );
  AND U23010 ( .A(a[13]), .B(b[95]), .Z(n13206) );
  XNOR U23011 ( .A(n13211), .B(n12568), .Z(n12570) );
  XOR U23012 ( .A(n13212), .B(n13213), .Z(n12568) );
  ANDN U23013 ( .B(n13214), .A(n13215), .Z(n13212) );
  AND U23014 ( .A(a[14]), .B(b[94]), .Z(n13211) );
  XNOR U23015 ( .A(n13216), .B(n12573), .Z(n12575) );
  XOR U23016 ( .A(n13217), .B(n13218), .Z(n12573) );
  ANDN U23017 ( .B(n13219), .A(n13220), .Z(n13217) );
  AND U23018 ( .A(a[15]), .B(b[93]), .Z(n13216) );
  XNOR U23019 ( .A(n13221), .B(n12578), .Z(n12580) );
  XOR U23020 ( .A(n13222), .B(n13223), .Z(n12578) );
  ANDN U23021 ( .B(n13224), .A(n13225), .Z(n13222) );
  AND U23022 ( .A(a[16]), .B(b[92]), .Z(n13221) );
  XNOR U23023 ( .A(n13226), .B(n12583), .Z(n12585) );
  XOR U23024 ( .A(n13227), .B(n13228), .Z(n12583) );
  ANDN U23025 ( .B(n13229), .A(n13230), .Z(n13227) );
  AND U23026 ( .A(a[17]), .B(b[91]), .Z(n13226) );
  XNOR U23027 ( .A(n13231), .B(n12588), .Z(n12590) );
  XOR U23028 ( .A(n13232), .B(n13233), .Z(n12588) );
  ANDN U23029 ( .B(n13234), .A(n13235), .Z(n13232) );
  AND U23030 ( .A(a[18]), .B(b[90]), .Z(n13231) );
  XNOR U23031 ( .A(n13236), .B(n12593), .Z(n12595) );
  XOR U23032 ( .A(n13237), .B(n13238), .Z(n12593) );
  ANDN U23033 ( .B(n13239), .A(n13240), .Z(n13237) );
  AND U23034 ( .A(a[19]), .B(b[89]), .Z(n13236) );
  XNOR U23035 ( .A(n13241), .B(n12598), .Z(n12600) );
  XOR U23036 ( .A(n13242), .B(n13243), .Z(n12598) );
  ANDN U23037 ( .B(n13244), .A(n13245), .Z(n13242) );
  AND U23038 ( .A(a[20]), .B(b[88]), .Z(n13241) );
  XNOR U23039 ( .A(n13246), .B(n12603), .Z(n12605) );
  XOR U23040 ( .A(n13247), .B(n13248), .Z(n12603) );
  ANDN U23041 ( .B(n13249), .A(n13250), .Z(n13247) );
  AND U23042 ( .A(a[21]), .B(b[87]), .Z(n13246) );
  XNOR U23043 ( .A(n13251), .B(n12608), .Z(n12610) );
  XOR U23044 ( .A(n13252), .B(n13253), .Z(n12608) );
  ANDN U23045 ( .B(n13254), .A(n13255), .Z(n13252) );
  AND U23046 ( .A(a[22]), .B(b[86]), .Z(n13251) );
  XNOR U23047 ( .A(n13256), .B(n12613), .Z(n12615) );
  XOR U23048 ( .A(n13257), .B(n13258), .Z(n12613) );
  ANDN U23049 ( .B(n13259), .A(n13260), .Z(n13257) );
  AND U23050 ( .A(a[23]), .B(b[85]), .Z(n13256) );
  XNOR U23051 ( .A(n13261), .B(n12618), .Z(n12620) );
  XOR U23052 ( .A(n13262), .B(n13263), .Z(n12618) );
  ANDN U23053 ( .B(n13264), .A(n13265), .Z(n13262) );
  AND U23054 ( .A(a[24]), .B(b[84]), .Z(n13261) );
  XNOR U23055 ( .A(n13266), .B(n12623), .Z(n12625) );
  XOR U23056 ( .A(n13267), .B(n13268), .Z(n12623) );
  ANDN U23057 ( .B(n13269), .A(n13270), .Z(n13267) );
  AND U23058 ( .A(a[25]), .B(b[83]), .Z(n13266) );
  XNOR U23059 ( .A(n13271), .B(n12628), .Z(n12630) );
  XOR U23060 ( .A(n13272), .B(n13273), .Z(n12628) );
  ANDN U23061 ( .B(n13274), .A(n13275), .Z(n13272) );
  AND U23062 ( .A(a[26]), .B(b[82]), .Z(n13271) );
  XNOR U23063 ( .A(n13276), .B(n12633), .Z(n12635) );
  XOR U23064 ( .A(n13277), .B(n13278), .Z(n12633) );
  ANDN U23065 ( .B(n13279), .A(n13280), .Z(n13277) );
  AND U23066 ( .A(a[27]), .B(b[81]), .Z(n13276) );
  XNOR U23067 ( .A(n13281), .B(n12638), .Z(n12640) );
  XOR U23068 ( .A(n13282), .B(n13283), .Z(n12638) );
  ANDN U23069 ( .B(n13284), .A(n13285), .Z(n13282) );
  AND U23070 ( .A(a[28]), .B(b[80]), .Z(n13281) );
  XNOR U23071 ( .A(n13286), .B(n12643), .Z(n12645) );
  XOR U23072 ( .A(n13287), .B(n13288), .Z(n12643) );
  ANDN U23073 ( .B(n13289), .A(n13290), .Z(n13287) );
  AND U23074 ( .A(a[29]), .B(b[79]), .Z(n13286) );
  XNOR U23075 ( .A(n13291), .B(n12648), .Z(n12650) );
  XOR U23076 ( .A(n13292), .B(n13293), .Z(n12648) );
  ANDN U23077 ( .B(n13294), .A(n13295), .Z(n13292) );
  AND U23078 ( .A(a[30]), .B(b[78]), .Z(n13291) );
  XNOR U23079 ( .A(n13296), .B(n12653), .Z(n12655) );
  XOR U23080 ( .A(n13297), .B(n13298), .Z(n12653) );
  ANDN U23081 ( .B(n13299), .A(n13300), .Z(n13297) );
  AND U23082 ( .A(a[31]), .B(b[77]), .Z(n13296) );
  XNOR U23083 ( .A(n13301), .B(n12658), .Z(n12660) );
  XOR U23084 ( .A(n13302), .B(n13303), .Z(n12658) );
  ANDN U23085 ( .B(n13304), .A(n13305), .Z(n13302) );
  AND U23086 ( .A(a[32]), .B(b[76]), .Z(n13301) );
  XNOR U23087 ( .A(n13306), .B(n12663), .Z(n12665) );
  XOR U23088 ( .A(n13307), .B(n13308), .Z(n12663) );
  ANDN U23089 ( .B(n13309), .A(n13310), .Z(n13307) );
  AND U23090 ( .A(a[33]), .B(b[75]), .Z(n13306) );
  XNOR U23091 ( .A(n13311), .B(n12668), .Z(n12670) );
  XOR U23092 ( .A(n13312), .B(n13313), .Z(n12668) );
  ANDN U23093 ( .B(n13314), .A(n13315), .Z(n13312) );
  AND U23094 ( .A(a[34]), .B(b[74]), .Z(n13311) );
  XNOR U23095 ( .A(n13316), .B(n12673), .Z(n12675) );
  XOR U23096 ( .A(n13317), .B(n13318), .Z(n12673) );
  ANDN U23097 ( .B(n13319), .A(n13320), .Z(n13317) );
  AND U23098 ( .A(a[35]), .B(b[73]), .Z(n13316) );
  XNOR U23099 ( .A(n13321), .B(n12678), .Z(n12680) );
  XOR U23100 ( .A(n13322), .B(n13323), .Z(n12678) );
  ANDN U23101 ( .B(n13324), .A(n13325), .Z(n13322) );
  AND U23102 ( .A(a[36]), .B(b[72]), .Z(n13321) );
  XNOR U23103 ( .A(n13326), .B(n12683), .Z(n12685) );
  XOR U23104 ( .A(n13327), .B(n13328), .Z(n12683) );
  ANDN U23105 ( .B(n13329), .A(n13330), .Z(n13327) );
  AND U23106 ( .A(a[37]), .B(b[71]), .Z(n13326) );
  XNOR U23107 ( .A(n13331), .B(n12688), .Z(n12690) );
  XOR U23108 ( .A(n13332), .B(n13333), .Z(n12688) );
  ANDN U23109 ( .B(n13334), .A(n13335), .Z(n13332) );
  AND U23110 ( .A(a[38]), .B(b[70]), .Z(n13331) );
  XNOR U23111 ( .A(n13336), .B(n12693), .Z(n12695) );
  XOR U23112 ( .A(n13337), .B(n13338), .Z(n12693) );
  ANDN U23113 ( .B(n13339), .A(n13340), .Z(n13337) );
  AND U23114 ( .A(a[39]), .B(b[69]), .Z(n13336) );
  XNOR U23115 ( .A(n13341), .B(n12698), .Z(n12700) );
  XOR U23116 ( .A(n13342), .B(n13343), .Z(n12698) );
  ANDN U23117 ( .B(n13344), .A(n13345), .Z(n13342) );
  AND U23118 ( .A(a[40]), .B(b[68]), .Z(n13341) );
  XNOR U23119 ( .A(n13346), .B(n12703), .Z(n12705) );
  XOR U23120 ( .A(n13347), .B(n13348), .Z(n12703) );
  ANDN U23121 ( .B(n13349), .A(n13350), .Z(n13347) );
  AND U23122 ( .A(a[41]), .B(b[67]), .Z(n13346) );
  XNOR U23123 ( .A(n13351), .B(n12708), .Z(n12710) );
  XOR U23124 ( .A(n13352), .B(n13353), .Z(n12708) );
  ANDN U23125 ( .B(n13354), .A(n13355), .Z(n13352) );
  AND U23126 ( .A(a[42]), .B(b[66]), .Z(n13351) );
  XNOR U23127 ( .A(n13356), .B(n12713), .Z(n12715) );
  XOR U23128 ( .A(n13357), .B(n13358), .Z(n12713) );
  ANDN U23129 ( .B(n13359), .A(n13360), .Z(n13357) );
  AND U23130 ( .A(a[43]), .B(b[65]), .Z(n13356) );
  XNOR U23131 ( .A(n13361), .B(n12718), .Z(n12720) );
  XOR U23132 ( .A(n13362), .B(n13363), .Z(n12718) );
  ANDN U23133 ( .B(n13364), .A(n13365), .Z(n13362) );
  AND U23134 ( .A(a[44]), .B(b[64]), .Z(n13361) );
  XNOR U23135 ( .A(n13366), .B(n12723), .Z(n12725) );
  XOR U23136 ( .A(n13367), .B(n13368), .Z(n12723) );
  ANDN U23137 ( .B(n13369), .A(n13370), .Z(n13367) );
  AND U23138 ( .A(a[45]), .B(b[63]), .Z(n13366) );
  XNOR U23139 ( .A(n13371), .B(n12728), .Z(n12730) );
  XOR U23140 ( .A(n13372), .B(n13373), .Z(n12728) );
  ANDN U23141 ( .B(n13374), .A(n13375), .Z(n13372) );
  AND U23142 ( .A(a[46]), .B(b[62]), .Z(n13371) );
  XNOR U23143 ( .A(n13376), .B(n12733), .Z(n12735) );
  XOR U23144 ( .A(n13377), .B(n13378), .Z(n12733) );
  ANDN U23145 ( .B(n13379), .A(n13380), .Z(n13377) );
  AND U23146 ( .A(a[47]), .B(b[61]), .Z(n13376) );
  XNOR U23147 ( .A(n13381), .B(n12738), .Z(n12740) );
  XOR U23148 ( .A(n13382), .B(n13383), .Z(n12738) );
  ANDN U23149 ( .B(n13384), .A(n13385), .Z(n13382) );
  AND U23150 ( .A(a[48]), .B(b[60]), .Z(n13381) );
  XNOR U23151 ( .A(n13386), .B(n12743), .Z(n12745) );
  XOR U23152 ( .A(n13387), .B(n13388), .Z(n12743) );
  ANDN U23153 ( .B(n13389), .A(n13390), .Z(n13387) );
  AND U23154 ( .A(a[49]), .B(b[59]), .Z(n13386) );
  XNOR U23155 ( .A(n13391), .B(n12748), .Z(n12750) );
  XOR U23156 ( .A(n13392), .B(n13393), .Z(n12748) );
  ANDN U23157 ( .B(n13394), .A(n13395), .Z(n13392) );
  AND U23158 ( .A(a[50]), .B(b[58]), .Z(n13391) );
  XNOR U23159 ( .A(n13396), .B(n12753), .Z(n12755) );
  XOR U23160 ( .A(n13397), .B(n13398), .Z(n12753) );
  ANDN U23161 ( .B(n13399), .A(n13400), .Z(n13397) );
  AND U23162 ( .A(a[51]), .B(b[57]), .Z(n13396) );
  XNOR U23163 ( .A(n13401), .B(n12758), .Z(n12760) );
  XOR U23164 ( .A(n13402), .B(n13403), .Z(n12758) );
  ANDN U23165 ( .B(n13404), .A(n13405), .Z(n13402) );
  AND U23166 ( .A(a[52]), .B(b[56]), .Z(n13401) );
  XNOR U23167 ( .A(n13406), .B(n12763), .Z(n12765) );
  XOR U23168 ( .A(n13407), .B(n13408), .Z(n12763) );
  ANDN U23169 ( .B(n13409), .A(n13410), .Z(n13407) );
  AND U23170 ( .A(a[53]), .B(b[55]), .Z(n13406) );
  XNOR U23171 ( .A(n13411), .B(n12768), .Z(n12770) );
  XOR U23172 ( .A(n13412), .B(n13413), .Z(n12768) );
  ANDN U23173 ( .B(n13414), .A(n13415), .Z(n13412) );
  AND U23174 ( .A(a[54]), .B(b[54]), .Z(n13411) );
  XNOR U23175 ( .A(n13416), .B(n12773), .Z(n12775) );
  XOR U23176 ( .A(n13417), .B(n13418), .Z(n12773) );
  ANDN U23177 ( .B(n13419), .A(n13420), .Z(n13417) );
  AND U23178 ( .A(a[55]), .B(b[53]), .Z(n13416) );
  XNOR U23179 ( .A(n13421), .B(n12778), .Z(n12780) );
  XOR U23180 ( .A(n13422), .B(n13423), .Z(n12778) );
  ANDN U23181 ( .B(n13424), .A(n13425), .Z(n13422) );
  AND U23182 ( .A(a[56]), .B(b[52]), .Z(n13421) );
  XNOR U23183 ( .A(n13426), .B(n12783), .Z(n12785) );
  XOR U23184 ( .A(n13427), .B(n13428), .Z(n12783) );
  ANDN U23185 ( .B(n13429), .A(n13430), .Z(n13427) );
  AND U23186 ( .A(a[57]), .B(b[51]), .Z(n13426) );
  XNOR U23187 ( .A(n13431), .B(n12788), .Z(n12790) );
  XOR U23188 ( .A(n13432), .B(n13433), .Z(n12788) );
  ANDN U23189 ( .B(n13434), .A(n13435), .Z(n13432) );
  AND U23190 ( .A(a[58]), .B(b[50]), .Z(n13431) );
  XNOR U23191 ( .A(n13436), .B(n12793), .Z(n12795) );
  XOR U23192 ( .A(n13437), .B(n13438), .Z(n12793) );
  ANDN U23193 ( .B(n13439), .A(n13440), .Z(n13437) );
  AND U23194 ( .A(a[59]), .B(b[49]), .Z(n13436) );
  XNOR U23195 ( .A(n13441), .B(n12798), .Z(n12800) );
  XOR U23196 ( .A(n13442), .B(n13443), .Z(n12798) );
  ANDN U23197 ( .B(n13444), .A(n13445), .Z(n13442) );
  AND U23198 ( .A(a[60]), .B(b[48]), .Z(n13441) );
  XNOR U23199 ( .A(n13446), .B(n12803), .Z(n12805) );
  XOR U23200 ( .A(n13447), .B(n13448), .Z(n12803) );
  ANDN U23201 ( .B(n13449), .A(n13450), .Z(n13447) );
  AND U23202 ( .A(a[61]), .B(b[47]), .Z(n13446) );
  XNOR U23203 ( .A(n13451), .B(n12808), .Z(n12810) );
  XOR U23204 ( .A(n13452), .B(n13453), .Z(n12808) );
  ANDN U23205 ( .B(n13454), .A(n13455), .Z(n13452) );
  AND U23206 ( .A(a[62]), .B(b[46]), .Z(n13451) );
  XNOR U23207 ( .A(n13456), .B(n12813), .Z(n12815) );
  XOR U23208 ( .A(n13457), .B(n13458), .Z(n12813) );
  ANDN U23209 ( .B(n13459), .A(n13460), .Z(n13457) );
  AND U23210 ( .A(a[63]), .B(b[45]), .Z(n13456) );
  XNOR U23211 ( .A(n13461), .B(n12818), .Z(n12820) );
  XOR U23212 ( .A(n13462), .B(n13463), .Z(n12818) );
  ANDN U23213 ( .B(n13464), .A(n13465), .Z(n13462) );
  AND U23214 ( .A(a[64]), .B(b[44]), .Z(n13461) );
  XNOR U23215 ( .A(n13466), .B(n12823), .Z(n12825) );
  XOR U23216 ( .A(n13467), .B(n13468), .Z(n12823) );
  ANDN U23217 ( .B(n13469), .A(n13470), .Z(n13467) );
  AND U23218 ( .A(a[65]), .B(b[43]), .Z(n13466) );
  XNOR U23219 ( .A(n13471), .B(n12828), .Z(n12830) );
  XOR U23220 ( .A(n13472), .B(n13473), .Z(n12828) );
  ANDN U23221 ( .B(n13474), .A(n13475), .Z(n13472) );
  AND U23222 ( .A(a[66]), .B(b[42]), .Z(n13471) );
  XNOR U23223 ( .A(n13476), .B(n12833), .Z(n12835) );
  XOR U23224 ( .A(n13477), .B(n13478), .Z(n12833) );
  ANDN U23225 ( .B(n13479), .A(n13480), .Z(n13477) );
  AND U23226 ( .A(a[67]), .B(b[41]), .Z(n13476) );
  XNOR U23227 ( .A(n13481), .B(n12838), .Z(n12840) );
  XOR U23228 ( .A(n13482), .B(n13483), .Z(n12838) );
  ANDN U23229 ( .B(n13484), .A(n13485), .Z(n13482) );
  AND U23230 ( .A(a[68]), .B(b[40]), .Z(n13481) );
  XNOR U23231 ( .A(n13486), .B(n12843), .Z(n12845) );
  XOR U23232 ( .A(n13487), .B(n13488), .Z(n12843) );
  ANDN U23233 ( .B(n13489), .A(n13490), .Z(n13487) );
  AND U23234 ( .A(a[69]), .B(b[39]), .Z(n13486) );
  XNOR U23235 ( .A(n13491), .B(n12848), .Z(n12850) );
  XOR U23236 ( .A(n13492), .B(n13493), .Z(n12848) );
  ANDN U23237 ( .B(n13494), .A(n13495), .Z(n13492) );
  AND U23238 ( .A(a[70]), .B(b[38]), .Z(n13491) );
  XNOR U23239 ( .A(n13496), .B(n12853), .Z(n12855) );
  XOR U23240 ( .A(n13497), .B(n13498), .Z(n12853) );
  ANDN U23241 ( .B(n13499), .A(n13500), .Z(n13497) );
  AND U23242 ( .A(a[71]), .B(b[37]), .Z(n13496) );
  XNOR U23243 ( .A(n13501), .B(n12858), .Z(n12860) );
  XOR U23244 ( .A(n13502), .B(n13503), .Z(n12858) );
  ANDN U23245 ( .B(n13504), .A(n13505), .Z(n13502) );
  AND U23246 ( .A(a[72]), .B(b[36]), .Z(n13501) );
  XNOR U23247 ( .A(n13506), .B(n12863), .Z(n12865) );
  XOR U23248 ( .A(n13507), .B(n13508), .Z(n12863) );
  ANDN U23249 ( .B(n13509), .A(n13510), .Z(n13507) );
  AND U23250 ( .A(a[73]), .B(b[35]), .Z(n13506) );
  XNOR U23251 ( .A(n13511), .B(n12868), .Z(n12870) );
  XOR U23252 ( .A(n13512), .B(n13513), .Z(n12868) );
  ANDN U23253 ( .B(n13514), .A(n13515), .Z(n13512) );
  AND U23254 ( .A(a[74]), .B(b[34]), .Z(n13511) );
  XNOR U23255 ( .A(n13516), .B(n12873), .Z(n12875) );
  XOR U23256 ( .A(n13517), .B(n13518), .Z(n12873) );
  ANDN U23257 ( .B(n13519), .A(n13520), .Z(n13517) );
  AND U23258 ( .A(a[75]), .B(b[33]), .Z(n13516) );
  XNOR U23259 ( .A(n13521), .B(n12878), .Z(n12880) );
  XOR U23260 ( .A(n13522), .B(n13523), .Z(n12878) );
  ANDN U23261 ( .B(n13524), .A(n13525), .Z(n13522) );
  AND U23262 ( .A(a[76]), .B(b[32]), .Z(n13521) );
  XNOR U23263 ( .A(n13526), .B(n12883), .Z(n12885) );
  XOR U23264 ( .A(n13527), .B(n13528), .Z(n12883) );
  ANDN U23265 ( .B(n13529), .A(n13530), .Z(n13527) );
  AND U23266 ( .A(a[77]), .B(b[31]), .Z(n13526) );
  XNOR U23267 ( .A(n13531), .B(n12888), .Z(n12890) );
  XOR U23268 ( .A(n13532), .B(n13533), .Z(n12888) );
  ANDN U23269 ( .B(n13534), .A(n13535), .Z(n13532) );
  AND U23270 ( .A(a[78]), .B(b[30]), .Z(n13531) );
  XNOR U23271 ( .A(n13536), .B(n12893), .Z(n12895) );
  XOR U23272 ( .A(n13537), .B(n13538), .Z(n12893) );
  ANDN U23273 ( .B(n13539), .A(n13540), .Z(n13537) );
  AND U23274 ( .A(a[79]), .B(b[29]), .Z(n13536) );
  XNOR U23275 ( .A(n13541), .B(n12898), .Z(n12900) );
  XOR U23276 ( .A(n13542), .B(n13543), .Z(n12898) );
  ANDN U23277 ( .B(n13544), .A(n13545), .Z(n13542) );
  AND U23278 ( .A(a[80]), .B(b[28]), .Z(n13541) );
  XNOR U23279 ( .A(n13546), .B(n12903), .Z(n12905) );
  XOR U23280 ( .A(n13547), .B(n13548), .Z(n12903) );
  ANDN U23281 ( .B(n13549), .A(n13550), .Z(n13547) );
  AND U23282 ( .A(a[81]), .B(b[27]), .Z(n13546) );
  XNOR U23283 ( .A(n13551), .B(n12908), .Z(n12910) );
  XOR U23284 ( .A(n13552), .B(n13553), .Z(n12908) );
  ANDN U23285 ( .B(n13554), .A(n13555), .Z(n13552) );
  AND U23286 ( .A(a[82]), .B(b[26]), .Z(n13551) );
  XNOR U23287 ( .A(n13556), .B(n12913), .Z(n12915) );
  XOR U23288 ( .A(n13557), .B(n13558), .Z(n12913) );
  ANDN U23289 ( .B(n13559), .A(n13560), .Z(n13557) );
  AND U23290 ( .A(a[83]), .B(b[25]), .Z(n13556) );
  XNOR U23291 ( .A(n13561), .B(n12918), .Z(n12920) );
  XOR U23292 ( .A(n13562), .B(n13563), .Z(n12918) );
  ANDN U23293 ( .B(n13564), .A(n13565), .Z(n13562) );
  AND U23294 ( .A(a[84]), .B(b[24]), .Z(n13561) );
  XNOR U23295 ( .A(n13566), .B(n12923), .Z(n12925) );
  XOR U23296 ( .A(n13567), .B(n13568), .Z(n12923) );
  ANDN U23297 ( .B(n13569), .A(n13570), .Z(n13567) );
  AND U23298 ( .A(a[85]), .B(b[23]), .Z(n13566) );
  XNOR U23299 ( .A(n13571), .B(n12928), .Z(n12930) );
  XOR U23300 ( .A(n13572), .B(n13573), .Z(n12928) );
  ANDN U23301 ( .B(n13574), .A(n13575), .Z(n13572) );
  AND U23302 ( .A(a[86]), .B(b[22]), .Z(n13571) );
  XNOR U23303 ( .A(n13576), .B(n12933), .Z(n12935) );
  XOR U23304 ( .A(n13577), .B(n13578), .Z(n12933) );
  ANDN U23305 ( .B(n13579), .A(n13580), .Z(n13577) );
  AND U23306 ( .A(a[87]), .B(b[21]), .Z(n13576) );
  XNOR U23307 ( .A(n13581), .B(n12938), .Z(n12940) );
  XOR U23308 ( .A(n13582), .B(n13583), .Z(n12938) );
  ANDN U23309 ( .B(n13584), .A(n13585), .Z(n13582) );
  AND U23310 ( .A(a[88]), .B(b[20]), .Z(n13581) );
  XNOR U23311 ( .A(n13586), .B(n12943), .Z(n12945) );
  XOR U23312 ( .A(n13587), .B(n13588), .Z(n12943) );
  ANDN U23313 ( .B(n13589), .A(n13590), .Z(n13587) );
  AND U23314 ( .A(a[89]), .B(b[19]), .Z(n13586) );
  XNOR U23315 ( .A(n13591), .B(n12948), .Z(n12950) );
  XOR U23316 ( .A(n13592), .B(n13593), .Z(n12948) );
  ANDN U23317 ( .B(n13594), .A(n13595), .Z(n13592) );
  AND U23318 ( .A(a[90]), .B(b[18]), .Z(n13591) );
  XNOR U23319 ( .A(n13596), .B(n12953), .Z(n12955) );
  XOR U23320 ( .A(n13597), .B(n13598), .Z(n12953) );
  ANDN U23321 ( .B(n13599), .A(n13600), .Z(n13597) );
  AND U23322 ( .A(a[91]), .B(b[17]), .Z(n13596) );
  XNOR U23323 ( .A(n13601), .B(n12958), .Z(n12960) );
  XOR U23324 ( .A(n13602), .B(n13603), .Z(n12958) );
  ANDN U23325 ( .B(n13604), .A(n13605), .Z(n13602) );
  AND U23326 ( .A(a[92]), .B(b[16]), .Z(n13601) );
  XNOR U23327 ( .A(n13606), .B(n12963), .Z(n12965) );
  XOR U23328 ( .A(n13607), .B(n13608), .Z(n12963) );
  ANDN U23329 ( .B(n13609), .A(n13610), .Z(n13607) );
  AND U23330 ( .A(a[93]), .B(b[15]), .Z(n13606) );
  XNOR U23331 ( .A(n13611), .B(n12968), .Z(n12970) );
  XOR U23332 ( .A(n13612), .B(n13613), .Z(n12968) );
  ANDN U23333 ( .B(n13614), .A(n13615), .Z(n13612) );
  AND U23334 ( .A(a[94]), .B(b[14]), .Z(n13611) );
  XNOR U23335 ( .A(n13616), .B(n12973), .Z(n12975) );
  XOR U23336 ( .A(n13617), .B(n13618), .Z(n12973) );
  ANDN U23337 ( .B(n13619), .A(n13620), .Z(n13617) );
  AND U23338 ( .A(a[95]), .B(b[13]), .Z(n13616) );
  XNOR U23339 ( .A(n13621), .B(n12978), .Z(n12980) );
  XOR U23340 ( .A(n13622), .B(n13623), .Z(n12978) );
  ANDN U23341 ( .B(n13624), .A(n13625), .Z(n13622) );
  AND U23342 ( .A(a[96]), .B(b[12]), .Z(n13621) );
  XNOR U23343 ( .A(n13626), .B(n12983), .Z(n12985) );
  XOR U23344 ( .A(n13627), .B(n13628), .Z(n12983) );
  ANDN U23345 ( .B(n13629), .A(n13630), .Z(n13627) );
  AND U23346 ( .A(a[97]), .B(b[11]), .Z(n13626) );
  XNOR U23347 ( .A(n13631), .B(n12988), .Z(n12990) );
  XOR U23348 ( .A(n13632), .B(n13633), .Z(n12988) );
  ANDN U23349 ( .B(n13634), .A(n13635), .Z(n13632) );
  AND U23350 ( .A(a[98]), .B(b[10]), .Z(n13631) );
  XNOR U23351 ( .A(n13636), .B(n12993), .Z(n12995) );
  XOR U23352 ( .A(n13637), .B(n13638), .Z(n12993) );
  ANDN U23353 ( .B(n13639), .A(n13640), .Z(n13637) );
  AND U23354 ( .A(b[9]), .B(a[99]), .Z(n13636) );
  XNOR U23355 ( .A(n13641), .B(n12998), .Z(n13000) );
  XOR U23356 ( .A(n13642), .B(n13643), .Z(n12998) );
  ANDN U23357 ( .B(n13644), .A(n13645), .Z(n13642) );
  AND U23358 ( .A(b[8]), .B(a[100]), .Z(n13641) );
  XNOR U23359 ( .A(n13646), .B(n13003), .Z(n13005) );
  XOR U23360 ( .A(n13647), .B(n13648), .Z(n13003) );
  ANDN U23361 ( .B(n13649), .A(n13650), .Z(n13647) );
  AND U23362 ( .A(b[7]), .B(a[101]), .Z(n13646) );
  XNOR U23363 ( .A(n13651), .B(n13008), .Z(n13010) );
  XOR U23364 ( .A(n13652), .B(n13653), .Z(n13008) );
  ANDN U23365 ( .B(n13654), .A(n13655), .Z(n13652) );
  AND U23366 ( .A(b[6]), .B(a[102]), .Z(n13651) );
  XNOR U23367 ( .A(n13656), .B(n13013), .Z(n13015) );
  XOR U23368 ( .A(n13657), .B(n13658), .Z(n13013) );
  ANDN U23369 ( .B(n13659), .A(n13660), .Z(n13657) );
  AND U23370 ( .A(b[5]), .B(a[103]), .Z(n13656) );
  XNOR U23371 ( .A(n13661), .B(n13018), .Z(n13020) );
  XOR U23372 ( .A(n13662), .B(n13663), .Z(n13018) );
  ANDN U23373 ( .B(n13664), .A(n13665), .Z(n13662) );
  AND U23374 ( .A(b[4]), .B(a[104]), .Z(n13661) );
  XNOR U23375 ( .A(n13666), .B(n13667), .Z(n13032) );
  NANDN U23376 ( .A(n13668), .B(n13669), .Z(n13667) );
  XNOR U23377 ( .A(n13670), .B(n13023), .Z(n13025) );
  XNOR U23378 ( .A(n13671), .B(n13672), .Z(n13023) );
  AND U23379 ( .A(n13673), .B(n13674), .Z(n13671) );
  AND U23380 ( .A(b[3]), .B(a[105]), .Z(n13670) );
  NAND U23381 ( .A(a[108]), .B(b[0]), .Z(n12392) );
  XNOR U23382 ( .A(n13038), .B(n13039), .Z(c[107]) );
  XNOR U23383 ( .A(n13668), .B(n13669), .Z(n13039) );
  XOR U23384 ( .A(n13666), .B(n13675), .Z(n13669) );
  NAND U23385 ( .A(b[1]), .B(a[106]), .Z(n13675) );
  XOR U23386 ( .A(n13674), .B(n13676), .Z(n13668) );
  XOR U23387 ( .A(n13666), .B(n13673), .Z(n13676) );
  XNOR U23388 ( .A(n13677), .B(n13672), .Z(n13673) );
  AND U23389 ( .A(b[2]), .B(a[105]), .Z(n13677) );
  NANDN U23390 ( .A(n13678), .B(n13679), .Z(n13666) );
  XOR U23391 ( .A(n13672), .B(n13664), .Z(n13680) );
  XNOR U23392 ( .A(n13663), .B(n13659), .Z(n13681) );
  XNOR U23393 ( .A(n13658), .B(n13654), .Z(n13682) );
  XNOR U23394 ( .A(n13653), .B(n13649), .Z(n13683) );
  XNOR U23395 ( .A(n13648), .B(n13644), .Z(n13684) );
  XNOR U23396 ( .A(n13643), .B(n13639), .Z(n13685) );
  XNOR U23397 ( .A(n13638), .B(n13634), .Z(n13686) );
  XNOR U23398 ( .A(n13633), .B(n13629), .Z(n13687) );
  XNOR U23399 ( .A(n13628), .B(n13624), .Z(n13688) );
  XNOR U23400 ( .A(n13623), .B(n13619), .Z(n13689) );
  XNOR U23401 ( .A(n13618), .B(n13614), .Z(n13690) );
  XNOR U23402 ( .A(n13613), .B(n13609), .Z(n13691) );
  XNOR U23403 ( .A(n13608), .B(n13604), .Z(n13692) );
  XNOR U23404 ( .A(n13603), .B(n13599), .Z(n13693) );
  XNOR U23405 ( .A(n13598), .B(n13594), .Z(n13694) );
  XNOR U23406 ( .A(n13593), .B(n13589), .Z(n13695) );
  XNOR U23407 ( .A(n13588), .B(n13584), .Z(n13696) );
  XNOR U23408 ( .A(n13583), .B(n13579), .Z(n13697) );
  XNOR U23409 ( .A(n13578), .B(n13574), .Z(n13698) );
  XNOR U23410 ( .A(n13573), .B(n13569), .Z(n13699) );
  XNOR U23411 ( .A(n13568), .B(n13564), .Z(n13700) );
  XNOR U23412 ( .A(n13563), .B(n13559), .Z(n13701) );
  XNOR U23413 ( .A(n13558), .B(n13554), .Z(n13702) );
  XNOR U23414 ( .A(n13553), .B(n13549), .Z(n13703) );
  XNOR U23415 ( .A(n13548), .B(n13544), .Z(n13704) );
  XNOR U23416 ( .A(n13543), .B(n13539), .Z(n13705) );
  XNOR U23417 ( .A(n13538), .B(n13534), .Z(n13706) );
  XNOR U23418 ( .A(n13533), .B(n13529), .Z(n13707) );
  XNOR U23419 ( .A(n13528), .B(n13524), .Z(n13708) );
  XNOR U23420 ( .A(n13523), .B(n13519), .Z(n13709) );
  XNOR U23421 ( .A(n13518), .B(n13514), .Z(n13710) );
  XNOR U23422 ( .A(n13513), .B(n13509), .Z(n13711) );
  XNOR U23423 ( .A(n13508), .B(n13504), .Z(n13712) );
  XNOR U23424 ( .A(n13503), .B(n13499), .Z(n13713) );
  XNOR U23425 ( .A(n13498), .B(n13494), .Z(n13714) );
  XNOR U23426 ( .A(n13493), .B(n13489), .Z(n13715) );
  XNOR U23427 ( .A(n13488), .B(n13484), .Z(n13716) );
  XNOR U23428 ( .A(n13483), .B(n13479), .Z(n13717) );
  XNOR U23429 ( .A(n13478), .B(n13474), .Z(n13718) );
  XNOR U23430 ( .A(n13473), .B(n13469), .Z(n13719) );
  XNOR U23431 ( .A(n13468), .B(n13464), .Z(n13720) );
  XNOR U23432 ( .A(n13463), .B(n13459), .Z(n13721) );
  XNOR U23433 ( .A(n13458), .B(n13454), .Z(n13722) );
  XNOR U23434 ( .A(n13453), .B(n13449), .Z(n13723) );
  XNOR U23435 ( .A(n13448), .B(n13444), .Z(n13724) );
  XNOR U23436 ( .A(n13443), .B(n13439), .Z(n13725) );
  XNOR U23437 ( .A(n13438), .B(n13434), .Z(n13726) );
  XNOR U23438 ( .A(n13433), .B(n13429), .Z(n13727) );
  XNOR U23439 ( .A(n13428), .B(n13424), .Z(n13728) );
  XNOR U23440 ( .A(n13423), .B(n13419), .Z(n13729) );
  XNOR U23441 ( .A(n13418), .B(n13414), .Z(n13730) );
  XNOR U23442 ( .A(n13413), .B(n13409), .Z(n13731) );
  XNOR U23443 ( .A(n13408), .B(n13404), .Z(n13732) );
  XNOR U23444 ( .A(n13403), .B(n13399), .Z(n13733) );
  XNOR U23445 ( .A(n13398), .B(n13394), .Z(n13734) );
  XNOR U23446 ( .A(n13393), .B(n13389), .Z(n13735) );
  XNOR U23447 ( .A(n13388), .B(n13384), .Z(n13736) );
  XNOR U23448 ( .A(n13383), .B(n13379), .Z(n13737) );
  XNOR U23449 ( .A(n13378), .B(n13374), .Z(n13738) );
  XNOR U23450 ( .A(n13373), .B(n13369), .Z(n13739) );
  XNOR U23451 ( .A(n13368), .B(n13364), .Z(n13740) );
  XNOR U23452 ( .A(n13363), .B(n13359), .Z(n13741) );
  XNOR U23453 ( .A(n13358), .B(n13354), .Z(n13742) );
  XNOR U23454 ( .A(n13353), .B(n13349), .Z(n13743) );
  XNOR U23455 ( .A(n13348), .B(n13344), .Z(n13744) );
  XNOR U23456 ( .A(n13343), .B(n13339), .Z(n13745) );
  XNOR U23457 ( .A(n13338), .B(n13334), .Z(n13746) );
  XNOR U23458 ( .A(n13333), .B(n13329), .Z(n13747) );
  XNOR U23459 ( .A(n13328), .B(n13324), .Z(n13748) );
  XNOR U23460 ( .A(n13323), .B(n13319), .Z(n13749) );
  XNOR U23461 ( .A(n13318), .B(n13314), .Z(n13750) );
  XNOR U23462 ( .A(n13313), .B(n13309), .Z(n13751) );
  XNOR U23463 ( .A(n13308), .B(n13304), .Z(n13752) );
  XNOR U23464 ( .A(n13303), .B(n13299), .Z(n13753) );
  XNOR U23465 ( .A(n13298), .B(n13294), .Z(n13754) );
  XNOR U23466 ( .A(n13293), .B(n13289), .Z(n13755) );
  XNOR U23467 ( .A(n13288), .B(n13284), .Z(n13756) );
  XNOR U23468 ( .A(n13283), .B(n13279), .Z(n13757) );
  XNOR U23469 ( .A(n13278), .B(n13274), .Z(n13758) );
  XNOR U23470 ( .A(n13273), .B(n13269), .Z(n13759) );
  XNOR U23471 ( .A(n13268), .B(n13264), .Z(n13760) );
  XNOR U23472 ( .A(n13263), .B(n13259), .Z(n13761) );
  XNOR U23473 ( .A(n13258), .B(n13254), .Z(n13762) );
  XNOR U23474 ( .A(n13253), .B(n13249), .Z(n13763) );
  XNOR U23475 ( .A(n13248), .B(n13244), .Z(n13764) );
  XNOR U23476 ( .A(n13243), .B(n13239), .Z(n13765) );
  XNOR U23477 ( .A(n13238), .B(n13234), .Z(n13766) );
  XNOR U23478 ( .A(n13233), .B(n13229), .Z(n13767) );
  XNOR U23479 ( .A(n13228), .B(n13224), .Z(n13768) );
  XNOR U23480 ( .A(n13223), .B(n13219), .Z(n13769) );
  XNOR U23481 ( .A(n13218), .B(n13214), .Z(n13770) );
  XNOR U23482 ( .A(n13213), .B(n13209), .Z(n13771) );
  XNOR U23483 ( .A(n13208), .B(n13204), .Z(n13772) );
  XNOR U23484 ( .A(n13203), .B(n13199), .Z(n13773) );
  XNOR U23485 ( .A(n13198), .B(n13194), .Z(n13774) );
  XNOR U23486 ( .A(n13193), .B(n13189), .Z(n13775) );
  XNOR U23487 ( .A(n13188), .B(n13184), .Z(n13776) );
  XNOR U23488 ( .A(n13183), .B(n13179), .Z(n13777) );
  XNOR U23489 ( .A(n13178), .B(n13174), .Z(n13778) );
  XNOR U23490 ( .A(n13173), .B(n13169), .Z(n13779) );
  XNOR U23491 ( .A(n13168), .B(n13164), .Z(n13780) );
  XNOR U23492 ( .A(n13163), .B(n13159), .Z(n13781) );
  XNOR U23493 ( .A(n13158), .B(n13154), .Z(n13782) );
  XNOR U23494 ( .A(n13153), .B(n13149), .Z(n13783) );
  XNOR U23495 ( .A(n13784), .B(n13148), .Z(n13149) );
  AND U23496 ( .A(a[0]), .B(b[107]), .Z(n13784) );
  XOR U23497 ( .A(n13785), .B(n13148), .Z(n13150) );
  XNOR U23498 ( .A(n13786), .B(n13787), .Z(n13148) );
  ANDN U23499 ( .B(n13788), .A(n13789), .Z(n13786) );
  AND U23500 ( .A(a[1]), .B(b[106]), .Z(n13785) );
  XNOR U23501 ( .A(n13790), .B(n13153), .Z(n13155) );
  XOR U23502 ( .A(n13791), .B(n13792), .Z(n13153) );
  ANDN U23503 ( .B(n13793), .A(n13794), .Z(n13791) );
  AND U23504 ( .A(a[2]), .B(b[105]), .Z(n13790) );
  XNOR U23505 ( .A(n13795), .B(n13158), .Z(n13160) );
  XOR U23506 ( .A(n13796), .B(n13797), .Z(n13158) );
  ANDN U23507 ( .B(n13798), .A(n13799), .Z(n13796) );
  AND U23508 ( .A(a[3]), .B(b[104]), .Z(n13795) );
  XNOR U23509 ( .A(n13800), .B(n13163), .Z(n13165) );
  XOR U23510 ( .A(n13801), .B(n13802), .Z(n13163) );
  ANDN U23511 ( .B(n13803), .A(n13804), .Z(n13801) );
  AND U23512 ( .A(a[4]), .B(b[103]), .Z(n13800) );
  XNOR U23513 ( .A(n13805), .B(n13168), .Z(n13170) );
  XOR U23514 ( .A(n13806), .B(n13807), .Z(n13168) );
  ANDN U23515 ( .B(n13808), .A(n13809), .Z(n13806) );
  AND U23516 ( .A(a[5]), .B(b[102]), .Z(n13805) );
  XNOR U23517 ( .A(n13810), .B(n13173), .Z(n13175) );
  XOR U23518 ( .A(n13811), .B(n13812), .Z(n13173) );
  ANDN U23519 ( .B(n13813), .A(n13814), .Z(n13811) );
  AND U23520 ( .A(a[6]), .B(b[101]), .Z(n13810) );
  XNOR U23521 ( .A(n13815), .B(n13178), .Z(n13180) );
  XOR U23522 ( .A(n13816), .B(n13817), .Z(n13178) );
  ANDN U23523 ( .B(n13818), .A(n13819), .Z(n13816) );
  AND U23524 ( .A(a[7]), .B(b[100]), .Z(n13815) );
  XNOR U23525 ( .A(n13820), .B(n13183), .Z(n13185) );
  XOR U23526 ( .A(n13821), .B(n13822), .Z(n13183) );
  ANDN U23527 ( .B(n13823), .A(n13824), .Z(n13821) );
  AND U23528 ( .A(a[8]), .B(b[99]), .Z(n13820) );
  XNOR U23529 ( .A(n13825), .B(n13188), .Z(n13190) );
  XOR U23530 ( .A(n13826), .B(n13827), .Z(n13188) );
  ANDN U23531 ( .B(n13828), .A(n13829), .Z(n13826) );
  AND U23532 ( .A(a[9]), .B(b[98]), .Z(n13825) );
  XNOR U23533 ( .A(n13830), .B(n13193), .Z(n13195) );
  XOR U23534 ( .A(n13831), .B(n13832), .Z(n13193) );
  ANDN U23535 ( .B(n13833), .A(n13834), .Z(n13831) );
  AND U23536 ( .A(a[10]), .B(b[97]), .Z(n13830) );
  XNOR U23537 ( .A(n13835), .B(n13198), .Z(n13200) );
  XOR U23538 ( .A(n13836), .B(n13837), .Z(n13198) );
  ANDN U23539 ( .B(n13838), .A(n13839), .Z(n13836) );
  AND U23540 ( .A(a[11]), .B(b[96]), .Z(n13835) );
  XNOR U23541 ( .A(n13840), .B(n13203), .Z(n13205) );
  XOR U23542 ( .A(n13841), .B(n13842), .Z(n13203) );
  ANDN U23543 ( .B(n13843), .A(n13844), .Z(n13841) );
  AND U23544 ( .A(a[12]), .B(b[95]), .Z(n13840) );
  XNOR U23545 ( .A(n13845), .B(n13208), .Z(n13210) );
  XOR U23546 ( .A(n13846), .B(n13847), .Z(n13208) );
  ANDN U23547 ( .B(n13848), .A(n13849), .Z(n13846) );
  AND U23548 ( .A(a[13]), .B(b[94]), .Z(n13845) );
  XNOR U23549 ( .A(n13850), .B(n13213), .Z(n13215) );
  XOR U23550 ( .A(n13851), .B(n13852), .Z(n13213) );
  ANDN U23551 ( .B(n13853), .A(n13854), .Z(n13851) );
  AND U23552 ( .A(a[14]), .B(b[93]), .Z(n13850) );
  XNOR U23553 ( .A(n13855), .B(n13218), .Z(n13220) );
  XOR U23554 ( .A(n13856), .B(n13857), .Z(n13218) );
  ANDN U23555 ( .B(n13858), .A(n13859), .Z(n13856) );
  AND U23556 ( .A(a[15]), .B(b[92]), .Z(n13855) );
  XNOR U23557 ( .A(n13860), .B(n13223), .Z(n13225) );
  XOR U23558 ( .A(n13861), .B(n13862), .Z(n13223) );
  ANDN U23559 ( .B(n13863), .A(n13864), .Z(n13861) );
  AND U23560 ( .A(a[16]), .B(b[91]), .Z(n13860) );
  XNOR U23561 ( .A(n13865), .B(n13228), .Z(n13230) );
  XOR U23562 ( .A(n13866), .B(n13867), .Z(n13228) );
  ANDN U23563 ( .B(n13868), .A(n13869), .Z(n13866) );
  AND U23564 ( .A(a[17]), .B(b[90]), .Z(n13865) );
  XNOR U23565 ( .A(n13870), .B(n13233), .Z(n13235) );
  XOR U23566 ( .A(n13871), .B(n13872), .Z(n13233) );
  ANDN U23567 ( .B(n13873), .A(n13874), .Z(n13871) );
  AND U23568 ( .A(a[18]), .B(b[89]), .Z(n13870) );
  XNOR U23569 ( .A(n13875), .B(n13238), .Z(n13240) );
  XOR U23570 ( .A(n13876), .B(n13877), .Z(n13238) );
  ANDN U23571 ( .B(n13878), .A(n13879), .Z(n13876) );
  AND U23572 ( .A(a[19]), .B(b[88]), .Z(n13875) );
  XNOR U23573 ( .A(n13880), .B(n13243), .Z(n13245) );
  XOR U23574 ( .A(n13881), .B(n13882), .Z(n13243) );
  ANDN U23575 ( .B(n13883), .A(n13884), .Z(n13881) );
  AND U23576 ( .A(a[20]), .B(b[87]), .Z(n13880) );
  XNOR U23577 ( .A(n13885), .B(n13248), .Z(n13250) );
  XOR U23578 ( .A(n13886), .B(n13887), .Z(n13248) );
  ANDN U23579 ( .B(n13888), .A(n13889), .Z(n13886) );
  AND U23580 ( .A(a[21]), .B(b[86]), .Z(n13885) );
  XNOR U23581 ( .A(n13890), .B(n13253), .Z(n13255) );
  XOR U23582 ( .A(n13891), .B(n13892), .Z(n13253) );
  ANDN U23583 ( .B(n13893), .A(n13894), .Z(n13891) );
  AND U23584 ( .A(a[22]), .B(b[85]), .Z(n13890) );
  XNOR U23585 ( .A(n13895), .B(n13258), .Z(n13260) );
  XOR U23586 ( .A(n13896), .B(n13897), .Z(n13258) );
  ANDN U23587 ( .B(n13898), .A(n13899), .Z(n13896) );
  AND U23588 ( .A(a[23]), .B(b[84]), .Z(n13895) );
  XNOR U23589 ( .A(n13900), .B(n13263), .Z(n13265) );
  XOR U23590 ( .A(n13901), .B(n13902), .Z(n13263) );
  ANDN U23591 ( .B(n13903), .A(n13904), .Z(n13901) );
  AND U23592 ( .A(a[24]), .B(b[83]), .Z(n13900) );
  XNOR U23593 ( .A(n13905), .B(n13268), .Z(n13270) );
  XOR U23594 ( .A(n13906), .B(n13907), .Z(n13268) );
  ANDN U23595 ( .B(n13908), .A(n13909), .Z(n13906) );
  AND U23596 ( .A(a[25]), .B(b[82]), .Z(n13905) );
  XNOR U23597 ( .A(n13910), .B(n13273), .Z(n13275) );
  XOR U23598 ( .A(n13911), .B(n13912), .Z(n13273) );
  ANDN U23599 ( .B(n13913), .A(n13914), .Z(n13911) );
  AND U23600 ( .A(a[26]), .B(b[81]), .Z(n13910) );
  XNOR U23601 ( .A(n13915), .B(n13278), .Z(n13280) );
  XOR U23602 ( .A(n13916), .B(n13917), .Z(n13278) );
  ANDN U23603 ( .B(n13918), .A(n13919), .Z(n13916) );
  AND U23604 ( .A(a[27]), .B(b[80]), .Z(n13915) );
  XNOR U23605 ( .A(n13920), .B(n13283), .Z(n13285) );
  XOR U23606 ( .A(n13921), .B(n13922), .Z(n13283) );
  ANDN U23607 ( .B(n13923), .A(n13924), .Z(n13921) );
  AND U23608 ( .A(a[28]), .B(b[79]), .Z(n13920) );
  XNOR U23609 ( .A(n13925), .B(n13288), .Z(n13290) );
  XOR U23610 ( .A(n13926), .B(n13927), .Z(n13288) );
  ANDN U23611 ( .B(n13928), .A(n13929), .Z(n13926) );
  AND U23612 ( .A(a[29]), .B(b[78]), .Z(n13925) );
  XNOR U23613 ( .A(n13930), .B(n13293), .Z(n13295) );
  XOR U23614 ( .A(n13931), .B(n13932), .Z(n13293) );
  ANDN U23615 ( .B(n13933), .A(n13934), .Z(n13931) );
  AND U23616 ( .A(a[30]), .B(b[77]), .Z(n13930) );
  XNOR U23617 ( .A(n13935), .B(n13298), .Z(n13300) );
  XOR U23618 ( .A(n13936), .B(n13937), .Z(n13298) );
  ANDN U23619 ( .B(n13938), .A(n13939), .Z(n13936) );
  AND U23620 ( .A(a[31]), .B(b[76]), .Z(n13935) );
  XNOR U23621 ( .A(n13940), .B(n13303), .Z(n13305) );
  XOR U23622 ( .A(n13941), .B(n13942), .Z(n13303) );
  ANDN U23623 ( .B(n13943), .A(n13944), .Z(n13941) );
  AND U23624 ( .A(a[32]), .B(b[75]), .Z(n13940) );
  XNOR U23625 ( .A(n13945), .B(n13308), .Z(n13310) );
  XOR U23626 ( .A(n13946), .B(n13947), .Z(n13308) );
  ANDN U23627 ( .B(n13948), .A(n13949), .Z(n13946) );
  AND U23628 ( .A(a[33]), .B(b[74]), .Z(n13945) );
  XNOR U23629 ( .A(n13950), .B(n13313), .Z(n13315) );
  XOR U23630 ( .A(n13951), .B(n13952), .Z(n13313) );
  ANDN U23631 ( .B(n13953), .A(n13954), .Z(n13951) );
  AND U23632 ( .A(a[34]), .B(b[73]), .Z(n13950) );
  XNOR U23633 ( .A(n13955), .B(n13318), .Z(n13320) );
  XOR U23634 ( .A(n13956), .B(n13957), .Z(n13318) );
  ANDN U23635 ( .B(n13958), .A(n13959), .Z(n13956) );
  AND U23636 ( .A(a[35]), .B(b[72]), .Z(n13955) );
  XNOR U23637 ( .A(n13960), .B(n13323), .Z(n13325) );
  XOR U23638 ( .A(n13961), .B(n13962), .Z(n13323) );
  ANDN U23639 ( .B(n13963), .A(n13964), .Z(n13961) );
  AND U23640 ( .A(a[36]), .B(b[71]), .Z(n13960) );
  XNOR U23641 ( .A(n13965), .B(n13328), .Z(n13330) );
  XOR U23642 ( .A(n13966), .B(n13967), .Z(n13328) );
  ANDN U23643 ( .B(n13968), .A(n13969), .Z(n13966) );
  AND U23644 ( .A(a[37]), .B(b[70]), .Z(n13965) );
  XNOR U23645 ( .A(n13970), .B(n13333), .Z(n13335) );
  XOR U23646 ( .A(n13971), .B(n13972), .Z(n13333) );
  ANDN U23647 ( .B(n13973), .A(n13974), .Z(n13971) );
  AND U23648 ( .A(a[38]), .B(b[69]), .Z(n13970) );
  XNOR U23649 ( .A(n13975), .B(n13338), .Z(n13340) );
  XOR U23650 ( .A(n13976), .B(n13977), .Z(n13338) );
  ANDN U23651 ( .B(n13978), .A(n13979), .Z(n13976) );
  AND U23652 ( .A(a[39]), .B(b[68]), .Z(n13975) );
  XNOR U23653 ( .A(n13980), .B(n13343), .Z(n13345) );
  XOR U23654 ( .A(n13981), .B(n13982), .Z(n13343) );
  ANDN U23655 ( .B(n13983), .A(n13984), .Z(n13981) );
  AND U23656 ( .A(a[40]), .B(b[67]), .Z(n13980) );
  XNOR U23657 ( .A(n13985), .B(n13348), .Z(n13350) );
  XOR U23658 ( .A(n13986), .B(n13987), .Z(n13348) );
  ANDN U23659 ( .B(n13988), .A(n13989), .Z(n13986) );
  AND U23660 ( .A(a[41]), .B(b[66]), .Z(n13985) );
  XNOR U23661 ( .A(n13990), .B(n13353), .Z(n13355) );
  XOR U23662 ( .A(n13991), .B(n13992), .Z(n13353) );
  ANDN U23663 ( .B(n13993), .A(n13994), .Z(n13991) );
  AND U23664 ( .A(a[42]), .B(b[65]), .Z(n13990) );
  XNOR U23665 ( .A(n13995), .B(n13358), .Z(n13360) );
  XOR U23666 ( .A(n13996), .B(n13997), .Z(n13358) );
  ANDN U23667 ( .B(n13998), .A(n13999), .Z(n13996) );
  AND U23668 ( .A(a[43]), .B(b[64]), .Z(n13995) );
  XNOR U23669 ( .A(n14000), .B(n13363), .Z(n13365) );
  XOR U23670 ( .A(n14001), .B(n14002), .Z(n13363) );
  ANDN U23671 ( .B(n14003), .A(n14004), .Z(n14001) );
  AND U23672 ( .A(a[44]), .B(b[63]), .Z(n14000) );
  XNOR U23673 ( .A(n14005), .B(n13368), .Z(n13370) );
  XOR U23674 ( .A(n14006), .B(n14007), .Z(n13368) );
  ANDN U23675 ( .B(n14008), .A(n14009), .Z(n14006) );
  AND U23676 ( .A(a[45]), .B(b[62]), .Z(n14005) );
  XNOR U23677 ( .A(n14010), .B(n13373), .Z(n13375) );
  XOR U23678 ( .A(n14011), .B(n14012), .Z(n13373) );
  ANDN U23679 ( .B(n14013), .A(n14014), .Z(n14011) );
  AND U23680 ( .A(a[46]), .B(b[61]), .Z(n14010) );
  XNOR U23681 ( .A(n14015), .B(n13378), .Z(n13380) );
  XOR U23682 ( .A(n14016), .B(n14017), .Z(n13378) );
  ANDN U23683 ( .B(n14018), .A(n14019), .Z(n14016) );
  AND U23684 ( .A(a[47]), .B(b[60]), .Z(n14015) );
  XNOR U23685 ( .A(n14020), .B(n13383), .Z(n13385) );
  XOR U23686 ( .A(n14021), .B(n14022), .Z(n13383) );
  ANDN U23687 ( .B(n14023), .A(n14024), .Z(n14021) );
  AND U23688 ( .A(a[48]), .B(b[59]), .Z(n14020) );
  XNOR U23689 ( .A(n14025), .B(n13388), .Z(n13390) );
  XOR U23690 ( .A(n14026), .B(n14027), .Z(n13388) );
  ANDN U23691 ( .B(n14028), .A(n14029), .Z(n14026) );
  AND U23692 ( .A(a[49]), .B(b[58]), .Z(n14025) );
  XNOR U23693 ( .A(n14030), .B(n13393), .Z(n13395) );
  XOR U23694 ( .A(n14031), .B(n14032), .Z(n13393) );
  ANDN U23695 ( .B(n14033), .A(n14034), .Z(n14031) );
  AND U23696 ( .A(a[50]), .B(b[57]), .Z(n14030) );
  XNOR U23697 ( .A(n14035), .B(n13398), .Z(n13400) );
  XOR U23698 ( .A(n14036), .B(n14037), .Z(n13398) );
  ANDN U23699 ( .B(n14038), .A(n14039), .Z(n14036) );
  AND U23700 ( .A(a[51]), .B(b[56]), .Z(n14035) );
  XNOR U23701 ( .A(n14040), .B(n13403), .Z(n13405) );
  XOR U23702 ( .A(n14041), .B(n14042), .Z(n13403) );
  ANDN U23703 ( .B(n14043), .A(n14044), .Z(n14041) );
  AND U23704 ( .A(a[52]), .B(b[55]), .Z(n14040) );
  XNOR U23705 ( .A(n14045), .B(n13408), .Z(n13410) );
  XOR U23706 ( .A(n14046), .B(n14047), .Z(n13408) );
  ANDN U23707 ( .B(n14048), .A(n14049), .Z(n14046) );
  AND U23708 ( .A(a[53]), .B(b[54]), .Z(n14045) );
  XNOR U23709 ( .A(n14050), .B(n13413), .Z(n13415) );
  XOR U23710 ( .A(n14051), .B(n14052), .Z(n13413) );
  ANDN U23711 ( .B(n14053), .A(n14054), .Z(n14051) );
  AND U23712 ( .A(a[54]), .B(b[53]), .Z(n14050) );
  XNOR U23713 ( .A(n14055), .B(n13418), .Z(n13420) );
  XOR U23714 ( .A(n14056), .B(n14057), .Z(n13418) );
  ANDN U23715 ( .B(n14058), .A(n14059), .Z(n14056) );
  AND U23716 ( .A(a[55]), .B(b[52]), .Z(n14055) );
  XNOR U23717 ( .A(n14060), .B(n13423), .Z(n13425) );
  XOR U23718 ( .A(n14061), .B(n14062), .Z(n13423) );
  ANDN U23719 ( .B(n14063), .A(n14064), .Z(n14061) );
  AND U23720 ( .A(a[56]), .B(b[51]), .Z(n14060) );
  XNOR U23721 ( .A(n14065), .B(n13428), .Z(n13430) );
  XOR U23722 ( .A(n14066), .B(n14067), .Z(n13428) );
  ANDN U23723 ( .B(n14068), .A(n14069), .Z(n14066) );
  AND U23724 ( .A(a[57]), .B(b[50]), .Z(n14065) );
  XNOR U23725 ( .A(n14070), .B(n13433), .Z(n13435) );
  XOR U23726 ( .A(n14071), .B(n14072), .Z(n13433) );
  ANDN U23727 ( .B(n14073), .A(n14074), .Z(n14071) );
  AND U23728 ( .A(a[58]), .B(b[49]), .Z(n14070) );
  XNOR U23729 ( .A(n14075), .B(n13438), .Z(n13440) );
  XOR U23730 ( .A(n14076), .B(n14077), .Z(n13438) );
  ANDN U23731 ( .B(n14078), .A(n14079), .Z(n14076) );
  AND U23732 ( .A(a[59]), .B(b[48]), .Z(n14075) );
  XNOR U23733 ( .A(n14080), .B(n13443), .Z(n13445) );
  XOR U23734 ( .A(n14081), .B(n14082), .Z(n13443) );
  ANDN U23735 ( .B(n14083), .A(n14084), .Z(n14081) );
  AND U23736 ( .A(a[60]), .B(b[47]), .Z(n14080) );
  XNOR U23737 ( .A(n14085), .B(n13448), .Z(n13450) );
  XOR U23738 ( .A(n14086), .B(n14087), .Z(n13448) );
  ANDN U23739 ( .B(n14088), .A(n14089), .Z(n14086) );
  AND U23740 ( .A(a[61]), .B(b[46]), .Z(n14085) );
  XNOR U23741 ( .A(n14090), .B(n13453), .Z(n13455) );
  XOR U23742 ( .A(n14091), .B(n14092), .Z(n13453) );
  ANDN U23743 ( .B(n14093), .A(n14094), .Z(n14091) );
  AND U23744 ( .A(a[62]), .B(b[45]), .Z(n14090) );
  XNOR U23745 ( .A(n14095), .B(n13458), .Z(n13460) );
  XOR U23746 ( .A(n14096), .B(n14097), .Z(n13458) );
  ANDN U23747 ( .B(n14098), .A(n14099), .Z(n14096) );
  AND U23748 ( .A(a[63]), .B(b[44]), .Z(n14095) );
  XNOR U23749 ( .A(n14100), .B(n13463), .Z(n13465) );
  XOR U23750 ( .A(n14101), .B(n14102), .Z(n13463) );
  ANDN U23751 ( .B(n14103), .A(n14104), .Z(n14101) );
  AND U23752 ( .A(a[64]), .B(b[43]), .Z(n14100) );
  XNOR U23753 ( .A(n14105), .B(n13468), .Z(n13470) );
  XOR U23754 ( .A(n14106), .B(n14107), .Z(n13468) );
  ANDN U23755 ( .B(n14108), .A(n14109), .Z(n14106) );
  AND U23756 ( .A(a[65]), .B(b[42]), .Z(n14105) );
  XNOR U23757 ( .A(n14110), .B(n13473), .Z(n13475) );
  XOR U23758 ( .A(n14111), .B(n14112), .Z(n13473) );
  ANDN U23759 ( .B(n14113), .A(n14114), .Z(n14111) );
  AND U23760 ( .A(a[66]), .B(b[41]), .Z(n14110) );
  XNOR U23761 ( .A(n14115), .B(n13478), .Z(n13480) );
  XOR U23762 ( .A(n14116), .B(n14117), .Z(n13478) );
  ANDN U23763 ( .B(n14118), .A(n14119), .Z(n14116) );
  AND U23764 ( .A(a[67]), .B(b[40]), .Z(n14115) );
  XNOR U23765 ( .A(n14120), .B(n13483), .Z(n13485) );
  XOR U23766 ( .A(n14121), .B(n14122), .Z(n13483) );
  ANDN U23767 ( .B(n14123), .A(n14124), .Z(n14121) );
  AND U23768 ( .A(a[68]), .B(b[39]), .Z(n14120) );
  XNOR U23769 ( .A(n14125), .B(n13488), .Z(n13490) );
  XOR U23770 ( .A(n14126), .B(n14127), .Z(n13488) );
  ANDN U23771 ( .B(n14128), .A(n14129), .Z(n14126) );
  AND U23772 ( .A(a[69]), .B(b[38]), .Z(n14125) );
  XNOR U23773 ( .A(n14130), .B(n13493), .Z(n13495) );
  XOR U23774 ( .A(n14131), .B(n14132), .Z(n13493) );
  ANDN U23775 ( .B(n14133), .A(n14134), .Z(n14131) );
  AND U23776 ( .A(a[70]), .B(b[37]), .Z(n14130) );
  XNOR U23777 ( .A(n14135), .B(n13498), .Z(n13500) );
  XOR U23778 ( .A(n14136), .B(n14137), .Z(n13498) );
  ANDN U23779 ( .B(n14138), .A(n14139), .Z(n14136) );
  AND U23780 ( .A(a[71]), .B(b[36]), .Z(n14135) );
  XNOR U23781 ( .A(n14140), .B(n13503), .Z(n13505) );
  XOR U23782 ( .A(n14141), .B(n14142), .Z(n13503) );
  ANDN U23783 ( .B(n14143), .A(n14144), .Z(n14141) );
  AND U23784 ( .A(a[72]), .B(b[35]), .Z(n14140) );
  XNOR U23785 ( .A(n14145), .B(n13508), .Z(n13510) );
  XOR U23786 ( .A(n14146), .B(n14147), .Z(n13508) );
  ANDN U23787 ( .B(n14148), .A(n14149), .Z(n14146) );
  AND U23788 ( .A(a[73]), .B(b[34]), .Z(n14145) );
  XNOR U23789 ( .A(n14150), .B(n13513), .Z(n13515) );
  XOR U23790 ( .A(n14151), .B(n14152), .Z(n13513) );
  ANDN U23791 ( .B(n14153), .A(n14154), .Z(n14151) );
  AND U23792 ( .A(a[74]), .B(b[33]), .Z(n14150) );
  XNOR U23793 ( .A(n14155), .B(n13518), .Z(n13520) );
  XOR U23794 ( .A(n14156), .B(n14157), .Z(n13518) );
  ANDN U23795 ( .B(n14158), .A(n14159), .Z(n14156) );
  AND U23796 ( .A(a[75]), .B(b[32]), .Z(n14155) );
  XNOR U23797 ( .A(n14160), .B(n13523), .Z(n13525) );
  XOR U23798 ( .A(n14161), .B(n14162), .Z(n13523) );
  ANDN U23799 ( .B(n14163), .A(n14164), .Z(n14161) );
  AND U23800 ( .A(a[76]), .B(b[31]), .Z(n14160) );
  XNOR U23801 ( .A(n14165), .B(n13528), .Z(n13530) );
  XOR U23802 ( .A(n14166), .B(n14167), .Z(n13528) );
  ANDN U23803 ( .B(n14168), .A(n14169), .Z(n14166) );
  AND U23804 ( .A(a[77]), .B(b[30]), .Z(n14165) );
  XNOR U23805 ( .A(n14170), .B(n13533), .Z(n13535) );
  XOR U23806 ( .A(n14171), .B(n14172), .Z(n13533) );
  ANDN U23807 ( .B(n14173), .A(n14174), .Z(n14171) );
  AND U23808 ( .A(a[78]), .B(b[29]), .Z(n14170) );
  XNOR U23809 ( .A(n14175), .B(n13538), .Z(n13540) );
  XOR U23810 ( .A(n14176), .B(n14177), .Z(n13538) );
  ANDN U23811 ( .B(n14178), .A(n14179), .Z(n14176) );
  AND U23812 ( .A(a[79]), .B(b[28]), .Z(n14175) );
  XNOR U23813 ( .A(n14180), .B(n13543), .Z(n13545) );
  XOR U23814 ( .A(n14181), .B(n14182), .Z(n13543) );
  ANDN U23815 ( .B(n14183), .A(n14184), .Z(n14181) );
  AND U23816 ( .A(a[80]), .B(b[27]), .Z(n14180) );
  XNOR U23817 ( .A(n14185), .B(n13548), .Z(n13550) );
  XOR U23818 ( .A(n14186), .B(n14187), .Z(n13548) );
  ANDN U23819 ( .B(n14188), .A(n14189), .Z(n14186) );
  AND U23820 ( .A(a[81]), .B(b[26]), .Z(n14185) );
  XNOR U23821 ( .A(n14190), .B(n13553), .Z(n13555) );
  XOR U23822 ( .A(n14191), .B(n14192), .Z(n13553) );
  ANDN U23823 ( .B(n14193), .A(n14194), .Z(n14191) );
  AND U23824 ( .A(a[82]), .B(b[25]), .Z(n14190) );
  XNOR U23825 ( .A(n14195), .B(n13558), .Z(n13560) );
  XOR U23826 ( .A(n14196), .B(n14197), .Z(n13558) );
  ANDN U23827 ( .B(n14198), .A(n14199), .Z(n14196) );
  AND U23828 ( .A(a[83]), .B(b[24]), .Z(n14195) );
  XNOR U23829 ( .A(n14200), .B(n13563), .Z(n13565) );
  XOR U23830 ( .A(n14201), .B(n14202), .Z(n13563) );
  ANDN U23831 ( .B(n14203), .A(n14204), .Z(n14201) );
  AND U23832 ( .A(a[84]), .B(b[23]), .Z(n14200) );
  XNOR U23833 ( .A(n14205), .B(n13568), .Z(n13570) );
  XOR U23834 ( .A(n14206), .B(n14207), .Z(n13568) );
  ANDN U23835 ( .B(n14208), .A(n14209), .Z(n14206) );
  AND U23836 ( .A(a[85]), .B(b[22]), .Z(n14205) );
  XNOR U23837 ( .A(n14210), .B(n13573), .Z(n13575) );
  XOR U23838 ( .A(n14211), .B(n14212), .Z(n13573) );
  ANDN U23839 ( .B(n14213), .A(n14214), .Z(n14211) );
  AND U23840 ( .A(a[86]), .B(b[21]), .Z(n14210) );
  XNOR U23841 ( .A(n14215), .B(n13578), .Z(n13580) );
  XOR U23842 ( .A(n14216), .B(n14217), .Z(n13578) );
  ANDN U23843 ( .B(n14218), .A(n14219), .Z(n14216) );
  AND U23844 ( .A(a[87]), .B(b[20]), .Z(n14215) );
  XNOR U23845 ( .A(n14220), .B(n13583), .Z(n13585) );
  XOR U23846 ( .A(n14221), .B(n14222), .Z(n13583) );
  ANDN U23847 ( .B(n14223), .A(n14224), .Z(n14221) );
  AND U23848 ( .A(a[88]), .B(b[19]), .Z(n14220) );
  XNOR U23849 ( .A(n14225), .B(n13588), .Z(n13590) );
  XOR U23850 ( .A(n14226), .B(n14227), .Z(n13588) );
  ANDN U23851 ( .B(n14228), .A(n14229), .Z(n14226) );
  AND U23852 ( .A(a[89]), .B(b[18]), .Z(n14225) );
  XNOR U23853 ( .A(n14230), .B(n13593), .Z(n13595) );
  XOR U23854 ( .A(n14231), .B(n14232), .Z(n13593) );
  ANDN U23855 ( .B(n14233), .A(n14234), .Z(n14231) );
  AND U23856 ( .A(a[90]), .B(b[17]), .Z(n14230) );
  XNOR U23857 ( .A(n14235), .B(n13598), .Z(n13600) );
  XOR U23858 ( .A(n14236), .B(n14237), .Z(n13598) );
  ANDN U23859 ( .B(n14238), .A(n14239), .Z(n14236) );
  AND U23860 ( .A(a[91]), .B(b[16]), .Z(n14235) );
  XNOR U23861 ( .A(n14240), .B(n13603), .Z(n13605) );
  XOR U23862 ( .A(n14241), .B(n14242), .Z(n13603) );
  ANDN U23863 ( .B(n14243), .A(n14244), .Z(n14241) );
  AND U23864 ( .A(a[92]), .B(b[15]), .Z(n14240) );
  XNOR U23865 ( .A(n14245), .B(n13608), .Z(n13610) );
  XOR U23866 ( .A(n14246), .B(n14247), .Z(n13608) );
  ANDN U23867 ( .B(n14248), .A(n14249), .Z(n14246) );
  AND U23868 ( .A(a[93]), .B(b[14]), .Z(n14245) );
  XNOR U23869 ( .A(n14250), .B(n13613), .Z(n13615) );
  XOR U23870 ( .A(n14251), .B(n14252), .Z(n13613) );
  ANDN U23871 ( .B(n14253), .A(n14254), .Z(n14251) );
  AND U23872 ( .A(a[94]), .B(b[13]), .Z(n14250) );
  XNOR U23873 ( .A(n14255), .B(n13618), .Z(n13620) );
  XOR U23874 ( .A(n14256), .B(n14257), .Z(n13618) );
  ANDN U23875 ( .B(n14258), .A(n14259), .Z(n14256) );
  AND U23876 ( .A(a[95]), .B(b[12]), .Z(n14255) );
  XNOR U23877 ( .A(n14260), .B(n13623), .Z(n13625) );
  XOR U23878 ( .A(n14261), .B(n14262), .Z(n13623) );
  ANDN U23879 ( .B(n14263), .A(n14264), .Z(n14261) );
  AND U23880 ( .A(a[96]), .B(b[11]), .Z(n14260) );
  XNOR U23881 ( .A(n14265), .B(n13628), .Z(n13630) );
  XOR U23882 ( .A(n14266), .B(n14267), .Z(n13628) );
  ANDN U23883 ( .B(n14268), .A(n14269), .Z(n14266) );
  AND U23884 ( .A(a[97]), .B(b[10]), .Z(n14265) );
  XNOR U23885 ( .A(n14270), .B(n13633), .Z(n13635) );
  XOR U23886 ( .A(n14271), .B(n14272), .Z(n13633) );
  ANDN U23887 ( .B(n14273), .A(n14274), .Z(n14271) );
  AND U23888 ( .A(b[9]), .B(a[98]), .Z(n14270) );
  XNOR U23889 ( .A(n14275), .B(n13638), .Z(n13640) );
  XOR U23890 ( .A(n14276), .B(n14277), .Z(n13638) );
  ANDN U23891 ( .B(n14278), .A(n14279), .Z(n14276) );
  AND U23892 ( .A(b[8]), .B(a[99]), .Z(n14275) );
  XNOR U23893 ( .A(n14280), .B(n13643), .Z(n13645) );
  XOR U23894 ( .A(n14281), .B(n14282), .Z(n13643) );
  ANDN U23895 ( .B(n14283), .A(n14284), .Z(n14281) );
  AND U23896 ( .A(b[7]), .B(a[100]), .Z(n14280) );
  XNOR U23897 ( .A(n14285), .B(n13648), .Z(n13650) );
  XOR U23898 ( .A(n14286), .B(n14287), .Z(n13648) );
  ANDN U23899 ( .B(n14288), .A(n14289), .Z(n14286) );
  AND U23900 ( .A(b[6]), .B(a[101]), .Z(n14285) );
  XNOR U23901 ( .A(n14290), .B(n13653), .Z(n13655) );
  XOR U23902 ( .A(n14291), .B(n14292), .Z(n13653) );
  ANDN U23903 ( .B(n14293), .A(n14294), .Z(n14291) );
  AND U23904 ( .A(b[5]), .B(a[102]), .Z(n14290) );
  XNOR U23905 ( .A(n14295), .B(n13658), .Z(n13660) );
  XOR U23906 ( .A(n14296), .B(n14297), .Z(n13658) );
  ANDN U23907 ( .B(n14298), .A(n14299), .Z(n14296) );
  AND U23908 ( .A(b[4]), .B(a[103]), .Z(n14295) );
  XNOR U23909 ( .A(n14300), .B(n14301), .Z(n13672) );
  NANDN U23910 ( .A(n14302), .B(n14303), .Z(n14301) );
  XNOR U23911 ( .A(n14304), .B(n13663), .Z(n13665) );
  XNOR U23912 ( .A(n14305), .B(n14306), .Z(n13663) );
  AND U23913 ( .A(n14307), .B(n14308), .Z(n14305) );
  AND U23914 ( .A(b[3]), .B(a[104]), .Z(n14304) );
  NAND U23915 ( .A(a[107]), .B(b[0]), .Z(n13038) );
  XNOR U23916 ( .A(n13678), .B(n13679), .Z(c[106]) );
  XNOR U23917 ( .A(n14302), .B(n14303), .Z(n13679) );
  XOR U23918 ( .A(n14300), .B(n14309), .Z(n14303) );
  NAND U23919 ( .A(b[1]), .B(a[105]), .Z(n14309) );
  XOR U23920 ( .A(n14308), .B(n14310), .Z(n14302) );
  XOR U23921 ( .A(n14300), .B(n14307), .Z(n14310) );
  XNOR U23922 ( .A(n14311), .B(n14306), .Z(n14307) );
  AND U23923 ( .A(b[2]), .B(a[104]), .Z(n14311) );
  NANDN U23924 ( .A(n14312), .B(n14313), .Z(n14300) );
  XOR U23925 ( .A(n14306), .B(n14298), .Z(n14314) );
  XNOR U23926 ( .A(n14297), .B(n14293), .Z(n14315) );
  XNOR U23927 ( .A(n14292), .B(n14288), .Z(n14316) );
  XNOR U23928 ( .A(n14287), .B(n14283), .Z(n14317) );
  XNOR U23929 ( .A(n14282), .B(n14278), .Z(n14318) );
  XNOR U23930 ( .A(n14277), .B(n14273), .Z(n14319) );
  XNOR U23931 ( .A(n14272), .B(n14268), .Z(n14320) );
  XNOR U23932 ( .A(n14267), .B(n14263), .Z(n14321) );
  XNOR U23933 ( .A(n14262), .B(n14258), .Z(n14322) );
  XNOR U23934 ( .A(n14257), .B(n14253), .Z(n14323) );
  XNOR U23935 ( .A(n14252), .B(n14248), .Z(n14324) );
  XNOR U23936 ( .A(n14247), .B(n14243), .Z(n14325) );
  XNOR U23937 ( .A(n14242), .B(n14238), .Z(n14326) );
  XNOR U23938 ( .A(n14237), .B(n14233), .Z(n14327) );
  XNOR U23939 ( .A(n14232), .B(n14228), .Z(n14328) );
  XNOR U23940 ( .A(n14227), .B(n14223), .Z(n14329) );
  XNOR U23941 ( .A(n14222), .B(n14218), .Z(n14330) );
  XNOR U23942 ( .A(n14217), .B(n14213), .Z(n14331) );
  XNOR U23943 ( .A(n14212), .B(n14208), .Z(n14332) );
  XNOR U23944 ( .A(n14207), .B(n14203), .Z(n14333) );
  XNOR U23945 ( .A(n14202), .B(n14198), .Z(n14334) );
  XNOR U23946 ( .A(n14197), .B(n14193), .Z(n14335) );
  XNOR U23947 ( .A(n14192), .B(n14188), .Z(n14336) );
  XNOR U23948 ( .A(n14187), .B(n14183), .Z(n14337) );
  XNOR U23949 ( .A(n14182), .B(n14178), .Z(n14338) );
  XNOR U23950 ( .A(n14177), .B(n14173), .Z(n14339) );
  XNOR U23951 ( .A(n14172), .B(n14168), .Z(n14340) );
  XNOR U23952 ( .A(n14167), .B(n14163), .Z(n14341) );
  XNOR U23953 ( .A(n14162), .B(n14158), .Z(n14342) );
  XNOR U23954 ( .A(n14157), .B(n14153), .Z(n14343) );
  XNOR U23955 ( .A(n14152), .B(n14148), .Z(n14344) );
  XNOR U23956 ( .A(n14147), .B(n14143), .Z(n14345) );
  XNOR U23957 ( .A(n14142), .B(n14138), .Z(n14346) );
  XNOR U23958 ( .A(n14137), .B(n14133), .Z(n14347) );
  XNOR U23959 ( .A(n14132), .B(n14128), .Z(n14348) );
  XNOR U23960 ( .A(n14127), .B(n14123), .Z(n14349) );
  XNOR U23961 ( .A(n14122), .B(n14118), .Z(n14350) );
  XNOR U23962 ( .A(n14117), .B(n14113), .Z(n14351) );
  XNOR U23963 ( .A(n14112), .B(n14108), .Z(n14352) );
  XNOR U23964 ( .A(n14107), .B(n14103), .Z(n14353) );
  XNOR U23965 ( .A(n14102), .B(n14098), .Z(n14354) );
  XNOR U23966 ( .A(n14097), .B(n14093), .Z(n14355) );
  XNOR U23967 ( .A(n14092), .B(n14088), .Z(n14356) );
  XNOR U23968 ( .A(n14087), .B(n14083), .Z(n14357) );
  XNOR U23969 ( .A(n14082), .B(n14078), .Z(n14358) );
  XNOR U23970 ( .A(n14077), .B(n14073), .Z(n14359) );
  XNOR U23971 ( .A(n14072), .B(n14068), .Z(n14360) );
  XNOR U23972 ( .A(n14067), .B(n14063), .Z(n14361) );
  XNOR U23973 ( .A(n14062), .B(n14058), .Z(n14362) );
  XNOR U23974 ( .A(n14057), .B(n14053), .Z(n14363) );
  XNOR U23975 ( .A(n14052), .B(n14048), .Z(n14364) );
  XNOR U23976 ( .A(n14047), .B(n14043), .Z(n14365) );
  XNOR U23977 ( .A(n14042), .B(n14038), .Z(n14366) );
  XNOR U23978 ( .A(n14037), .B(n14033), .Z(n14367) );
  XNOR U23979 ( .A(n14032), .B(n14028), .Z(n14368) );
  XNOR U23980 ( .A(n14027), .B(n14023), .Z(n14369) );
  XNOR U23981 ( .A(n14022), .B(n14018), .Z(n14370) );
  XNOR U23982 ( .A(n14017), .B(n14013), .Z(n14371) );
  XNOR U23983 ( .A(n14012), .B(n14008), .Z(n14372) );
  XNOR U23984 ( .A(n14007), .B(n14003), .Z(n14373) );
  XNOR U23985 ( .A(n14002), .B(n13998), .Z(n14374) );
  XNOR U23986 ( .A(n13997), .B(n13993), .Z(n14375) );
  XNOR U23987 ( .A(n13992), .B(n13988), .Z(n14376) );
  XNOR U23988 ( .A(n13987), .B(n13983), .Z(n14377) );
  XNOR U23989 ( .A(n13982), .B(n13978), .Z(n14378) );
  XNOR U23990 ( .A(n13977), .B(n13973), .Z(n14379) );
  XNOR U23991 ( .A(n13972), .B(n13968), .Z(n14380) );
  XNOR U23992 ( .A(n13967), .B(n13963), .Z(n14381) );
  XNOR U23993 ( .A(n13962), .B(n13958), .Z(n14382) );
  XNOR U23994 ( .A(n13957), .B(n13953), .Z(n14383) );
  XNOR U23995 ( .A(n13952), .B(n13948), .Z(n14384) );
  XNOR U23996 ( .A(n13947), .B(n13943), .Z(n14385) );
  XNOR U23997 ( .A(n13942), .B(n13938), .Z(n14386) );
  XNOR U23998 ( .A(n13937), .B(n13933), .Z(n14387) );
  XNOR U23999 ( .A(n13932), .B(n13928), .Z(n14388) );
  XNOR U24000 ( .A(n13927), .B(n13923), .Z(n14389) );
  XNOR U24001 ( .A(n13922), .B(n13918), .Z(n14390) );
  XNOR U24002 ( .A(n13917), .B(n13913), .Z(n14391) );
  XNOR U24003 ( .A(n13912), .B(n13908), .Z(n14392) );
  XNOR U24004 ( .A(n13907), .B(n13903), .Z(n14393) );
  XNOR U24005 ( .A(n13902), .B(n13898), .Z(n14394) );
  XNOR U24006 ( .A(n13897), .B(n13893), .Z(n14395) );
  XNOR U24007 ( .A(n13892), .B(n13888), .Z(n14396) );
  XNOR U24008 ( .A(n13887), .B(n13883), .Z(n14397) );
  XNOR U24009 ( .A(n13882), .B(n13878), .Z(n14398) );
  XNOR U24010 ( .A(n13877), .B(n13873), .Z(n14399) );
  XNOR U24011 ( .A(n13872), .B(n13868), .Z(n14400) );
  XNOR U24012 ( .A(n13867), .B(n13863), .Z(n14401) );
  XNOR U24013 ( .A(n13862), .B(n13858), .Z(n14402) );
  XNOR U24014 ( .A(n13857), .B(n13853), .Z(n14403) );
  XNOR U24015 ( .A(n13852), .B(n13848), .Z(n14404) );
  XNOR U24016 ( .A(n13847), .B(n13843), .Z(n14405) );
  XNOR U24017 ( .A(n13842), .B(n13838), .Z(n14406) );
  XNOR U24018 ( .A(n13837), .B(n13833), .Z(n14407) );
  XNOR U24019 ( .A(n13832), .B(n13828), .Z(n14408) );
  XNOR U24020 ( .A(n13827), .B(n13823), .Z(n14409) );
  XNOR U24021 ( .A(n13822), .B(n13818), .Z(n14410) );
  XNOR U24022 ( .A(n13817), .B(n13813), .Z(n14411) );
  XNOR U24023 ( .A(n13812), .B(n13808), .Z(n14412) );
  XNOR U24024 ( .A(n13807), .B(n13803), .Z(n14413) );
  XNOR U24025 ( .A(n13802), .B(n13798), .Z(n14414) );
  XNOR U24026 ( .A(n13797), .B(n13793), .Z(n14415) );
  XNOR U24027 ( .A(n13792), .B(n13788), .Z(n14416) );
  XOR U24028 ( .A(n14417), .B(n13787), .Z(n13788) );
  AND U24029 ( .A(a[0]), .B(b[106]), .Z(n14417) );
  XNOR U24030 ( .A(n14418), .B(n13787), .Z(n13789) );
  XNOR U24031 ( .A(n14419), .B(n14420), .Z(n13787) );
  ANDN U24032 ( .B(n14421), .A(n14422), .Z(n14419) );
  AND U24033 ( .A(a[1]), .B(b[105]), .Z(n14418) );
  XNOR U24034 ( .A(n14423), .B(n13792), .Z(n13794) );
  XOR U24035 ( .A(n14424), .B(n14425), .Z(n13792) );
  ANDN U24036 ( .B(n14426), .A(n14427), .Z(n14424) );
  AND U24037 ( .A(a[2]), .B(b[104]), .Z(n14423) );
  XNOR U24038 ( .A(n14428), .B(n13797), .Z(n13799) );
  XOR U24039 ( .A(n14429), .B(n14430), .Z(n13797) );
  ANDN U24040 ( .B(n14431), .A(n14432), .Z(n14429) );
  AND U24041 ( .A(a[3]), .B(b[103]), .Z(n14428) );
  XNOR U24042 ( .A(n14433), .B(n13802), .Z(n13804) );
  XOR U24043 ( .A(n14434), .B(n14435), .Z(n13802) );
  ANDN U24044 ( .B(n14436), .A(n14437), .Z(n14434) );
  AND U24045 ( .A(a[4]), .B(b[102]), .Z(n14433) );
  XNOR U24046 ( .A(n14438), .B(n13807), .Z(n13809) );
  XOR U24047 ( .A(n14439), .B(n14440), .Z(n13807) );
  ANDN U24048 ( .B(n14441), .A(n14442), .Z(n14439) );
  AND U24049 ( .A(a[5]), .B(b[101]), .Z(n14438) );
  XNOR U24050 ( .A(n14443), .B(n13812), .Z(n13814) );
  XOR U24051 ( .A(n14444), .B(n14445), .Z(n13812) );
  ANDN U24052 ( .B(n14446), .A(n14447), .Z(n14444) );
  AND U24053 ( .A(a[6]), .B(b[100]), .Z(n14443) );
  XNOR U24054 ( .A(n14448), .B(n13817), .Z(n13819) );
  XOR U24055 ( .A(n14449), .B(n14450), .Z(n13817) );
  ANDN U24056 ( .B(n14451), .A(n14452), .Z(n14449) );
  AND U24057 ( .A(a[7]), .B(b[99]), .Z(n14448) );
  XNOR U24058 ( .A(n14453), .B(n13822), .Z(n13824) );
  XOR U24059 ( .A(n14454), .B(n14455), .Z(n13822) );
  ANDN U24060 ( .B(n14456), .A(n14457), .Z(n14454) );
  AND U24061 ( .A(a[8]), .B(b[98]), .Z(n14453) );
  XNOR U24062 ( .A(n14458), .B(n13827), .Z(n13829) );
  XOR U24063 ( .A(n14459), .B(n14460), .Z(n13827) );
  ANDN U24064 ( .B(n14461), .A(n14462), .Z(n14459) );
  AND U24065 ( .A(a[9]), .B(b[97]), .Z(n14458) );
  XNOR U24066 ( .A(n14463), .B(n13832), .Z(n13834) );
  XOR U24067 ( .A(n14464), .B(n14465), .Z(n13832) );
  ANDN U24068 ( .B(n14466), .A(n14467), .Z(n14464) );
  AND U24069 ( .A(a[10]), .B(b[96]), .Z(n14463) );
  XNOR U24070 ( .A(n14468), .B(n13837), .Z(n13839) );
  XOR U24071 ( .A(n14469), .B(n14470), .Z(n13837) );
  ANDN U24072 ( .B(n14471), .A(n14472), .Z(n14469) );
  AND U24073 ( .A(a[11]), .B(b[95]), .Z(n14468) );
  XNOR U24074 ( .A(n14473), .B(n13842), .Z(n13844) );
  XOR U24075 ( .A(n14474), .B(n14475), .Z(n13842) );
  ANDN U24076 ( .B(n14476), .A(n14477), .Z(n14474) );
  AND U24077 ( .A(a[12]), .B(b[94]), .Z(n14473) );
  XNOR U24078 ( .A(n14478), .B(n13847), .Z(n13849) );
  XOR U24079 ( .A(n14479), .B(n14480), .Z(n13847) );
  ANDN U24080 ( .B(n14481), .A(n14482), .Z(n14479) );
  AND U24081 ( .A(a[13]), .B(b[93]), .Z(n14478) );
  XNOR U24082 ( .A(n14483), .B(n13852), .Z(n13854) );
  XOR U24083 ( .A(n14484), .B(n14485), .Z(n13852) );
  ANDN U24084 ( .B(n14486), .A(n14487), .Z(n14484) );
  AND U24085 ( .A(a[14]), .B(b[92]), .Z(n14483) );
  XNOR U24086 ( .A(n14488), .B(n13857), .Z(n13859) );
  XOR U24087 ( .A(n14489), .B(n14490), .Z(n13857) );
  ANDN U24088 ( .B(n14491), .A(n14492), .Z(n14489) );
  AND U24089 ( .A(a[15]), .B(b[91]), .Z(n14488) );
  XNOR U24090 ( .A(n14493), .B(n13862), .Z(n13864) );
  XOR U24091 ( .A(n14494), .B(n14495), .Z(n13862) );
  ANDN U24092 ( .B(n14496), .A(n14497), .Z(n14494) );
  AND U24093 ( .A(a[16]), .B(b[90]), .Z(n14493) );
  XNOR U24094 ( .A(n14498), .B(n13867), .Z(n13869) );
  XOR U24095 ( .A(n14499), .B(n14500), .Z(n13867) );
  ANDN U24096 ( .B(n14501), .A(n14502), .Z(n14499) );
  AND U24097 ( .A(a[17]), .B(b[89]), .Z(n14498) );
  XNOR U24098 ( .A(n14503), .B(n13872), .Z(n13874) );
  XOR U24099 ( .A(n14504), .B(n14505), .Z(n13872) );
  ANDN U24100 ( .B(n14506), .A(n14507), .Z(n14504) );
  AND U24101 ( .A(a[18]), .B(b[88]), .Z(n14503) );
  XNOR U24102 ( .A(n14508), .B(n13877), .Z(n13879) );
  XOR U24103 ( .A(n14509), .B(n14510), .Z(n13877) );
  ANDN U24104 ( .B(n14511), .A(n14512), .Z(n14509) );
  AND U24105 ( .A(a[19]), .B(b[87]), .Z(n14508) );
  XNOR U24106 ( .A(n14513), .B(n13882), .Z(n13884) );
  XOR U24107 ( .A(n14514), .B(n14515), .Z(n13882) );
  ANDN U24108 ( .B(n14516), .A(n14517), .Z(n14514) );
  AND U24109 ( .A(a[20]), .B(b[86]), .Z(n14513) );
  XNOR U24110 ( .A(n14518), .B(n13887), .Z(n13889) );
  XOR U24111 ( .A(n14519), .B(n14520), .Z(n13887) );
  ANDN U24112 ( .B(n14521), .A(n14522), .Z(n14519) );
  AND U24113 ( .A(a[21]), .B(b[85]), .Z(n14518) );
  XNOR U24114 ( .A(n14523), .B(n13892), .Z(n13894) );
  XOR U24115 ( .A(n14524), .B(n14525), .Z(n13892) );
  ANDN U24116 ( .B(n14526), .A(n14527), .Z(n14524) );
  AND U24117 ( .A(a[22]), .B(b[84]), .Z(n14523) );
  XNOR U24118 ( .A(n14528), .B(n13897), .Z(n13899) );
  XOR U24119 ( .A(n14529), .B(n14530), .Z(n13897) );
  ANDN U24120 ( .B(n14531), .A(n14532), .Z(n14529) );
  AND U24121 ( .A(a[23]), .B(b[83]), .Z(n14528) );
  XNOR U24122 ( .A(n14533), .B(n13902), .Z(n13904) );
  XOR U24123 ( .A(n14534), .B(n14535), .Z(n13902) );
  ANDN U24124 ( .B(n14536), .A(n14537), .Z(n14534) );
  AND U24125 ( .A(a[24]), .B(b[82]), .Z(n14533) );
  XNOR U24126 ( .A(n14538), .B(n13907), .Z(n13909) );
  XOR U24127 ( .A(n14539), .B(n14540), .Z(n13907) );
  ANDN U24128 ( .B(n14541), .A(n14542), .Z(n14539) );
  AND U24129 ( .A(a[25]), .B(b[81]), .Z(n14538) );
  XNOR U24130 ( .A(n14543), .B(n13912), .Z(n13914) );
  XOR U24131 ( .A(n14544), .B(n14545), .Z(n13912) );
  ANDN U24132 ( .B(n14546), .A(n14547), .Z(n14544) );
  AND U24133 ( .A(a[26]), .B(b[80]), .Z(n14543) );
  XNOR U24134 ( .A(n14548), .B(n13917), .Z(n13919) );
  XOR U24135 ( .A(n14549), .B(n14550), .Z(n13917) );
  ANDN U24136 ( .B(n14551), .A(n14552), .Z(n14549) );
  AND U24137 ( .A(a[27]), .B(b[79]), .Z(n14548) );
  XNOR U24138 ( .A(n14553), .B(n13922), .Z(n13924) );
  XOR U24139 ( .A(n14554), .B(n14555), .Z(n13922) );
  ANDN U24140 ( .B(n14556), .A(n14557), .Z(n14554) );
  AND U24141 ( .A(a[28]), .B(b[78]), .Z(n14553) );
  XNOR U24142 ( .A(n14558), .B(n13927), .Z(n13929) );
  XOR U24143 ( .A(n14559), .B(n14560), .Z(n13927) );
  ANDN U24144 ( .B(n14561), .A(n14562), .Z(n14559) );
  AND U24145 ( .A(a[29]), .B(b[77]), .Z(n14558) );
  XNOR U24146 ( .A(n14563), .B(n13932), .Z(n13934) );
  XOR U24147 ( .A(n14564), .B(n14565), .Z(n13932) );
  ANDN U24148 ( .B(n14566), .A(n14567), .Z(n14564) );
  AND U24149 ( .A(a[30]), .B(b[76]), .Z(n14563) );
  XNOR U24150 ( .A(n14568), .B(n13937), .Z(n13939) );
  XOR U24151 ( .A(n14569), .B(n14570), .Z(n13937) );
  ANDN U24152 ( .B(n14571), .A(n14572), .Z(n14569) );
  AND U24153 ( .A(a[31]), .B(b[75]), .Z(n14568) );
  XNOR U24154 ( .A(n14573), .B(n13942), .Z(n13944) );
  XOR U24155 ( .A(n14574), .B(n14575), .Z(n13942) );
  ANDN U24156 ( .B(n14576), .A(n14577), .Z(n14574) );
  AND U24157 ( .A(a[32]), .B(b[74]), .Z(n14573) );
  XNOR U24158 ( .A(n14578), .B(n13947), .Z(n13949) );
  XOR U24159 ( .A(n14579), .B(n14580), .Z(n13947) );
  ANDN U24160 ( .B(n14581), .A(n14582), .Z(n14579) );
  AND U24161 ( .A(a[33]), .B(b[73]), .Z(n14578) );
  XNOR U24162 ( .A(n14583), .B(n13952), .Z(n13954) );
  XOR U24163 ( .A(n14584), .B(n14585), .Z(n13952) );
  ANDN U24164 ( .B(n14586), .A(n14587), .Z(n14584) );
  AND U24165 ( .A(a[34]), .B(b[72]), .Z(n14583) );
  XNOR U24166 ( .A(n14588), .B(n13957), .Z(n13959) );
  XOR U24167 ( .A(n14589), .B(n14590), .Z(n13957) );
  ANDN U24168 ( .B(n14591), .A(n14592), .Z(n14589) );
  AND U24169 ( .A(a[35]), .B(b[71]), .Z(n14588) );
  XNOR U24170 ( .A(n14593), .B(n13962), .Z(n13964) );
  XOR U24171 ( .A(n14594), .B(n14595), .Z(n13962) );
  ANDN U24172 ( .B(n14596), .A(n14597), .Z(n14594) );
  AND U24173 ( .A(a[36]), .B(b[70]), .Z(n14593) );
  XNOR U24174 ( .A(n14598), .B(n13967), .Z(n13969) );
  XOR U24175 ( .A(n14599), .B(n14600), .Z(n13967) );
  ANDN U24176 ( .B(n14601), .A(n14602), .Z(n14599) );
  AND U24177 ( .A(a[37]), .B(b[69]), .Z(n14598) );
  XNOR U24178 ( .A(n14603), .B(n13972), .Z(n13974) );
  XOR U24179 ( .A(n14604), .B(n14605), .Z(n13972) );
  ANDN U24180 ( .B(n14606), .A(n14607), .Z(n14604) );
  AND U24181 ( .A(a[38]), .B(b[68]), .Z(n14603) );
  XNOR U24182 ( .A(n14608), .B(n13977), .Z(n13979) );
  XOR U24183 ( .A(n14609), .B(n14610), .Z(n13977) );
  ANDN U24184 ( .B(n14611), .A(n14612), .Z(n14609) );
  AND U24185 ( .A(a[39]), .B(b[67]), .Z(n14608) );
  XNOR U24186 ( .A(n14613), .B(n13982), .Z(n13984) );
  XOR U24187 ( .A(n14614), .B(n14615), .Z(n13982) );
  ANDN U24188 ( .B(n14616), .A(n14617), .Z(n14614) );
  AND U24189 ( .A(a[40]), .B(b[66]), .Z(n14613) );
  XNOR U24190 ( .A(n14618), .B(n13987), .Z(n13989) );
  XOR U24191 ( .A(n14619), .B(n14620), .Z(n13987) );
  ANDN U24192 ( .B(n14621), .A(n14622), .Z(n14619) );
  AND U24193 ( .A(a[41]), .B(b[65]), .Z(n14618) );
  XNOR U24194 ( .A(n14623), .B(n13992), .Z(n13994) );
  XOR U24195 ( .A(n14624), .B(n14625), .Z(n13992) );
  ANDN U24196 ( .B(n14626), .A(n14627), .Z(n14624) );
  AND U24197 ( .A(a[42]), .B(b[64]), .Z(n14623) );
  XNOR U24198 ( .A(n14628), .B(n13997), .Z(n13999) );
  XOR U24199 ( .A(n14629), .B(n14630), .Z(n13997) );
  ANDN U24200 ( .B(n14631), .A(n14632), .Z(n14629) );
  AND U24201 ( .A(a[43]), .B(b[63]), .Z(n14628) );
  XNOR U24202 ( .A(n14633), .B(n14002), .Z(n14004) );
  XOR U24203 ( .A(n14634), .B(n14635), .Z(n14002) );
  ANDN U24204 ( .B(n14636), .A(n14637), .Z(n14634) );
  AND U24205 ( .A(a[44]), .B(b[62]), .Z(n14633) );
  XNOR U24206 ( .A(n14638), .B(n14007), .Z(n14009) );
  XOR U24207 ( .A(n14639), .B(n14640), .Z(n14007) );
  ANDN U24208 ( .B(n14641), .A(n14642), .Z(n14639) );
  AND U24209 ( .A(a[45]), .B(b[61]), .Z(n14638) );
  XNOR U24210 ( .A(n14643), .B(n14012), .Z(n14014) );
  XOR U24211 ( .A(n14644), .B(n14645), .Z(n14012) );
  ANDN U24212 ( .B(n14646), .A(n14647), .Z(n14644) );
  AND U24213 ( .A(a[46]), .B(b[60]), .Z(n14643) );
  XNOR U24214 ( .A(n14648), .B(n14017), .Z(n14019) );
  XOR U24215 ( .A(n14649), .B(n14650), .Z(n14017) );
  ANDN U24216 ( .B(n14651), .A(n14652), .Z(n14649) );
  AND U24217 ( .A(a[47]), .B(b[59]), .Z(n14648) );
  XNOR U24218 ( .A(n14653), .B(n14022), .Z(n14024) );
  XOR U24219 ( .A(n14654), .B(n14655), .Z(n14022) );
  ANDN U24220 ( .B(n14656), .A(n14657), .Z(n14654) );
  AND U24221 ( .A(a[48]), .B(b[58]), .Z(n14653) );
  XNOR U24222 ( .A(n14658), .B(n14027), .Z(n14029) );
  XOR U24223 ( .A(n14659), .B(n14660), .Z(n14027) );
  ANDN U24224 ( .B(n14661), .A(n14662), .Z(n14659) );
  AND U24225 ( .A(a[49]), .B(b[57]), .Z(n14658) );
  XNOR U24226 ( .A(n14663), .B(n14032), .Z(n14034) );
  XOR U24227 ( .A(n14664), .B(n14665), .Z(n14032) );
  ANDN U24228 ( .B(n14666), .A(n14667), .Z(n14664) );
  AND U24229 ( .A(a[50]), .B(b[56]), .Z(n14663) );
  XNOR U24230 ( .A(n14668), .B(n14037), .Z(n14039) );
  XOR U24231 ( .A(n14669), .B(n14670), .Z(n14037) );
  ANDN U24232 ( .B(n14671), .A(n14672), .Z(n14669) );
  AND U24233 ( .A(a[51]), .B(b[55]), .Z(n14668) );
  XNOR U24234 ( .A(n14673), .B(n14042), .Z(n14044) );
  XOR U24235 ( .A(n14674), .B(n14675), .Z(n14042) );
  ANDN U24236 ( .B(n14676), .A(n14677), .Z(n14674) );
  AND U24237 ( .A(a[52]), .B(b[54]), .Z(n14673) );
  XNOR U24238 ( .A(n14678), .B(n14047), .Z(n14049) );
  XOR U24239 ( .A(n14679), .B(n14680), .Z(n14047) );
  ANDN U24240 ( .B(n14681), .A(n14682), .Z(n14679) );
  AND U24241 ( .A(a[53]), .B(b[53]), .Z(n14678) );
  XNOR U24242 ( .A(n14683), .B(n14052), .Z(n14054) );
  XOR U24243 ( .A(n14684), .B(n14685), .Z(n14052) );
  ANDN U24244 ( .B(n14686), .A(n14687), .Z(n14684) );
  AND U24245 ( .A(a[54]), .B(b[52]), .Z(n14683) );
  XNOR U24246 ( .A(n14688), .B(n14057), .Z(n14059) );
  XOR U24247 ( .A(n14689), .B(n14690), .Z(n14057) );
  ANDN U24248 ( .B(n14691), .A(n14692), .Z(n14689) );
  AND U24249 ( .A(a[55]), .B(b[51]), .Z(n14688) );
  XNOR U24250 ( .A(n14693), .B(n14062), .Z(n14064) );
  XOR U24251 ( .A(n14694), .B(n14695), .Z(n14062) );
  ANDN U24252 ( .B(n14696), .A(n14697), .Z(n14694) );
  AND U24253 ( .A(a[56]), .B(b[50]), .Z(n14693) );
  XNOR U24254 ( .A(n14698), .B(n14067), .Z(n14069) );
  XOR U24255 ( .A(n14699), .B(n14700), .Z(n14067) );
  ANDN U24256 ( .B(n14701), .A(n14702), .Z(n14699) );
  AND U24257 ( .A(a[57]), .B(b[49]), .Z(n14698) );
  XNOR U24258 ( .A(n14703), .B(n14072), .Z(n14074) );
  XOR U24259 ( .A(n14704), .B(n14705), .Z(n14072) );
  ANDN U24260 ( .B(n14706), .A(n14707), .Z(n14704) );
  AND U24261 ( .A(a[58]), .B(b[48]), .Z(n14703) );
  XNOR U24262 ( .A(n14708), .B(n14077), .Z(n14079) );
  XOR U24263 ( .A(n14709), .B(n14710), .Z(n14077) );
  ANDN U24264 ( .B(n14711), .A(n14712), .Z(n14709) );
  AND U24265 ( .A(a[59]), .B(b[47]), .Z(n14708) );
  XNOR U24266 ( .A(n14713), .B(n14082), .Z(n14084) );
  XOR U24267 ( .A(n14714), .B(n14715), .Z(n14082) );
  ANDN U24268 ( .B(n14716), .A(n14717), .Z(n14714) );
  AND U24269 ( .A(a[60]), .B(b[46]), .Z(n14713) );
  XNOR U24270 ( .A(n14718), .B(n14087), .Z(n14089) );
  XOR U24271 ( .A(n14719), .B(n14720), .Z(n14087) );
  ANDN U24272 ( .B(n14721), .A(n14722), .Z(n14719) );
  AND U24273 ( .A(a[61]), .B(b[45]), .Z(n14718) );
  XNOR U24274 ( .A(n14723), .B(n14092), .Z(n14094) );
  XOR U24275 ( .A(n14724), .B(n14725), .Z(n14092) );
  ANDN U24276 ( .B(n14726), .A(n14727), .Z(n14724) );
  AND U24277 ( .A(a[62]), .B(b[44]), .Z(n14723) );
  XNOR U24278 ( .A(n14728), .B(n14097), .Z(n14099) );
  XOR U24279 ( .A(n14729), .B(n14730), .Z(n14097) );
  ANDN U24280 ( .B(n14731), .A(n14732), .Z(n14729) );
  AND U24281 ( .A(a[63]), .B(b[43]), .Z(n14728) );
  XNOR U24282 ( .A(n14733), .B(n14102), .Z(n14104) );
  XOR U24283 ( .A(n14734), .B(n14735), .Z(n14102) );
  ANDN U24284 ( .B(n14736), .A(n14737), .Z(n14734) );
  AND U24285 ( .A(a[64]), .B(b[42]), .Z(n14733) );
  XNOR U24286 ( .A(n14738), .B(n14107), .Z(n14109) );
  XOR U24287 ( .A(n14739), .B(n14740), .Z(n14107) );
  ANDN U24288 ( .B(n14741), .A(n14742), .Z(n14739) );
  AND U24289 ( .A(a[65]), .B(b[41]), .Z(n14738) );
  XNOR U24290 ( .A(n14743), .B(n14112), .Z(n14114) );
  XOR U24291 ( .A(n14744), .B(n14745), .Z(n14112) );
  ANDN U24292 ( .B(n14746), .A(n14747), .Z(n14744) );
  AND U24293 ( .A(a[66]), .B(b[40]), .Z(n14743) );
  XNOR U24294 ( .A(n14748), .B(n14117), .Z(n14119) );
  XOR U24295 ( .A(n14749), .B(n14750), .Z(n14117) );
  ANDN U24296 ( .B(n14751), .A(n14752), .Z(n14749) );
  AND U24297 ( .A(a[67]), .B(b[39]), .Z(n14748) );
  XNOR U24298 ( .A(n14753), .B(n14122), .Z(n14124) );
  XOR U24299 ( .A(n14754), .B(n14755), .Z(n14122) );
  ANDN U24300 ( .B(n14756), .A(n14757), .Z(n14754) );
  AND U24301 ( .A(a[68]), .B(b[38]), .Z(n14753) );
  XNOR U24302 ( .A(n14758), .B(n14127), .Z(n14129) );
  XOR U24303 ( .A(n14759), .B(n14760), .Z(n14127) );
  ANDN U24304 ( .B(n14761), .A(n14762), .Z(n14759) );
  AND U24305 ( .A(a[69]), .B(b[37]), .Z(n14758) );
  XNOR U24306 ( .A(n14763), .B(n14132), .Z(n14134) );
  XOR U24307 ( .A(n14764), .B(n14765), .Z(n14132) );
  ANDN U24308 ( .B(n14766), .A(n14767), .Z(n14764) );
  AND U24309 ( .A(a[70]), .B(b[36]), .Z(n14763) );
  XNOR U24310 ( .A(n14768), .B(n14137), .Z(n14139) );
  XOR U24311 ( .A(n14769), .B(n14770), .Z(n14137) );
  ANDN U24312 ( .B(n14771), .A(n14772), .Z(n14769) );
  AND U24313 ( .A(a[71]), .B(b[35]), .Z(n14768) );
  XNOR U24314 ( .A(n14773), .B(n14142), .Z(n14144) );
  XOR U24315 ( .A(n14774), .B(n14775), .Z(n14142) );
  ANDN U24316 ( .B(n14776), .A(n14777), .Z(n14774) );
  AND U24317 ( .A(a[72]), .B(b[34]), .Z(n14773) );
  XNOR U24318 ( .A(n14778), .B(n14147), .Z(n14149) );
  XOR U24319 ( .A(n14779), .B(n14780), .Z(n14147) );
  ANDN U24320 ( .B(n14781), .A(n14782), .Z(n14779) );
  AND U24321 ( .A(a[73]), .B(b[33]), .Z(n14778) );
  XNOR U24322 ( .A(n14783), .B(n14152), .Z(n14154) );
  XOR U24323 ( .A(n14784), .B(n14785), .Z(n14152) );
  ANDN U24324 ( .B(n14786), .A(n14787), .Z(n14784) );
  AND U24325 ( .A(a[74]), .B(b[32]), .Z(n14783) );
  XNOR U24326 ( .A(n14788), .B(n14157), .Z(n14159) );
  XOR U24327 ( .A(n14789), .B(n14790), .Z(n14157) );
  ANDN U24328 ( .B(n14791), .A(n14792), .Z(n14789) );
  AND U24329 ( .A(a[75]), .B(b[31]), .Z(n14788) );
  XNOR U24330 ( .A(n14793), .B(n14162), .Z(n14164) );
  XOR U24331 ( .A(n14794), .B(n14795), .Z(n14162) );
  ANDN U24332 ( .B(n14796), .A(n14797), .Z(n14794) );
  AND U24333 ( .A(a[76]), .B(b[30]), .Z(n14793) );
  XNOR U24334 ( .A(n14798), .B(n14167), .Z(n14169) );
  XOR U24335 ( .A(n14799), .B(n14800), .Z(n14167) );
  ANDN U24336 ( .B(n14801), .A(n14802), .Z(n14799) );
  AND U24337 ( .A(a[77]), .B(b[29]), .Z(n14798) );
  XNOR U24338 ( .A(n14803), .B(n14172), .Z(n14174) );
  XOR U24339 ( .A(n14804), .B(n14805), .Z(n14172) );
  ANDN U24340 ( .B(n14806), .A(n14807), .Z(n14804) );
  AND U24341 ( .A(a[78]), .B(b[28]), .Z(n14803) );
  XNOR U24342 ( .A(n14808), .B(n14177), .Z(n14179) );
  XOR U24343 ( .A(n14809), .B(n14810), .Z(n14177) );
  ANDN U24344 ( .B(n14811), .A(n14812), .Z(n14809) );
  AND U24345 ( .A(a[79]), .B(b[27]), .Z(n14808) );
  XNOR U24346 ( .A(n14813), .B(n14182), .Z(n14184) );
  XOR U24347 ( .A(n14814), .B(n14815), .Z(n14182) );
  ANDN U24348 ( .B(n14816), .A(n14817), .Z(n14814) );
  AND U24349 ( .A(a[80]), .B(b[26]), .Z(n14813) );
  XNOR U24350 ( .A(n14818), .B(n14187), .Z(n14189) );
  XOR U24351 ( .A(n14819), .B(n14820), .Z(n14187) );
  ANDN U24352 ( .B(n14821), .A(n14822), .Z(n14819) );
  AND U24353 ( .A(a[81]), .B(b[25]), .Z(n14818) );
  XNOR U24354 ( .A(n14823), .B(n14192), .Z(n14194) );
  XOR U24355 ( .A(n14824), .B(n14825), .Z(n14192) );
  ANDN U24356 ( .B(n14826), .A(n14827), .Z(n14824) );
  AND U24357 ( .A(a[82]), .B(b[24]), .Z(n14823) );
  XNOR U24358 ( .A(n14828), .B(n14197), .Z(n14199) );
  XOR U24359 ( .A(n14829), .B(n14830), .Z(n14197) );
  ANDN U24360 ( .B(n14831), .A(n14832), .Z(n14829) );
  AND U24361 ( .A(a[83]), .B(b[23]), .Z(n14828) );
  XNOR U24362 ( .A(n14833), .B(n14202), .Z(n14204) );
  XOR U24363 ( .A(n14834), .B(n14835), .Z(n14202) );
  ANDN U24364 ( .B(n14836), .A(n14837), .Z(n14834) );
  AND U24365 ( .A(a[84]), .B(b[22]), .Z(n14833) );
  XNOR U24366 ( .A(n14838), .B(n14207), .Z(n14209) );
  XOR U24367 ( .A(n14839), .B(n14840), .Z(n14207) );
  ANDN U24368 ( .B(n14841), .A(n14842), .Z(n14839) );
  AND U24369 ( .A(a[85]), .B(b[21]), .Z(n14838) );
  XNOR U24370 ( .A(n14843), .B(n14212), .Z(n14214) );
  XOR U24371 ( .A(n14844), .B(n14845), .Z(n14212) );
  ANDN U24372 ( .B(n14846), .A(n14847), .Z(n14844) );
  AND U24373 ( .A(a[86]), .B(b[20]), .Z(n14843) );
  XNOR U24374 ( .A(n14848), .B(n14217), .Z(n14219) );
  XOR U24375 ( .A(n14849), .B(n14850), .Z(n14217) );
  ANDN U24376 ( .B(n14851), .A(n14852), .Z(n14849) );
  AND U24377 ( .A(a[87]), .B(b[19]), .Z(n14848) );
  XNOR U24378 ( .A(n14853), .B(n14222), .Z(n14224) );
  XOR U24379 ( .A(n14854), .B(n14855), .Z(n14222) );
  ANDN U24380 ( .B(n14856), .A(n14857), .Z(n14854) );
  AND U24381 ( .A(a[88]), .B(b[18]), .Z(n14853) );
  XNOR U24382 ( .A(n14858), .B(n14227), .Z(n14229) );
  XOR U24383 ( .A(n14859), .B(n14860), .Z(n14227) );
  ANDN U24384 ( .B(n14861), .A(n14862), .Z(n14859) );
  AND U24385 ( .A(a[89]), .B(b[17]), .Z(n14858) );
  XNOR U24386 ( .A(n14863), .B(n14232), .Z(n14234) );
  XOR U24387 ( .A(n14864), .B(n14865), .Z(n14232) );
  ANDN U24388 ( .B(n14866), .A(n14867), .Z(n14864) );
  AND U24389 ( .A(a[90]), .B(b[16]), .Z(n14863) );
  XNOR U24390 ( .A(n14868), .B(n14237), .Z(n14239) );
  XOR U24391 ( .A(n14869), .B(n14870), .Z(n14237) );
  ANDN U24392 ( .B(n14871), .A(n14872), .Z(n14869) );
  AND U24393 ( .A(a[91]), .B(b[15]), .Z(n14868) );
  XNOR U24394 ( .A(n14873), .B(n14242), .Z(n14244) );
  XOR U24395 ( .A(n14874), .B(n14875), .Z(n14242) );
  ANDN U24396 ( .B(n14876), .A(n14877), .Z(n14874) );
  AND U24397 ( .A(a[92]), .B(b[14]), .Z(n14873) );
  XNOR U24398 ( .A(n14878), .B(n14247), .Z(n14249) );
  XOR U24399 ( .A(n14879), .B(n14880), .Z(n14247) );
  ANDN U24400 ( .B(n14881), .A(n14882), .Z(n14879) );
  AND U24401 ( .A(a[93]), .B(b[13]), .Z(n14878) );
  XNOR U24402 ( .A(n14883), .B(n14252), .Z(n14254) );
  XOR U24403 ( .A(n14884), .B(n14885), .Z(n14252) );
  ANDN U24404 ( .B(n14886), .A(n14887), .Z(n14884) );
  AND U24405 ( .A(a[94]), .B(b[12]), .Z(n14883) );
  XNOR U24406 ( .A(n14888), .B(n14257), .Z(n14259) );
  XOR U24407 ( .A(n14889), .B(n14890), .Z(n14257) );
  ANDN U24408 ( .B(n14891), .A(n14892), .Z(n14889) );
  AND U24409 ( .A(a[95]), .B(b[11]), .Z(n14888) );
  XNOR U24410 ( .A(n14893), .B(n14262), .Z(n14264) );
  XOR U24411 ( .A(n14894), .B(n14895), .Z(n14262) );
  ANDN U24412 ( .B(n14896), .A(n14897), .Z(n14894) );
  AND U24413 ( .A(a[96]), .B(b[10]), .Z(n14893) );
  XNOR U24414 ( .A(n14898), .B(n14267), .Z(n14269) );
  XOR U24415 ( .A(n14899), .B(n14900), .Z(n14267) );
  ANDN U24416 ( .B(n14901), .A(n14902), .Z(n14899) );
  AND U24417 ( .A(b[9]), .B(a[97]), .Z(n14898) );
  XNOR U24418 ( .A(n14903), .B(n14272), .Z(n14274) );
  XOR U24419 ( .A(n14904), .B(n14905), .Z(n14272) );
  ANDN U24420 ( .B(n14906), .A(n14907), .Z(n14904) );
  AND U24421 ( .A(b[8]), .B(a[98]), .Z(n14903) );
  XNOR U24422 ( .A(n14908), .B(n14277), .Z(n14279) );
  XOR U24423 ( .A(n14909), .B(n14910), .Z(n14277) );
  ANDN U24424 ( .B(n14911), .A(n14912), .Z(n14909) );
  AND U24425 ( .A(b[7]), .B(a[99]), .Z(n14908) );
  XNOR U24426 ( .A(n14913), .B(n14282), .Z(n14284) );
  XOR U24427 ( .A(n14914), .B(n14915), .Z(n14282) );
  ANDN U24428 ( .B(n14916), .A(n14917), .Z(n14914) );
  AND U24429 ( .A(b[6]), .B(a[100]), .Z(n14913) );
  XNOR U24430 ( .A(n14918), .B(n14287), .Z(n14289) );
  XOR U24431 ( .A(n14919), .B(n14920), .Z(n14287) );
  ANDN U24432 ( .B(n14921), .A(n14922), .Z(n14919) );
  AND U24433 ( .A(b[5]), .B(a[101]), .Z(n14918) );
  XNOR U24434 ( .A(n14923), .B(n14292), .Z(n14294) );
  XOR U24435 ( .A(n14924), .B(n14925), .Z(n14292) );
  ANDN U24436 ( .B(n14926), .A(n14927), .Z(n14924) );
  AND U24437 ( .A(b[4]), .B(a[102]), .Z(n14923) );
  XNOR U24438 ( .A(n14928), .B(n14929), .Z(n14306) );
  NANDN U24439 ( .A(n14930), .B(n14931), .Z(n14929) );
  XNOR U24440 ( .A(n14932), .B(n14297), .Z(n14299) );
  XNOR U24441 ( .A(n14933), .B(n14934), .Z(n14297) );
  AND U24442 ( .A(n14935), .B(n14936), .Z(n14933) );
  AND U24443 ( .A(b[3]), .B(a[103]), .Z(n14932) );
  NAND U24444 ( .A(a[106]), .B(b[0]), .Z(n13678) );
  XNOR U24445 ( .A(n14312), .B(n14313), .Z(c[105]) );
  XNOR U24446 ( .A(n14930), .B(n14931), .Z(n14313) );
  XOR U24447 ( .A(n14928), .B(n14937), .Z(n14931) );
  NAND U24448 ( .A(b[1]), .B(a[104]), .Z(n14937) );
  XOR U24449 ( .A(n14936), .B(n14938), .Z(n14930) );
  XOR U24450 ( .A(n14928), .B(n14935), .Z(n14938) );
  XNOR U24451 ( .A(n14939), .B(n14934), .Z(n14935) );
  AND U24452 ( .A(b[2]), .B(a[103]), .Z(n14939) );
  NANDN U24453 ( .A(n14940), .B(n14941), .Z(n14928) );
  XOR U24454 ( .A(n14934), .B(n14926), .Z(n14942) );
  XNOR U24455 ( .A(n14925), .B(n14921), .Z(n14943) );
  XNOR U24456 ( .A(n14920), .B(n14916), .Z(n14944) );
  XNOR U24457 ( .A(n14915), .B(n14911), .Z(n14945) );
  XNOR U24458 ( .A(n14910), .B(n14906), .Z(n14946) );
  XNOR U24459 ( .A(n14905), .B(n14901), .Z(n14947) );
  XNOR U24460 ( .A(n14900), .B(n14896), .Z(n14948) );
  XNOR U24461 ( .A(n14895), .B(n14891), .Z(n14949) );
  XNOR U24462 ( .A(n14890), .B(n14886), .Z(n14950) );
  XNOR U24463 ( .A(n14885), .B(n14881), .Z(n14951) );
  XNOR U24464 ( .A(n14880), .B(n14876), .Z(n14952) );
  XNOR U24465 ( .A(n14875), .B(n14871), .Z(n14953) );
  XNOR U24466 ( .A(n14870), .B(n14866), .Z(n14954) );
  XNOR U24467 ( .A(n14865), .B(n14861), .Z(n14955) );
  XNOR U24468 ( .A(n14860), .B(n14856), .Z(n14956) );
  XNOR U24469 ( .A(n14855), .B(n14851), .Z(n14957) );
  XNOR U24470 ( .A(n14850), .B(n14846), .Z(n14958) );
  XNOR U24471 ( .A(n14845), .B(n14841), .Z(n14959) );
  XNOR U24472 ( .A(n14840), .B(n14836), .Z(n14960) );
  XNOR U24473 ( .A(n14835), .B(n14831), .Z(n14961) );
  XNOR U24474 ( .A(n14830), .B(n14826), .Z(n14962) );
  XNOR U24475 ( .A(n14825), .B(n14821), .Z(n14963) );
  XNOR U24476 ( .A(n14820), .B(n14816), .Z(n14964) );
  XNOR U24477 ( .A(n14815), .B(n14811), .Z(n14965) );
  XNOR U24478 ( .A(n14810), .B(n14806), .Z(n14966) );
  XNOR U24479 ( .A(n14805), .B(n14801), .Z(n14967) );
  XNOR U24480 ( .A(n14800), .B(n14796), .Z(n14968) );
  XNOR U24481 ( .A(n14795), .B(n14791), .Z(n14969) );
  XNOR U24482 ( .A(n14790), .B(n14786), .Z(n14970) );
  XNOR U24483 ( .A(n14785), .B(n14781), .Z(n14971) );
  XNOR U24484 ( .A(n14780), .B(n14776), .Z(n14972) );
  XNOR U24485 ( .A(n14775), .B(n14771), .Z(n14973) );
  XNOR U24486 ( .A(n14770), .B(n14766), .Z(n14974) );
  XNOR U24487 ( .A(n14765), .B(n14761), .Z(n14975) );
  XNOR U24488 ( .A(n14760), .B(n14756), .Z(n14976) );
  XNOR U24489 ( .A(n14755), .B(n14751), .Z(n14977) );
  XNOR U24490 ( .A(n14750), .B(n14746), .Z(n14978) );
  XNOR U24491 ( .A(n14745), .B(n14741), .Z(n14979) );
  XNOR U24492 ( .A(n14740), .B(n14736), .Z(n14980) );
  XNOR U24493 ( .A(n14735), .B(n14731), .Z(n14981) );
  XNOR U24494 ( .A(n14730), .B(n14726), .Z(n14982) );
  XNOR U24495 ( .A(n14725), .B(n14721), .Z(n14983) );
  XNOR U24496 ( .A(n14720), .B(n14716), .Z(n14984) );
  XNOR U24497 ( .A(n14715), .B(n14711), .Z(n14985) );
  XNOR U24498 ( .A(n14710), .B(n14706), .Z(n14986) );
  XNOR U24499 ( .A(n14705), .B(n14701), .Z(n14987) );
  XNOR U24500 ( .A(n14700), .B(n14696), .Z(n14988) );
  XNOR U24501 ( .A(n14695), .B(n14691), .Z(n14989) );
  XNOR U24502 ( .A(n14690), .B(n14686), .Z(n14990) );
  XNOR U24503 ( .A(n14685), .B(n14681), .Z(n14991) );
  XNOR U24504 ( .A(n14680), .B(n14676), .Z(n14992) );
  XNOR U24505 ( .A(n14675), .B(n14671), .Z(n14993) );
  XNOR U24506 ( .A(n14670), .B(n14666), .Z(n14994) );
  XNOR U24507 ( .A(n14665), .B(n14661), .Z(n14995) );
  XNOR U24508 ( .A(n14660), .B(n14656), .Z(n14996) );
  XNOR U24509 ( .A(n14655), .B(n14651), .Z(n14997) );
  XNOR U24510 ( .A(n14650), .B(n14646), .Z(n14998) );
  XNOR U24511 ( .A(n14645), .B(n14641), .Z(n14999) );
  XNOR U24512 ( .A(n14640), .B(n14636), .Z(n15000) );
  XNOR U24513 ( .A(n14635), .B(n14631), .Z(n15001) );
  XNOR U24514 ( .A(n14630), .B(n14626), .Z(n15002) );
  XNOR U24515 ( .A(n14625), .B(n14621), .Z(n15003) );
  XNOR U24516 ( .A(n14620), .B(n14616), .Z(n15004) );
  XNOR U24517 ( .A(n14615), .B(n14611), .Z(n15005) );
  XNOR U24518 ( .A(n14610), .B(n14606), .Z(n15006) );
  XNOR U24519 ( .A(n14605), .B(n14601), .Z(n15007) );
  XNOR U24520 ( .A(n14600), .B(n14596), .Z(n15008) );
  XNOR U24521 ( .A(n14595), .B(n14591), .Z(n15009) );
  XNOR U24522 ( .A(n14590), .B(n14586), .Z(n15010) );
  XNOR U24523 ( .A(n14585), .B(n14581), .Z(n15011) );
  XNOR U24524 ( .A(n14580), .B(n14576), .Z(n15012) );
  XNOR U24525 ( .A(n14575), .B(n14571), .Z(n15013) );
  XNOR U24526 ( .A(n14570), .B(n14566), .Z(n15014) );
  XNOR U24527 ( .A(n14565), .B(n14561), .Z(n15015) );
  XNOR U24528 ( .A(n14560), .B(n14556), .Z(n15016) );
  XNOR U24529 ( .A(n14555), .B(n14551), .Z(n15017) );
  XNOR U24530 ( .A(n14550), .B(n14546), .Z(n15018) );
  XNOR U24531 ( .A(n14545), .B(n14541), .Z(n15019) );
  XNOR U24532 ( .A(n14540), .B(n14536), .Z(n15020) );
  XNOR U24533 ( .A(n14535), .B(n14531), .Z(n15021) );
  XNOR U24534 ( .A(n14530), .B(n14526), .Z(n15022) );
  XNOR U24535 ( .A(n14525), .B(n14521), .Z(n15023) );
  XNOR U24536 ( .A(n14520), .B(n14516), .Z(n15024) );
  XNOR U24537 ( .A(n14515), .B(n14511), .Z(n15025) );
  XNOR U24538 ( .A(n14510), .B(n14506), .Z(n15026) );
  XNOR U24539 ( .A(n14505), .B(n14501), .Z(n15027) );
  XNOR U24540 ( .A(n14500), .B(n14496), .Z(n15028) );
  XNOR U24541 ( .A(n14495), .B(n14491), .Z(n15029) );
  XNOR U24542 ( .A(n14490), .B(n14486), .Z(n15030) );
  XNOR U24543 ( .A(n14485), .B(n14481), .Z(n15031) );
  XNOR U24544 ( .A(n14480), .B(n14476), .Z(n15032) );
  XNOR U24545 ( .A(n14475), .B(n14471), .Z(n15033) );
  XNOR U24546 ( .A(n14470), .B(n14466), .Z(n15034) );
  XNOR U24547 ( .A(n14465), .B(n14461), .Z(n15035) );
  XNOR U24548 ( .A(n14460), .B(n14456), .Z(n15036) );
  XNOR U24549 ( .A(n14455), .B(n14451), .Z(n15037) );
  XNOR U24550 ( .A(n14450), .B(n14446), .Z(n15038) );
  XNOR U24551 ( .A(n14445), .B(n14441), .Z(n15039) );
  XNOR U24552 ( .A(n14440), .B(n14436), .Z(n15040) );
  XNOR U24553 ( .A(n14435), .B(n14431), .Z(n15041) );
  XNOR U24554 ( .A(n14430), .B(n14426), .Z(n15042) );
  XNOR U24555 ( .A(n14425), .B(n14421), .Z(n15043) );
  XNOR U24556 ( .A(n15044), .B(n14420), .Z(n14421) );
  AND U24557 ( .A(a[0]), .B(b[105]), .Z(n15044) );
  XOR U24558 ( .A(n15045), .B(n14420), .Z(n14422) );
  XNOR U24559 ( .A(n15046), .B(n15047), .Z(n14420) );
  ANDN U24560 ( .B(n15048), .A(n15049), .Z(n15046) );
  AND U24561 ( .A(a[1]), .B(b[104]), .Z(n15045) );
  XNOR U24562 ( .A(n15050), .B(n14425), .Z(n14427) );
  XOR U24563 ( .A(n15051), .B(n15052), .Z(n14425) );
  ANDN U24564 ( .B(n15053), .A(n15054), .Z(n15051) );
  AND U24565 ( .A(a[2]), .B(b[103]), .Z(n15050) );
  XNOR U24566 ( .A(n15055), .B(n14430), .Z(n14432) );
  XOR U24567 ( .A(n15056), .B(n15057), .Z(n14430) );
  ANDN U24568 ( .B(n15058), .A(n15059), .Z(n15056) );
  AND U24569 ( .A(a[3]), .B(b[102]), .Z(n15055) );
  XNOR U24570 ( .A(n15060), .B(n14435), .Z(n14437) );
  XOR U24571 ( .A(n15061), .B(n15062), .Z(n14435) );
  ANDN U24572 ( .B(n15063), .A(n15064), .Z(n15061) );
  AND U24573 ( .A(a[4]), .B(b[101]), .Z(n15060) );
  XNOR U24574 ( .A(n15065), .B(n14440), .Z(n14442) );
  XOR U24575 ( .A(n15066), .B(n15067), .Z(n14440) );
  ANDN U24576 ( .B(n15068), .A(n15069), .Z(n15066) );
  AND U24577 ( .A(a[5]), .B(b[100]), .Z(n15065) );
  XNOR U24578 ( .A(n15070), .B(n14445), .Z(n14447) );
  XOR U24579 ( .A(n15071), .B(n15072), .Z(n14445) );
  ANDN U24580 ( .B(n15073), .A(n15074), .Z(n15071) );
  AND U24581 ( .A(a[6]), .B(b[99]), .Z(n15070) );
  XNOR U24582 ( .A(n15075), .B(n14450), .Z(n14452) );
  XOR U24583 ( .A(n15076), .B(n15077), .Z(n14450) );
  ANDN U24584 ( .B(n15078), .A(n15079), .Z(n15076) );
  AND U24585 ( .A(a[7]), .B(b[98]), .Z(n15075) );
  XNOR U24586 ( .A(n15080), .B(n14455), .Z(n14457) );
  XOR U24587 ( .A(n15081), .B(n15082), .Z(n14455) );
  ANDN U24588 ( .B(n15083), .A(n15084), .Z(n15081) );
  AND U24589 ( .A(a[8]), .B(b[97]), .Z(n15080) );
  XNOR U24590 ( .A(n15085), .B(n14460), .Z(n14462) );
  XOR U24591 ( .A(n15086), .B(n15087), .Z(n14460) );
  ANDN U24592 ( .B(n15088), .A(n15089), .Z(n15086) );
  AND U24593 ( .A(a[9]), .B(b[96]), .Z(n15085) );
  XNOR U24594 ( .A(n15090), .B(n14465), .Z(n14467) );
  XOR U24595 ( .A(n15091), .B(n15092), .Z(n14465) );
  ANDN U24596 ( .B(n15093), .A(n15094), .Z(n15091) );
  AND U24597 ( .A(a[10]), .B(b[95]), .Z(n15090) );
  XNOR U24598 ( .A(n15095), .B(n14470), .Z(n14472) );
  XOR U24599 ( .A(n15096), .B(n15097), .Z(n14470) );
  ANDN U24600 ( .B(n15098), .A(n15099), .Z(n15096) );
  AND U24601 ( .A(a[11]), .B(b[94]), .Z(n15095) );
  XNOR U24602 ( .A(n15100), .B(n14475), .Z(n14477) );
  XOR U24603 ( .A(n15101), .B(n15102), .Z(n14475) );
  ANDN U24604 ( .B(n15103), .A(n15104), .Z(n15101) );
  AND U24605 ( .A(a[12]), .B(b[93]), .Z(n15100) );
  XNOR U24606 ( .A(n15105), .B(n14480), .Z(n14482) );
  XOR U24607 ( .A(n15106), .B(n15107), .Z(n14480) );
  ANDN U24608 ( .B(n15108), .A(n15109), .Z(n15106) );
  AND U24609 ( .A(a[13]), .B(b[92]), .Z(n15105) );
  XNOR U24610 ( .A(n15110), .B(n14485), .Z(n14487) );
  XOR U24611 ( .A(n15111), .B(n15112), .Z(n14485) );
  ANDN U24612 ( .B(n15113), .A(n15114), .Z(n15111) );
  AND U24613 ( .A(a[14]), .B(b[91]), .Z(n15110) );
  XNOR U24614 ( .A(n15115), .B(n14490), .Z(n14492) );
  XOR U24615 ( .A(n15116), .B(n15117), .Z(n14490) );
  ANDN U24616 ( .B(n15118), .A(n15119), .Z(n15116) );
  AND U24617 ( .A(a[15]), .B(b[90]), .Z(n15115) );
  XNOR U24618 ( .A(n15120), .B(n14495), .Z(n14497) );
  XOR U24619 ( .A(n15121), .B(n15122), .Z(n14495) );
  ANDN U24620 ( .B(n15123), .A(n15124), .Z(n15121) );
  AND U24621 ( .A(a[16]), .B(b[89]), .Z(n15120) );
  XNOR U24622 ( .A(n15125), .B(n14500), .Z(n14502) );
  XOR U24623 ( .A(n15126), .B(n15127), .Z(n14500) );
  ANDN U24624 ( .B(n15128), .A(n15129), .Z(n15126) );
  AND U24625 ( .A(a[17]), .B(b[88]), .Z(n15125) );
  XNOR U24626 ( .A(n15130), .B(n14505), .Z(n14507) );
  XOR U24627 ( .A(n15131), .B(n15132), .Z(n14505) );
  ANDN U24628 ( .B(n15133), .A(n15134), .Z(n15131) );
  AND U24629 ( .A(a[18]), .B(b[87]), .Z(n15130) );
  XNOR U24630 ( .A(n15135), .B(n14510), .Z(n14512) );
  XOR U24631 ( .A(n15136), .B(n15137), .Z(n14510) );
  ANDN U24632 ( .B(n15138), .A(n15139), .Z(n15136) );
  AND U24633 ( .A(a[19]), .B(b[86]), .Z(n15135) );
  XNOR U24634 ( .A(n15140), .B(n14515), .Z(n14517) );
  XOR U24635 ( .A(n15141), .B(n15142), .Z(n14515) );
  ANDN U24636 ( .B(n15143), .A(n15144), .Z(n15141) );
  AND U24637 ( .A(a[20]), .B(b[85]), .Z(n15140) );
  XNOR U24638 ( .A(n15145), .B(n14520), .Z(n14522) );
  XOR U24639 ( .A(n15146), .B(n15147), .Z(n14520) );
  ANDN U24640 ( .B(n15148), .A(n15149), .Z(n15146) );
  AND U24641 ( .A(a[21]), .B(b[84]), .Z(n15145) );
  XNOR U24642 ( .A(n15150), .B(n14525), .Z(n14527) );
  XOR U24643 ( .A(n15151), .B(n15152), .Z(n14525) );
  ANDN U24644 ( .B(n15153), .A(n15154), .Z(n15151) );
  AND U24645 ( .A(a[22]), .B(b[83]), .Z(n15150) );
  XNOR U24646 ( .A(n15155), .B(n14530), .Z(n14532) );
  XOR U24647 ( .A(n15156), .B(n15157), .Z(n14530) );
  ANDN U24648 ( .B(n15158), .A(n15159), .Z(n15156) );
  AND U24649 ( .A(a[23]), .B(b[82]), .Z(n15155) );
  XNOR U24650 ( .A(n15160), .B(n14535), .Z(n14537) );
  XOR U24651 ( .A(n15161), .B(n15162), .Z(n14535) );
  ANDN U24652 ( .B(n15163), .A(n15164), .Z(n15161) );
  AND U24653 ( .A(a[24]), .B(b[81]), .Z(n15160) );
  XNOR U24654 ( .A(n15165), .B(n14540), .Z(n14542) );
  XOR U24655 ( .A(n15166), .B(n15167), .Z(n14540) );
  ANDN U24656 ( .B(n15168), .A(n15169), .Z(n15166) );
  AND U24657 ( .A(a[25]), .B(b[80]), .Z(n15165) );
  XNOR U24658 ( .A(n15170), .B(n14545), .Z(n14547) );
  XOR U24659 ( .A(n15171), .B(n15172), .Z(n14545) );
  ANDN U24660 ( .B(n15173), .A(n15174), .Z(n15171) );
  AND U24661 ( .A(a[26]), .B(b[79]), .Z(n15170) );
  XNOR U24662 ( .A(n15175), .B(n14550), .Z(n14552) );
  XOR U24663 ( .A(n15176), .B(n15177), .Z(n14550) );
  ANDN U24664 ( .B(n15178), .A(n15179), .Z(n15176) );
  AND U24665 ( .A(a[27]), .B(b[78]), .Z(n15175) );
  XNOR U24666 ( .A(n15180), .B(n14555), .Z(n14557) );
  XOR U24667 ( .A(n15181), .B(n15182), .Z(n14555) );
  ANDN U24668 ( .B(n15183), .A(n15184), .Z(n15181) );
  AND U24669 ( .A(a[28]), .B(b[77]), .Z(n15180) );
  XNOR U24670 ( .A(n15185), .B(n14560), .Z(n14562) );
  XOR U24671 ( .A(n15186), .B(n15187), .Z(n14560) );
  ANDN U24672 ( .B(n15188), .A(n15189), .Z(n15186) );
  AND U24673 ( .A(a[29]), .B(b[76]), .Z(n15185) );
  XNOR U24674 ( .A(n15190), .B(n14565), .Z(n14567) );
  XOR U24675 ( .A(n15191), .B(n15192), .Z(n14565) );
  ANDN U24676 ( .B(n15193), .A(n15194), .Z(n15191) );
  AND U24677 ( .A(a[30]), .B(b[75]), .Z(n15190) );
  XNOR U24678 ( .A(n15195), .B(n14570), .Z(n14572) );
  XOR U24679 ( .A(n15196), .B(n15197), .Z(n14570) );
  ANDN U24680 ( .B(n15198), .A(n15199), .Z(n15196) );
  AND U24681 ( .A(a[31]), .B(b[74]), .Z(n15195) );
  XNOR U24682 ( .A(n15200), .B(n14575), .Z(n14577) );
  XOR U24683 ( .A(n15201), .B(n15202), .Z(n14575) );
  ANDN U24684 ( .B(n15203), .A(n15204), .Z(n15201) );
  AND U24685 ( .A(a[32]), .B(b[73]), .Z(n15200) );
  XNOR U24686 ( .A(n15205), .B(n14580), .Z(n14582) );
  XOR U24687 ( .A(n15206), .B(n15207), .Z(n14580) );
  ANDN U24688 ( .B(n15208), .A(n15209), .Z(n15206) );
  AND U24689 ( .A(a[33]), .B(b[72]), .Z(n15205) );
  XNOR U24690 ( .A(n15210), .B(n14585), .Z(n14587) );
  XOR U24691 ( .A(n15211), .B(n15212), .Z(n14585) );
  ANDN U24692 ( .B(n15213), .A(n15214), .Z(n15211) );
  AND U24693 ( .A(a[34]), .B(b[71]), .Z(n15210) );
  XNOR U24694 ( .A(n15215), .B(n14590), .Z(n14592) );
  XOR U24695 ( .A(n15216), .B(n15217), .Z(n14590) );
  ANDN U24696 ( .B(n15218), .A(n15219), .Z(n15216) );
  AND U24697 ( .A(a[35]), .B(b[70]), .Z(n15215) );
  XNOR U24698 ( .A(n15220), .B(n14595), .Z(n14597) );
  XOR U24699 ( .A(n15221), .B(n15222), .Z(n14595) );
  ANDN U24700 ( .B(n15223), .A(n15224), .Z(n15221) );
  AND U24701 ( .A(a[36]), .B(b[69]), .Z(n15220) );
  XNOR U24702 ( .A(n15225), .B(n14600), .Z(n14602) );
  XOR U24703 ( .A(n15226), .B(n15227), .Z(n14600) );
  ANDN U24704 ( .B(n15228), .A(n15229), .Z(n15226) );
  AND U24705 ( .A(a[37]), .B(b[68]), .Z(n15225) );
  XNOR U24706 ( .A(n15230), .B(n14605), .Z(n14607) );
  XOR U24707 ( .A(n15231), .B(n15232), .Z(n14605) );
  ANDN U24708 ( .B(n15233), .A(n15234), .Z(n15231) );
  AND U24709 ( .A(a[38]), .B(b[67]), .Z(n15230) );
  XNOR U24710 ( .A(n15235), .B(n14610), .Z(n14612) );
  XOR U24711 ( .A(n15236), .B(n15237), .Z(n14610) );
  ANDN U24712 ( .B(n15238), .A(n15239), .Z(n15236) );
  AND U24713 ( .A(a[39]), .B(b[66]), .Z(n15235) );
  XNOR U24714 ( .A(n15240), .B(n14615), .Z(n14617) );
  XOR U24715 ( .A(n15241), .B(n15242), .Z(n14615) );
  ANDN U24716 ( .B(n15243), .A(n15244), .Z(n15241) );
  AND U24717 ( .A(a[40]), .B(b[65]), .Z(n15240) );
  XNOR U24718 ( .A(n15245), .B(n14620), .Z(n14622) );
  XOR U24719 ( .A(n15246), .B(n15247), .Z(n14620) );
  ANDN U24720 ( .B(n15248), .A(n15249), .Z(n15246) );
  AND U24721 ( .A(a[41]), .B(b[64]), .Z(n15245) );
  XNOR U24722 ( .A(n15250), .B(n14625), .Z(n14627) );
  XOR U24723 ( .A(n15251), .B(n15252), .Z(n14625) );
  ANDN U24724 ( .B(n15253), .A(n15254), .Z(n15251) );
  AND U24725 ( .A(a[42]), .B(b[63]), .Z(n15250) );
  XNOR U24726 ( .A(n15255), .B(n14630), .Z(n14632) );
  XOR U24727 ( .A(n15256), .B(n15257), .Z(n14630) );
  ANDN U24728 ( .B(n15258), .A(n15259), .Z(n15256) );
  AND U24729 ( .A(a[43]), .B(b[62]), .Z(n15255) );
  XNOR U24730 ( .A(n15260), .B(n14635), .Z(n14637) );
  XOR U24731 ( .A(n15261), .B(n15262), .Z(n14635) );
  ANDN U24732 ( .B(n15263), .A(n15264), .Z(n15261) );
  AND U24733 ( .A(a[44]), .B(b[61]), .Z(n15260) );
  XNOR U24734 ( .A(n15265), .B(n14640), .Z(n14642) );
  XOR U24735 ( .A(n15266), .B(n15267), .Z(n14640) );
  ANDN U24736 ( .B(n15268), .A(n15269), .Z(n15266) );
  AND U24737 ( .A(a[45]), .B(b[60]), .Z(n15265) );
  XNOR U24738 ( .A(n15270), .B(n14645), .Z(n14647) );
  XOR U24739 ( .A(n15271), .B(n15272), .Z(n14645) );
  ANDN U24740 ( .B(n15273), .A(n15274), .Z(n15271) );
  AND U24741 ( .A(a[46]), .B(b[59]), .Z(n15270) );
  XNOR U24742 ( .A(n15275), .B(n14650), .Z(n14652) );
  XOR U24743 ( .A(n15276), .B(n15277), .Z(n14650) );
  ANDN U24744 ( .B(n15278), .A(n15279), .Z(n15276) );
  AND U24745 ( .A(a[47]), .B(b[58]), .Z(n15275) );
  XNOR U24746 ( .A(n15280), .B(n14655), .Z(n14657) );
  XOR U24747 ( .A(n15281), .B(n15282), .Z(n14655) );
  ANDN U24748 ( .B(n15283), .A(n15284), .Z(n15281) );
  AND U24749 ( .A(a[48]), .B(b[57]), .Z(n15280) );
  XNOR U24750 ( .A(n15285), .B(n14660), .Z(n14662) );
  XOR U24751 ( .A(n15286), .B(n15287), .Z(n14660) );
  ANDN U24752 ( .B(n15288), .A(n15289), .Z(n15286) );
  AND U24753 ( .A(a[49]), .B(b[56]), .Z(n15285) );
  XNOR U24754 ( .A(n15290), .B(n14665), .Z(n14667) );
  XOR U24755 ( .A(n15291), .B(n15292), .Z(n14665) );
  ANDN U24756 ( .B(n15293), .A(n15294), .Z(n15291) );
  AND U24757 ( .A(a[50]), .B(b[55]), .Z(n15290) );
  XNOR U24758 ( .A(n15295), .B(n14670), .Z(n14672) );
  XOR U24759 ( .A(n15296), .B(n15297), .Z(n14670) );
  ANDN U24760 ( .B(n15298), .A(n15299), .Z(n15296) );
  AND U24761 ( .A(a[51]), .B(b[54]), .Z(n15295) );
  XNOR U24762 ( .A(n15300), .B(n14675), .Z(n14677) );
  XOR U24763 ( .A(n15301), .B(n15302), .Z(n14675) );
  ANDN U24764 ( .B(n15303), .A(n15304), .Z(n15301) );
  AND U24765 ( .A(a[52]), .B(b[53]), .Z(n15300) );
  XNOR U24766 ( .A(n15305), .B(n14680), .Z(n14682) );
  XOR U24767 ( .A(n15306), .B(n15307), .Z(n14680) );
  ANDN U24768 ( .B(n15308), .A(n15309), .Z(n15306) );
  AND U24769 ( .A(a[53]), .B(b[52]), .Z(n15305) );
  XNOR U24770 ( .A(n15310), .B(n14685), .Z(n14687) );
  XOR U24771 ( .A(n15311), .B(n15312), .Z(n14685) );
  ANDN U24772 ( .B(n15313), .A(n15314), .Z(n15311) );
  AND U24773 ( .A(a[54]), .B(b[51]), .Z(n15310) );
  XNOR U24774 ( .A(n15315), .B(n14690), .Z(n14692) );
  XOR U24775 ( .A(n15316), .B(n15317), .Z(n14690) );
  ANDN U24776 ( .B(n15318), .A(n15319), .Z(n15316) );
  AND U24777 ( .A(a[55]), .B(b[50]), .Z(n15315) );
  XNOR U24778 ( .A(n15320), .B(n14695), .Z(n14697) );
  XOR U24779 ( .A(n15321), .B(n15322), .Z(n14695) );
  ANDN U24780 ( .B(n15323), .A(n15324), .Z(n15321) );
  AND U24781 ( .A(a[56]), .B(b[49]), .Z(n15320) );
  XNOR U24782 ( .A(n15325), .B(n14700), .Z(n14702) );
  XOR U24783 ( .A(n15326), .B(n15327), .Z(n14700) );
  ANDN U24784 ( .B(n15328), .A(n15329), .Z(n15326) );
  AND U24785 ( .A(a[57]), .B(b[48]), .Z(n15325) );
  XNOR U24786 ( .A(n15330), .B(n14705), .Z(n14707) );
  XOR U24787 ( .A(n15331), .B(n15332), .Z(n14705) );
  ANDN U24788 ( .B(n15333), .A(n15334), .Z(n15331) );
  AND U24789 ( .A(a[58]), .B(b[47]), .Z(n15330) );
  XNOR U24790 ( .A(n15335), .B(n14710), .Z(n14712) );
  XOR U24791 ( .A(n15336), .B(n15337), .Z(n14710) );
  ANDN U24792 ( .B(n15338), .A(n15339), .Z(n15336) );
  AND U24793 ( .A(a[59]), .B(b[46]), .Z(n15335) );
  XNOR U24794 ( .A(n15340), .B(n14715), .Z(n14717) );
  XOR U24795 ( .A(n15341), .B(n15342), .Z(n14715) );
  ANDN U24796 ( .B(n15343), .A(n15344), .Z(n15341) );
  AND U24797 ( .A(a[60]), .B(b[45]), .Z(n15340) );
  XNOR U24798 ( .A(n15345), .B(n14720), .Z(n14722) );
  XOR U24799 ( .A(n15346), .B(n15347), .Z(n14720) );
  ANDN U24800 ( .B(n15348), .A(n15349), .Z(n15346) );
  AND U24801 ( .A(a[61]), .B(b[44]), .Z(n15345) );
  XNOR U24802 ( .A(n15350), .B(n14725), .Z(n14727) );
  XOR U24803 ( .A(n15351), .B(n15352), .Z(n14725) );
  ANDN U24804 ( .B(n15353), .A(n15354), .Z(n15351) );
  AND U24805 ( .A(a[62]), .B(b[43]), .Z(n15350) );
  XNOR U24806 ( .A(n15355), .B(n14730), .Z(n14732) );
  XOR U24807 ( .A(n15356), .B(n15357), .Z(n14730) );
  ANDN U24808 ( .B(n15358), .A(n15359), .Z(n15356) );
  AND U24809 ( .A(a[63]), .B(b[42]), .Z(n15355) );
  XNOR U24810 ( .A(n15360), .B(n14735), .Z(n14737) );
  XOR U24811 ( .A(n15361), .B(n15362), .Z(n14735) );
  ANDN U24812 ( .B(n15363), .A(n15364), .Z(n15361) );
  AND U24813 ( .A(a[64]), .B(b[41]), .Z(n15360) );
  XNOR U24814 ( .A(n15365), .B(n14740), .Z(n14742) );
  XOR U24815 ( .A(n15366), .B(n15367), .Z(n14740) );
  ANDN U24816 ( .B(n15368), .A(n15369), .Z(n15366) );
  AND U24817 ( .A(a[65]), .B(b[40]), .Z(n15365) );
  XNOR U24818 ( .A(n15370), .B(n14745), .Z(n14747) );
  XOR U24819 ( .A(n15371), .B(n15372), .Z(n14745) );
  ANDN U24820 ( .B(n15373), .A(n15374), .Z(n15371) );
  AND U24821 ( .A(a[66]), .B(b[39]), .Z(n15370) );
  XNOR U24822 ( .A(n15375), .B(n14750), .Z(n14752) );
  XOR U24823 ( .A(n15376), .B(n15377), .Z(n14750) );
  ANDN U24824 ( .B(n15378), .A(n15379), .Z(n15376) );
  AND U24825 ( .A(a[67]), .B(b[38]), .Z(n15375) );
  XNOR U24826 ( .A(n15380), .B(n14755), .Z(n14757) );
  XOR U24827 ( .A(n15381), .B(n15382), .Z(n14755) );
  ANDN U24828 ( .B(n15383), .A(n15384), .Z(n15381) );
  AND U24829 ( .A(a[68]), .B(b[37]), .Z(n15380) );
  XNOR U24830 ( .A(n15385), .B(n14760), .Z(n14762) );
  XOR U24831 ( .A(n15386), .B(n15387), .Z(n14760) );
  ANDN U24832 ( .B(n15388), .A(n15389), .Z(n15386) );
  AND U24833 ( .A(a[69]), .B(b[36]), .Z(n15385) );
  XNOR U24834 ( .A(n15390), .B(n14765), .Z(n14767) );
  XOR U24835 ( .A(n15391), .B(n15392), .Z(n14765) );
  ANDN U24836 ( .B(n15393), .A(n15394), .Z(n15391) );
  AND U24837 ( .A(a[70]), .B(b[35]), .Z(n15390) );
  XNOR U24838 ( .A(n15395), .B(n14770), .Z(n14772) );
  XOR U24839 ( .A(n15396), .B(n15397), .Z(n14770) );
  ANDN U24840 ( .B(n15398), .A(n15399), .Z(n15396) );
  AND U24841 ( .A(a[71]), .B(b[34]), .Z(n15395) );
  XNOR U24842 ( .A(n15400), .B(n14775), .Z(n14777) );
  XOR U24843 ( .A(n15401), .B(n15402), .Z(n14775) );
  ANDN U24844 ( .B(n15403), .A(n15404), .Z(n15401) );
  AND U24845 ( .A(a[72]), .B(b[33]), .Z(n15400) );
  XNOR U24846 ( .A(n15405), .B(n14780), .Z(n14782) );
  XOR U24847 ( .A(n15406), .B(n15407), .Z(n14780) );
  ANDN U24848 ( .B(n15408), .A(n15409), .Z(n15406) );
  AND U24849 ( .A(a[73]), .B(b[32]), .Z(n15405) );
  XNOR U24850 ( .A(n15410), .B(n14785), .Z(n14787) );
  XOR U24851 ( .A(n15411), .B(n15412), .Z(n14785) );
  ANDN U24852 ( .B(n15413), .A(n15414), .Z(n15411) );
  AND U24853 ( .A(a[74]), .B(b[31]), .Z(n15410) );
  XNOR U24854 ( .A(n15415), .B(n14790), .Z(n14792) );
  XOR U24855 ( .A(n15416), .B(n15417), .Z(n14790) );
  ANDN U24856 ( .B(n15418), .A(n15419), .Z(n15416) );
  AND U24857 ( .A(a[75]), .B(b[30]), .Z(n15415) );
  XNOR U24858 ( .A(n15420), .B(n14795), .Z(n14797) );
  XOR U24859 ( .A(n15421), .B(n15422), .Z(n14795) );
  ANDN U24860 ( .B(n15423), .A(n15424), .Z(n15421) );
  AND U24861 ( .A(a[76]), .B(b[29]), .Z(n15420) );
  XNOR U24862 ( .A(n15425), .B(n14800), .Z(n14802) );
  XOR U24863 ( .A(n15426), .B(n15427), .Z(n14800) );
  ANDN U24864 ( .B(n15428), .A(n15429), .Z(n15426) );
  AND U24865 ( .A(a[77]), .B(b[28]), .Z(n15425) );
  XNOR U24866 ( .A(n15430), .B(n14805), .Z(n14807) );
  XOR U24867 ( .A(n15431), .B(n15432), .Z(n14805) );
  ANDN U24868 ( .B(n15433), .A(n15434), .Z(n15431) );
  AND U24869 ( .A(a[78]), .B(b[27]), .Z(n15430) );
  XNOR U24870 ( .A(n15435), .B(n14810), .Z(n14812) );
  XOR U24871 ( .A(n15436), .B(n15437), .Z(n14810) );
  ANDN U24872 ( .B(n15438), .A(n15439), .Z(n15436) );
  AND U24873 ( .A(a[79]), .B(b[26]), .Z(n15435) );
  XNOR U24874 ( .A(n15440), .B(n14815), .Z(n14817) );
  XOR U24875 ( .A(n15441), .B(n15442), .Z(n14815) );
  ANDN U24876 ( .B(n15443), .A(n15444), .Z(n15441) );
  AND U24877 ( .A(a[80]), .B(b[25]), .Z(n15440) );
  XNOR U24878 ( .A(n15445), .B(n14820), .Z(n14822) );
  XOR U24879 ( .A(n15446), .B(n15447), .Z(n14820) );
  ANDN U24880 ( .B(n15448), .A(n15449), .Z(n15446) );
  AND U24881 ( .A(a[81]), .B(b[24]), .Z(n15445) );
  XNOR U24882 ( .A(n15450), .B(n14825), .Z(n14827) );
  XOR U24883 ( .A(n15451), .B(n15452), .Z(n14825) );
  ANDN U24884 ( .B(n15453), .A(n15454), .Z(n15451) );
  AND U24885 ( .A(a[82]), .B(b[23]), .Z(n15450) );
  XNOR U24886 ( .A(n15455), .B(n14830), .Z(n14832) );
  XOR U24887 ( .A(n15456), .B(n15457), .Z(n14830) );
  ANDN U24888 ( .B(n15458), .A(n15459), .Z(n15456) );
  AND U24889 ( .A(a[83]), .B(b[22]), .Z(n15455) );
  XNOR U24890 ( .A(n15460), .B(n14835), .Z(n14837) );
  XOR U24891 ( .A(n15461), .B(n15462), .Z(n14835) );
  ANDN U24892 ( .B(n15463), .A(n15464), .Z(n15461) );
  AND U24893 ( .A(a[84]), .B(b[21]), .Z(n15460) );
  XNOR U24894 ( .A(n15465), .B(n14840), .Z(n14842) );
  XOR U24895 ( .A(n15466), .B(n15467), .Z(n14840) );
  ANDN U24896 ( .B(n15468), .A(n15469), .Z(n15466) );
  AND U24897 ( .A(a[85]), .B(b[20]), .Z(n15465) );
  XNOR U24898 ( .A(n15470), .B(n14845), .Z(n14847) );
  XOR U24899 ( .A(n15471), .B(n15472), .Z(n14845) );
  ANDN U24900 ( .B(n15473), .A(n15474), .Z(n15471) );
  AND U24901 ( .A(a[86]), .B(b[19]), .Z(n15470) );
  XNOR U24902 ( .A(n15475), .B(n14850), .Z(n14852) );
  XOR U24903 ( .A(n15476), .B(n15477), .Z(n14850) );
  ANDN U24904 ( .B(n15478), .A(n15479), .Z(n15476) );
  AND U24905 ( .A(a[87]), .B(b[18]), .Z(n15475) );
  XNOR U24906 ( .A(n15480), .B(n14855), .Z(n14857) );
  XOR U24907 ( .A(n15481), .B(n15482), .Z(n14855) );
  ANDN U24908 ( .B(n15483), .A(n15484), .Z(n15481) );
  AND U24909 ( .A(a[88]), .B(b[17]), .Z(n15480) );
  XNOR U24910 ( .A(n15485), .B(n14860), .Z(n14862) );
  XOR U24911 ( .A(n15486), .B(n15487), .Z(n14860) );
  ANDN U24912 ( .B(n15488), .A(n15489), .Z(n15486) );
  AND U24913 ( .A(a[89]), .B(b[16]), .Z(n15485) );
  XNOR U24914 ( .A(n15490), .B(n14865), .Z(n14867) );
  XOR U24915 ( .A(n15491), .B(n15492), .Z(n14865) );
  ANDN U24916 ( .B(n15493), .A(n15494), .Z(n15491) );
  AND U24917 ( .A(a[90]), .B(b[15]), .Z(n15490) );
  XNOR U24918 ( .A(n15495), .B(n14870), .Z(n14872) );
  XOR U24919 ( .A(n15496), .B(n15497), .Z(n14870) );
  ANDN U24920 ( .B(n15498), .A(n15499), .Z(n15496) );
  AND U24921 ( .A(a[91]), .B(b[14]), .Z(n15495) );
  XNOR U24922 ( .A(n15500), .B(n14875), .Z(n14877) );
  XOR U24923 ( .A(n15501), .B(n15502), .Z(n14875) );
  ANDN U24924 ( .B(n15503), .A(n15504), .Z(n15501) );
  AND U24925 ( .A(a[92]), .B(b[13]), .Z(n15500) );
  XNOR U24926 ( .A(n15505), .B(n14880), .Z(n14882) );
  XOR U24927 ( .A(n15506), .B(n15507), .Z(n14880) );
  ANDN U24928 ( .B(n15508), .A(n15509), .Z(n15506) );
  AND U24929 ( .A(a[93]), .B(b[12]), .Z(n15505) );
  XNOR U24930 ( .A(n15510), .B(n14885), .Z(n14887) );
  XOR U24931 ( .A(n15511), .B(n15512), .Z(n14885) );
  ANDN U24932 ( .B(n15513), .A(n15514), .Z(n15511) );
  AND U24933 ( .A(a[94]), .B(b[11]), .Z(n15510) );
  XNOR U24934 ( .A(n15515), .B(n14890), .Z(n14892) );
  XOR U24935 ( .A(n15516), .B(n15517), .Z(n14890) );
  ANDN U24936 ( .B(n15518), .A(n15519), .Z(n15516) );
  AND U24937 ( .A(a[95]), .B(b[10]), .Z(n15515) );
  XNOR U24938 ( .A(n15520), .B(n14895), .Z(n14897) );
  XOR U24939 ( .A(n15521), .B(n15522), .Z(n14895) );
  ANDN U24940 ( .B(n15523), .A(n15524), .Z(n15521) );
  AND U24941 ( .A(b[9]), .B(a[96]), .Z(n15520) );
  XNOR U24942 ( .A(n15525), .B(n14900), .Z(n14902) );
  XOR U24943 ( .A(n15526), .B(n15527), .Z(n14900) );
  ANDN U24944 ( .B(n15528), .A(n15529), .Z(n15526) );
  AND U24945 ( .A(b[8]), .B(a[97]), .Z(n15525) );
  XNOR U24946 ( .A(n15530), .B(n14905), .Z(n14907) );
  XOR U24947 ( .A(n15531), .B(n15532), .Z(n14905) );
  ANDN U24948 ( .B(n15533), .A(n15534), .Z(n15531) );
  AND U24949 ( .A(b[7]), .B(a[98]), .Z(n15530) );
  XNOR U24950 ( .A(n15535), .B(n14910), .Z(n14912) );
  XOR U24951 ( .A(n15536), .B(n15537), .Z(n14910) );
  ANDN U24952 ( .B(n15538), .A(n15539), .Z(n15536) );
  AND U24953 ( .A(b[6]), .B(a[99]), .Z(n15535) );
  XNOR U24954 ( .A(n15540), .B(n14915), .Z(n14917) );
  XOR U24955 ( .A(n15541), .B(n15542), .Z(n14915) );
  ANDN U24956 ( .B(n15543), .A(n15544), .Z(n15541) );
  AND U24957 ( .A(b[5]), .B(a[100]), .Z(n15540) );
  XNOR U24958 ( .A(n15545), .B(n14920), .Z(n14922) );
  XOR U24959 ( .A(n15546), .B(n15547), .Z(n14920) );
  ANDN U24960 ( .B(n15548), .A(n15549), .Z(n15546) );
  AND U24961 ( .A(b[4]), .B(a[101]), .Z(n15545) );
  XNOR U24962 ( .A(n15550), .B(n15551), .Z(n14934) );
  NANDN U24963 ( .A(n15552), .B(n15553), .Z(n15551) );
  XNOR U24964 ( .A(n15554), .B(n14925), .Z(n14927) );
  XNOR U24965 ( .A(n15555), .B(n15556), .Z(n14925) );
  AND U24966 ( .A(n15557), .B(n15558), .Z(n15555) );
  AND U24967 ( .A(b[3]), .B(a[102]), .Z(n15554) );
  NAND U24968 ( .A(a[105]), .B(b[0]), .Z(n14312) );
  XNOR U24969 ( .A(n14940), .B(n14941), .Z(c[104]) );
  XNOR U24970 ( .A(n15552), .B(n15553), .Z(n14941) );
  XOR U24971 ( .A(n15550), .B(n15559), .Z(n15553) );
  NAND U24972 ( .A(b[1]), .B(a[103]), .Z(n15559) );
  XOR U24973 ( .A(n15558), .B(n15560), .Z(n15552) );
  XOR U24974 ( .A(n15550), .B(n15557), .Z(n15560) );
  XNOR U24975 ( .A(n15561), .B(n15556), .Z(n15557) );
  AND U24976 ( .A(b[2]), .B(a[102]), .Z(n15561) );
  NANDN U24977 ( .A(n15562), .B(n15563), .Z(n15550) );
  XOR U24978 ( .A(n15556), .B(n15548), .Z(n15564) );
  XNOR U24979 ( .A(n15547), .B(n15543), .Z(n15565) );
  XNOR U24980 ( .A(n15542), .B(n15538), .Z(n15566) );
  XNOR U24981 ( .A(n15537), .B(n15533), .Z(n15567) );
  XNOR U24982 ( .A(n15532), .B(n15528), .Z(n15568) );
  XNOR U24983 ( .A(n15527), .B(n15523), .Z(n15569) );
  XNOR U24984 ( .A(n15522), .B(n15518), .Z(n15570) );
  XNOR U24985 ( .A(n15517), .B(n15513), .Z(n15571) );
  XNOR U24986 ( .A(n15512), .B(n15508), .Z(n15572) );
  XNOR U24987 ( .A(n15507), .B(n15503), .Z(n15573) );
  XNOR U24988 ( .A(n15502), .B(n15498), .Z(n15574) );
  XNOR U24989 ( .A(n15497), .B(n15493), .Z(n15575) );
  XNOR U24990 ( .A(n15492), .B(n15488), .Z(n15576) );
  XNOR U24991 ( .A(n15487), .B(n15483), .Z(n15577) );
  XNOR U24992 ( .A(n15482), .B(n15478), .Z(n15578) );
  XNOR U24993 ( .A(n15477), .B(n15473), .Z(n15579) );
  XNOR U24994 ( .A(n15472), .B(n15468), .Z(n15580) );
  XNOR U24995 ( .A(n15467), .B(n15463), .Z(n15581) );
  XNOR U24996 ( .A(n15462), .B(n15458), .Z(n15582) );
  XNOR U24997 ( .A(n15457), .B(n15453), .Z(n15583) );
  XNOR U24998 ( .A(n15452), .B(n15448), .Z(n15584) );
  XNOR U24999 ( .A(n15447), .B(n15443), .Z(n15585) );
  XNOR U25000 ( .A(n15442), .B(n15438), .Z(n15586) );
  XNOR U25001 ( .A(n15437), .B(n15433), .Z(n15587) );
  XNOR U25002 ( .A(n15432), .B(n15428), .Z(n15588) );
  XNOR U25003 ( .A(n15427), .B(n15423), .Z(n15589) );
  XNOR U25004 ( .A(n15422), .B(n15418), .Z(n15590) );
  XNOR U25005 ( .A(n15417), .B(n15413), .Z(n15591) );
  XNOR U25006 ( .A(n15412), .B(n15408), .Z(n15592) );
  XNOR U25007 ( .A(n15407), .B(n15403), .Z(n15593) );
  XNOR U25008 ( .A(n15402), .B(n15398), .Z(n15594) );
  XNOR U25009 ( .A(n15397), .B(n15393), .Z(n15595) );
  XNOR U25010 ( .A(n15392), .B(n15388), .Z(n15596) );
  XNOR U25011 ( .A(n15387), .B(n15383), .Z(n15597) );
  XNOR U25012 ( .A(n15382), .B(n15378), .Z(n15598) );
  XNOR U25013 ( .A(n15377), .B(n15373), .Z(n15599) );
  XNOR U25014 ( .A(n15372), .B(n15368), .Z(n15600) );
  XNOR U25015 ( .A(n15367), .B(n15363), .Z(n15601) );
  XNOR U25016 ( .A(n15362), .B(n15358), .Z(n15602) );
  XNOR U25017 ( .A(n15357), .B(n15353), .Z(n15603) );
  XNOR U25018 ( .A(n15352), .B(n15348), .Z(n15604) );
  XNOR U25019 ( .A(n15347), .B(n15343), .Z(n15605) );
  XNOR U25020 ( .A(n15342), .B(n15338), .Z(n15606) );
  XNOR U25021 ( .A(n15337), .B(n15333), .Z(n15607) );
  XNOR U25022 ( .A(n15332), .B(n15328), .Z(n15608) );
  XNOR U25023 ( .A(n15327), .B(n15323), .Z(n15609) );
  XNOR U25024 ( .A(n15322), .B(n15318), .Z(n15610) );
  XNOR U25025 ( .A(n15317), .B(n15313), .Z(n15611) );
  XNOR U25026 ( .A(n15312), .B(n15308), .Z(n15612) );
  XNOR U25027 ( .A(n15307), .B(n15303), .Z(n15613) );
  XNOR U25028 ( .A(n15302), .B(n15298), .Z(n15614) );
  XNOR U25029 ( .A(n15297), .B(n15293), .Z(n15615) );
  XNOR U25030 ( .A(n15292), .B(n15288), .Z(n15616) );
  XNOR U25031 ( .A(n15287), .B(n15283), .Z(n15617) );
  XNOR U25032 ( .A(n15282), .B(n15278), .Z(n15618) );
  XNOR U25033 ( .A(n15277), .B(n15273), .Z(n15619) );
  XNOR U25034 ( .A(n15272), .B(n15268), .Z(n15620) );
  XNOR U25035 ( .A(n15267), .B(n15263), .Z(n15621) );
  XNOR U25036 ( .A(n15262), .B(n15258), .Z(n15622) );
  XNOR U25037 ( .A(n15257), .B(n15253), .Z(n15623) );
  XNOR U25038 ( .A(n15252), .B(n15248), .Z(n15624) );
  XNOR U25039 ( .A(n15247), .B(n15243), .Z(n15625) );
  XNOR U25040 ( .A(n15242), .B(n15238), .Z(n15626) );
  XNOR U25041 ( .A(n15237), .B(n15233), .Z(n15627) );
  XNOR U25042 ( .A(n15232), .B(n15228), .Z(n15628) );
  XNOR U25043 ( .A(n15227), .B(n15223), .Z(n15629) );
  XNOR U25044 ( .A(n15222), .B(n15218), .Z(n15630) );
  XNOR U25045 ( .A(n15217), .B(n15213), .Z(n15631) );
  XNOR U25046 ( .A(n15212), .B(n15208), .Z(n15632) );
  XNOR U25047 ( .A(n15207), .B(n15203), .Z(n15633) );
  XNOR U25048 ( .A(n15202), .B(n15198), .Z(n15634) );
  XNOR U25049 ( .A(n15197), .B(n15193), .Z(n15635) );
  XNOR U25050 ( .A(n15192), .B(n15188), .Z(n15636) );
  XNOR U25051 ( .A(n15187), .B(n15183), .Z(n15637) );
  XNOR U25052 ( .A(n15182), .B(n15178), .Z(n15638) );
  XNOR U25053 ( .A(n15177), .B(n15173), .Z(n15639) );
  XNOR U25054 ( .A(n15172), .B(n15168), .Z(n15640) );
  XNOR U25055 ( .A(n15167), .B(n15163), .Z(n15641) );
  XNOR U25056 ( .A(n15162), .B(n15158), .Z(n15642) );
  XNOR U25057 ( .A(n15157), .B(n15153), .Z(n15643) );
  XNOR U25058 ( .A(n15152), .B(n15148), .Z(n15644) );
  XNOR U25059 ( .A(n15147), .B(n15143), .Z(n15645) );
  XNOR U25060 ( .A(n15142), .B(n15138), .Z(n15646) );
  XNOR U25061 ( .A(n15137), .B(n15133), .Z(n15647) );
  XNOR U25062 ( .A(n15132), .B(n15128), .Z(n15648) );
  XNOR U25063 ( .A(n15127), .B(n15123), .Z(n15649) );
  XNOR U25064 ( .A(n15122), .B(n15118), .Z(n15650) );
  XNOR U25065 ( .A(n15117), .B(n15113), .Z(n15651) );
  XNOR U25066 ( .A(n15112), .B(n15108), .Z(n15652) );
  XNOR U25067 ( .A(n15107), .B(n15103), .Z(n15653) );
  XNOR U25068 ( .A(n15102), .B(n15098), .Z(n15654) );
  XNOR U25069 ( .A(n15097), .B(n15093), .Z(n15655) );
  XNOR U25070 ( .A(n15092), .B(n15088), .Z(n15656) );
  XNOR U25071 ( .A(n15087), .B(n15083), .Z(n15657) );
  XNOR U25072 ( .A(n15082), .B(n15078), .Z(n15658) );
  XNOR U25073 ( .A(n15077), .B(n15073), .Z(n15659) );
  XNOR U25074 ( .A(n15072), .B(n15068), .Z(n15660) );
  XNOR U25075 ( .A(n15067), .B(n15063), .Z(n15661) );
  XNOR U25076 ( .A(n15062), .B(n15058), .Z(n15662) );
  XNOR U25077 ( .A(n15057), .B(n15053), .Z(n15663) );
  XNOR U25078 ( .A(n15052), .B(n15048), .Z(n15664) );
  XOR U25079 ( .A(n15665), .B(n15047), .Z(n15048) );
  AND U25080 ( .A(a[0]), .B(b[104]), .Z(n15665) );
  XNOR U25081 ( .A(n15666), .B(n15047), .Z(n15049) );
  XNOR U25082 ( .A(n15667), .B(n15668), .Z(n15047) );
  ANDN U25083 ( .B(n15669), .A(n15670), .Z(n15667) );
  AND U25084 ( .A(a[1]), .B(b[103]), .Z(n15666) );
  XNOR U25085 ( .A(n15671), .B(n15052), .Z(n15054) );
  XOR U25086 ( .A(n15672), .B(n15673), .Z(n15052) );
  ANDN U25087 ( .B(n15674), .A(n15675), .Z(n15672) );
  AND U25088 ( .A(a[2]), .B(b[102]), .Z(n15671) );
  XNOR U25089 ( .A(n15676), .B(n15057), .Z(n15059) );
  XOR U25090 ( .A(n15677), .B(n15678), .Z(n15057) );
  ANDN U25091 ( .B(n15679), .A(n15680), .Z(n15677) );
  AND U25092 ( .A(a[3]), .B(b[101]), .Z(n15676) );
  XNOR U25093 ( .A(n15681), .B(n15062), .Z(n15064) );
  XOR U25094 ( .A(n15682), .B(n15683), .Z(n15062) );
  ANDN U25095 ( .B(n15684), .A(n15685), .Z(n15682) );
  AND U25096 ( .A(a[4]), .B(b[100]), .Z(n15681) );
  XNOR U25097 ( .A(n15686), .B(n15067), .Z(n15069) );
  XOR U25098 ( .A(n15687), .B(n15688), .Z(n15067) );
  ANDN U25099 ( .B(n15689), .A(n15690), .Z(n15687) );
  AND U25100 ( .A(a[5]), .B(b[99]), .Z(n15686) );
  XNOR U25101 ( .A(n15691), .B(n15072), .Z(n15074) );
  XOR U25102 ( .A(n15692), .B(n15693), .Z(n15072) );
  ANDN U25103 ( .B(n15694), .A(n15695), .Z(n15692) );
  AND U25104 ( .A(a[6]), .B(b[98]), .Z(n15691) );
  XNOR U25105 ( .A(n15696), .B(n15077), .Z(n15079) );
  XOR U25106 ( .A(n15697), .B(n15698), .Z(n15077) );
  ANDN U25107 ( .B(n15699), .A(n15700), .Z(n15697) );
  AND U25108 ( .A(a[7]), .B(b[97]), .Z(n15696) );
  XNOR U25109 ( .A(n15701), .B(n15082), .Z(n15084) );
  XOR U25110 ( .A(n15702), .B(n15703), .Z(n15082) );
  ANDN U25111 ( .B(n15704), .A(n15705), .Z(n15702) );
  AND U25112 ( .A(a[8]), .B(b[96]), .Z(n15701) );
  XNOR U25113 ( .A(n15706), .B(n15087), .Z(n15089) );
  XOR U25114 ( .A(n15707), .B(n15708), .Z(n15087) );
  ANDN U25115 ( .B(n15709), .A(n15710), .Z(n15707) );
  AND U25116 ( .A(a[9]), .B(b[95]), .Z(n15706) );
  XNOR U25117 ( .A(n15711), .B(n15092), .Z(n15094) );
  XOR U25118 ( .A(n15712), .B(n15713), .Z(n15092) );
  ANDN U25119 ( .B(n15714), .A(n15715), .Z(n15712) );
  AND U25120 ( .A(a[10]), .B(b[94]), .Z(n15711) );
  XNOR U25121 ( .A(n15716), .B(n15097), .Z(n15099) );
  XOR U25122 ( .A(n15717), .B(n15718), .Z(n15097) );
  ANDN U25123 ( .B(n15719), .A(n15720), .Z(n15717) );
  AND U25124 ( .A(a[11]), .B(b[93]), .Z(n15716) );
  XNOR U25125 ( .A(n15721), .B(n15102), .Z(n15104) );
  XOR U25126 ( .A(n15722), .B(n15723), .Z(n15102) );
  ANDN U25127 ( .B(n15724), .A(n15725), .Z(n15722) );
  AND U25128 ( .A(a[12]), .B(b[92]), .Z(n15721) );
  XNOR U25129 ( .A(n15726), .B(n15107), .Z(n15109) );
  XOR U25130 ( .A(n15727), .B(n15728), .Z(n15107) );
  ANDN U25131 ( .B(n15729), .A(n15730), .Z(n15727) );
  AND U25132 ( .A(a[13]), .B(b[91]), .Z(n15726) );
  XNOR U25133 ( .A(n15731), .B(n15112), .Z(n15114) );
  XOR U25134 ( .A(n15732), .B(n15733), .Z(n15112) );
  ANDN U25135 ( .B(n15734), .A(n15735), .Z(n15732) );
  AND U25136 ( .A(a[14]), .B(b[90]), .Z(n15731) );
  XNOR U25137 ( .A(n15736), .B(n15117), .Z(n15119) );
  XOR U25138 ( .A(n15737), .B(n15738), .Z(n15117) );
  ANDN U25139 ( .B(n15739), .A(n15740), .Z(n15737) );
  AND U25140 ( .A(a[15]), .B(b[89]), .Z(n15736) );
  XNOR U25141 ( .A(n15741), .B(n15122), .Z(n15124) );
  XOR U25142 ( .A(n15742), .B(n15743), .Z(n15122) );
  ANDN U25143 ( .B(n15744), .A(n15745), .Z(n15742) );
  AND U25144 ( .A(a[16]), .B(b[88]), .Z(n15741) );
  XNOR U25145 ( .A(n15746), .B(n15127), .Z(n15129) );
  XOR U25146 ( .A(n15747), .B(n15748), .Z(n15127) );
  ANDN U25147 ( .B(n15749), .A(n15750), .Z(n15747) );
  AND U25148 ( .A(a[17]), .B(b[87]), .Z(n15746) );
  XNOR U25149 ( .A(n15751), .B(n15132), .Z(n15134) );
  XOR U25150 ( .A(n15752), .B(n15753), .Z(n15132) );
  ANDN U25151 ( .B(n15754), .A(n15755), .Z(n15752) );
  AND U25152 ( .A(a[18]), .B(b[86]), .Z(n15751) );
  XNOR U25153 ( .A(n15756), .B(n15137), .Z(n15139) );
  XOR U25154 ( .A(n15757), .B(n15758), .Z(n15137) );
  ANDN U25155 ( .B(n15759), .A(n15760), .Z(n15757) );
  AND U25156 ( .A(a[19]), .B(b[85]), .Z(n15756) );
  XNOR U25157 ( .A(n15761), .B(n15142), .Z(n15144) );
  XOR U25158 ( .A(n15762), .B(n15763), .Z(n15142) );
  ANDN U25159 ( .B(n15764), .A(n15765), .Z(n15762) );
  AND U25160 ( .A(a[20]), .B(b[84]), .Z(n15761) );
  XNOR U25161 ( .A(n15766), .B(n15147), .Z(n15149) );
  XOR U25162 ( .A(n15767), .B(n15768), .Z(n15147) );
  ANDN U25163 ( .B(n15769), .A(n15770), .Z(n15767) );
  AND U25164 ( .A(a[21]), .B(b[83]), .Z(n15766) );
  XNOR U25165 ( .A(n15771), .B(n15152), .Z(n15154) );
  XOR U25166 ( .A(n15772), .B(n15773), .Z(n15152) );
  ANDN U25167 ( .B(n15774), .A(n15775), .Z(n15772) );
  AND U25168 ( .A(a[22]), .B(b[82]), .Z(n15771) );
  XNOR U25169 ( .A(n15776), .B(n15157), .Z(n15159) );
  XOR U25170 ( .A(n15777), .B(n15778), .Z(n15157) );
  ANDN U25171 ( .B(n15779), .A(n15780), .Z(n15777) );
  AND U25172 ( .A(a[23]), .B(b[81]), .Z(n15776) );
  XNOR U25173 ( .A(n15781), .B(n15162), .Z(n15164) );
  XOR U25174 ( .A(n15782), .B(n15783), .Z(n15162) );
  ANDN U25175 ( .B(n15784), .A(n15785), .Z(n15782) );
  AND U25176 ( .A(a[24]), .B(b[80]), .Z(n15781) );
  XNOR U25177 ( .A(n15786), .B(n15167), .Z(n15169) );
  XOR U25178 ( .A(n15787), .B(n15788), .Z(n15167) );
  ANDN U25179 ( .B(n15789), .A(n15790), .Z(n15787) );
  AND U25180 ( .A(a[25]), .B(b[79]), .Z(n15786) );
  XNOR U25181 ( .A(n15791), .B(n15172), .Z(n15174) );
  XOR U25182 ( .A(n15792), .B(n15793), .Z(n15172) );
  ANDN U25183 ( .B(n15794), .A(n15795), .Z(n15792) );
  AND U25184 ( .A(a[26]), .B(b[78]), .Z(n15791) );
  XNOR U25185 ( .A(n15796), .B(n15177), .Z(n15179) );
  XOR U25186 ( .A(n15797), .B(n15798), .Z(n15177) );
  ANDN U25187 ( .B(n15799), .A(n15800), .Z(n15797) );
  AND U25188 ( .A(a[27]), .B(b[77]), .Z(n15796) );
  XNOR U25189 ( .A(n15801), .B(n15182), .Z(n15184) );
  XOR U25190 ( .A(n15802), .B(n15803), .Z(n15182) );
  ANDN U25191 ( .B(n15804), .A(n15805), .Z(n15802) );
  AND U25192 ( .A(a[28]), .B(b[76]), .Z(n15801) );
  XNOR U25193 ( .A(n15806), .B(n15187), .Z(n15189) );
  XOR U25194 ( .A(n15807), .B(n15808), .Z(n15187) );
  ANDN U25195 ( .B(n15809), .A(n15810), .Z(n15807) );
  AND U25196 ( .A(a[29]), .B(b[75]), .Z(n15806) );
  XNOR U25197 ( .A(n15811), .B(n15192), .Z(n15194) );
  XOR U25198 ( .A(n15812), .B(n15813), .Z(n15192) );
  ANDN U25199 ( .B(n15814), .A(n15815), .Z(n15812) );
  AND U25200 ( .A(a[30]), .B(b[74]), .Z(n15811) );
  XNOR U25201 ( .A(n15816), .B(n15197), .Z(n15199) );
  XOR U25202 ( .A(n15817), .B(n15818), .Z(n15197) );
  ANDN U25203 ( .B(n15819), .A(n15820), .Z(n15817) );
  AND U25204 ( .A(a[31]), .B(b[73]), .Z(n15816) );
  XNOR U25205 ( .A(n15821), .B(n15202), .Z(n15204) );
  XOR U25206 ( .A(n15822), .B(n15823), .Z(n15202) );
  ANDN U25207 ( .B(n15824), .A(n15825), .Z(n15822) );
  AND U25208 ( .A(a[32]), .B(b[72]), .Z(n15821) );
  XNOR U25209 ( .A(n15826), .B(n15207), .Z(n15209) );
  XOR U25210 ( .A(n15827), .B(n15828), .Z(n15207) );
  ANDN U25211 ( .B(n15829), .A(n15830), .Z(n15827) );
  AND U25212 ( .A(a[33]), .B(b[71]), .Z(n15826) );
  XNOR U25213 ( .A(n15831), .B(n15212), .Z(n15214) );
  XOR U25214 ( .A(n15832), .B(n15833), .Z(n15212) );
  ANDN U25215 ( .B(n15834), .A(n15835), .Z(n15832) );
  AND U25216 ( .A(a[34]), .B(b[70]), .Z(n15831) );
  XNOR U25217 ( .A(n15836), .B(n15217), .Z(n15219) );
  XOR U25218 ( .A(n15837), .B(n15838), .Z(n15217) );
  ANDN U25219 ( .B(n15839), .A(n15840), .Z(n15837) );
  AND U25220 ( .A(a[35]), .B(b[69]), .Z(n15836) );
  XNOR U25221 ( .A(n15841), .B(n15222), .Z(n15224) );
  XOR U25222 ( .A(n15842), .B(n15843), .Z(n15222) );
  ANDN U25223 ( .B(n15844), .A(n15845), .Z(n15842) );
  AND U25224 ( .A(a[36]), .B(b[68]), .Z(n15841) );
  XNOR U25225 ( .A(n15846), .B(n15227), .Z(n15229) );
  XOR U25226 ( .A(n15847), .B(n15848), .Z(n15227) );
  ANDN U25227 ( .B(n15849), .A(n15850), .Z(n15847) );
  AND U25228 ( .A(a[37]), .B(b[67]), .Z(n15846) );
  XNOR U25229 ( .A(n15851), .B(n15232), .Z(n15234) );
  XOR U25230 ( .A(n15852), .B(n15853), .Z(n15232) );
  ANDN U25231 ( .B(n15854), .A(n15855), .Z(n15852) );
  AND U25232 ( .A(a[38]), .B(b[66]), .Z(n15851) );
  XNOR U25233 ( .A(n15856), .B(n15237), .Z(n15239) );
  XOR U25234 ( .A(n15857), .B(n15858), .Z(n15237) );
  ANDN U25235 ( .B(n15859), .A(n15860), .Z(n15857) );
  AND U25236 ( .A(a[39]), .B(b[65]), .Z(n15856) );
  XNOR U25237 ( .A(n15861), .B(n15242), .Z(n15244) );
  XOR U25238 ( .A(n15862), .B(n15863), .Z(n15242) );
  ANDN U25239 ( .B(n15864), .A(n15865), .Z(n15862) );
  AND U25240 ( .A(a[40]), .B(b[64]), .Z(n15861) );
  XNOR U25241 ( .A(n15866), .B(n15247), .Z(n15249) );
  XOR U25242 ( .A(n15867), .B(n15868), .Z(n15247) );
  ANDN U25243 ( .B(n15869), .A(n15870), .Z(n15867) );
  AND U25244 ( .A(a[41]), .B(b[63]), .Z(n15866) );
  XNOR U25245 ( .A(n15871), .B(n15252), .Z(n15254) );
  XOR U25246 ( .A(n15872), .B(n15873), .Z(n15252) );
  ANDN U25247 ( .B(n15874), .A(n15875), .Z(n15872) );
  AND U25248 ( .A(a[42]), .B(b[62]), .Z(n15871) );
  XNOR U25249 ( .A(n15876), .B(n15257), .Z(n15259) );
  XOR U25250 ( .A(n15877), .B(n15878), .Z(n15257) );
  ANDN U25251 ( .B(n15879), .A(n15880), .Z(n15877) );
  AND U25252 ( .A(a[43]), .B(b[61]), .Z(n15876) );
  XNOR U25253 ( .A(n15881), .B(n15262), .Z(n15264) );
  XOR U25254 ( .A(n15882), .B(n15883), .Z(n15262) );
  ANDN U25255 ( .B(n15884), .A(n15885), .Z(n15882) );
  AND U25256 ( .A(a[44]), .B(b[60]), .Z(n15881) );
  XNOR U25257 ( .A(n15886), .B(n15267), .Z(n15269) );
  XOR U25258 ( .A(n15887), .B(n15888), .Z(n15267) );
  ANDN U25259 ( .B(n15889), .A(n15890), .Z(n15887) );
  AND U25260 ( .A(a[45]), .B(b[59]), .Z(n15886) );
  XNOR U25261 ( .A(n15891), .B(n15272), .Z(n15274) );
  XOR U25262 ( .A(n15892), .B(n15893), .Z(n15272) );
  ANDN U25263 ( .B(n15894), .A(n15895), .Z(n15892) );
  AND U25264 ( .A(a[46]), .B(b[58]), .Z(n15891) );
  XNOR U25265 ( .A(n15896), .B(n15277), .Z(n15279) );
  XOR U25266 ( .A(n15897), .B(n15898), .Z(n15277) );
  ANDN U25267 ( .B(n15899), .A(n15900), .Z(n15897) );
  AND U25268 ( .A(a[47]), .B(b[57]), .Z(n15896) );
  XNOR U25269 ( .A(n15901), .B(n15282), .Z(n15284) );
  XOR U25270 ( .A(n15902), .B(n15903), .Z(n15282) );
  ANDN U25271 ( .B(n15904), .A(n15905), .Z(n15902) );
  AND U25272 ( .A(a[48]), .B(b[56]), .Z(n15901) );
  XNOR U25273 ( .A(n15906), .B(n15287), .Z(n15289) );
  XOR U25274 ( .A(n15907), .B(n15908), .Z(n15287) );
  ANDN U25275 ( .B(n15909), .A(n15910), .Z(n15907) );
  AND U25276 ( .A(a[49]), .B(b[55]), .Z(n15906) );
  XNOR U25277 ( .A(n15911), .B(n15292), .Z(n15294) );
  XOR U25278 ( .A(n15912), .B(n15913), .Z(n15292) );
  ANDN U25279 ( .B(n15914), .A(n15915), .Z(n15912) );
  AND U25280 ( .A(a[50]), .B(b[54]), .Z(n15911) );
  XNOR U25281 ( .A(n15916), .B(n15297), .Z(n15299) );
  XOR U25282 ( .A(n15917), .B(n15918), .Z(n15297) );
  ANDN U25283 ( .B(n15919), .A(n15920), .Z(n15917) );
  AND U25284 ( .A(a[51]), .B(b[53]), .Z(n15916) );
  XNOR U25285 ( .A(n15921), .B(n15302), .Z(n15304) );
  XOR U25286 ( .A(n15922), .B(n15923), .Z(n15302) );
  ANDN U25287 ( .B(n15924), .A(n15925), .Z(n15922) );
  AND U25288 ( .A(a[52]), .B(b[52]), .Z(n15921) );
  XNOR U25289 ( .A(n15926), .B(n15307), .Z(n15309) );
  XOR U25290 ( .A(n15927), .B(n15928), .Z(n15307) );
  ANDN U25291 ( .B(n15929), .A(n15930), .Z(n15927) );
  AND U25292 ( .A(a[53]), .B(b[51]), .Z(n15926) );
  XNOR U25293 ( .A(n15931), .B(n15312), .Z(n15314) );
  XOR U25294 ( .A(n15932), .B(n15933), .Z(n15312) );
  ANDN U25295 ( .B(n15934), .A(n15935), .Z(n15932) );
  AND U25296 ( .A(a[54]), .B(b[50]), .Z(n15931) );
  XNOR U25297 ( .A(n15936), .B(n15317), .Z(n15319) );
  XOR U25298 ( .A(n15937), .B(n15938), .Z(n15317) );
  ANDN U25299 ( .B(n15939), .A(n15940), .Z(n15937) );
  AND U25300 ( .A(a[55]), .B(b[49]), .Z(n15936) );
  XNOR U25301 ( .A(n15941), .B(n15322), .Z(n15324) );
  XOR U25302 ( .A(n15942), .B(n15943), .Z(n15322) );
  ANDN U25303 ( .B(n15944), .A(n15945), .Z(n15942) );
  AND U25304 ( .A(a[56]), .B(b[48]), .Z(n15941) );
  XNOR U25305 ( .A(n15946), .B(n15327), .Z(n15329) );
  XOR U25306 ( .A(n15947), .B(n15948), .Z(n15327) );
  ANDN U25307 ( .B(n15949), .A(n15950), .Z(n15947) );
  AND U25308 ( .A(a[57]), .B(b[47]), .Z(n15946) );
  XNOR U25309 ( .A(n15951), .B(n15332), .Z(n15334) );
  XOR U25310 ( .A(n15952), .B(n15953), .Z(n15332) );
  ANDN U25311 ( .B(n15954), .A(n15955), .Z(n15952) );
  AND U25312 ( .A(a[58]), .B(b[46]), .Z(n15951) );
  XNOR U25313 ( .A(n15956), .B(n15337), .Z(n15339) );
  XOR U25314 ( .A(n15957), .B(n15958), .Z(n15337) );
  ANDN U25315 ( .B(n15959), .A(n15960), .Z(n15957) );
  AND U25316 ( .A(a[59]), .B(b[45]), .Z(n15956) );
  XNOR U25317 ( .A(n15961), .B(n15342), .Z(n15344) );
  XOR U25318 ( .A(n15962), .B(n15963), .Z(n15342) );
  ANDN U25319 ( .B(n15964), .A(n15965), .Z(n15962) );
  AND U25320 ( .A(a[60]), .B(b[44]), .Z(n15961) );
  XNOR U25321 ( .A(n15966), .B(n15347), .Z(n15349) );
  XOR U25322 ( .A(n15967), .B(n15968), .Z(n15347) );
  ANDN U25323 ( .B(n15969), .A(n15970), .Z(n15967) );
  AND U25324 ( .A(a[61]), .B(b[43]), .Z(n15966) );
  XNOR U25325 ( .A(n15971), .B(n15352), .Z(n15354) );
  XOR U25326 ( .A(n15972), .B(n15973), .Z(n15352) );
  ANDN U25327 ( .B(n15974), .A(n15975), .Z(n15972) );
  AND U25328 ( .A(a[62]), .B(b[42]), .Z(n15971) );
  XNOR U25329 ( .A(n15976), .B(n15357), .Z(n15359) );
  XOR U25330 ( .A(n15977), .B(n15978), .Z(n15357) );
  ANDN U25331 ( .B(n15979), .A(n15980), .Z(n15977) );
  AND U25332 ( .A(a[63]), .B(b[41]), .Z(n15976) );
  XNOR U25333 ( .A(n15981), .B(n15362), .Z(n15364) );
  XOR U25334 ( .A(n15982), .B(n15983), .Z(n15362) );
  ANDN U25335 ( .B(n15984), .A(n15985), .Z(n15982) );
  AND U25336 ( .A(a[64]), .B(b[40]), .Z(n15981) );
  XNOR U25337 ( .A(n15986), .B(n15367), .Z(n15369) );
  XOR U25338 ( .A(n15987), .B(n15988), .Z(n15367) );
  ANDN U25339 ( .B(n15989), .A(n15990), .Z(n15987) );
  AND U25340 ( .A(a[65]), .B(b[39]), .Z(n15986) );
  XNOR U25341 ( .A(n15991), .B(n15372), .Z(n15374) );
  XOR U25342 ( .A(n15992), .B(n15993), .Z(n15372) );
  ANDN U25343 ( .B(n15994), .A(n15995), .Z(n15992) );
  AND U25344 ( .A(a[66]), .B(b[38]), .Z(n15991) );
  XNOR U25345 ( .A(n15996), .B(n15377), .Z(n15379) );
  XOR U25346 ( .A(n15997), .B(n15998), .Z(n15377) );
  ANDN U25347 ( .B(n15999), .A(n16000), .Z(n15997) );
  AND U25348 ( .A(a[67]), .B(b[37]), .Z(n15996) );
  XNOR U25349 ( .A(n16001), .B(n15382), .Z(n15384) );
  XOR U25350 ( .A(n16002), .B(n16003), .Z(n15382) );
  ANDN U25351 ( .B(n16004), .A(n16005), .Z(n16002) );
  AND U25352 ( .A(a[68]), .B(b[36]), .Z(n16001) );
  XNOR U25353 ( .A(n16006), .B(n15387), .Z(n15389) );
  XOR U25354 ( .A(n16007), .B(n16008), .Z(n15387) );
  ANDN U25355 ( .B(n16009), .A(n16010), .Z(n16007) );
  AND U25356 ( .A(a[69]), .B(b[35]), .Z(n16006) );
  XNOR U25357 ( .A(n16011), .B(n15392), .Z(n15394) );
  XOR U25358 ( .A(n16012), .B(n16013), .Z(n15392) );
  ANDN U25359 ( .B(n16014), .A(n16015), .Z(n16012) );
  AND U25360 ( .A(a[70]), .B(b[34]), .Z(n16011) );
  XNOR U25361 ( .A(n16016), .B(n15397), .Z(n15399) );
  XOR U25362 ( .A(n16017), .B(n16018), .Z(n15397) );
  ANDN U25363 ( .B(n16019), .A(n16020), .Z(n16017) );
  AND U25364 ( .A(a[71]), .B(b[33]), .Z(n16016) );
  XNOR U25365 ( .A(n16021), .B(n15402), .Z(n15404) );
  XOR U25366 ( .A(n16022), .B(n16023), .Z(n15402) );
  ANDN U25367 ( .B(n16024), .A(n16025), .Z(n16022) );
  AND U25368 ( .A(a[72]), .B(b[32]), .Z(n16021) );
  XNOR U25369 ( .A(n16026), .B(n15407), .Z(n15409) );
  XOR U25370 ( .A(n16027), .B(n16028), .Z(n15407) );
  ANDN U25371 ( .B(n16029), .A(n16030), .Z(n16027) );
  AND U25372 ( .A(a[73]), .B(b[31]), .Z(n16026) );
  XNOR U25373 ( .A(n16031), .B(n15412), .Z(n15414) );
  XOR U25374 ( .A(n16032), .B(n16033), .Z(n15412) );
  ANDN U25375 ( .B(n16034), .A(n16035), .Z(n16032) );
  AND U25376 ( .A(a[74]), .B(b[30]), .Z(n16031) );
  XNOR U25377 ( .A(n16036), .B(n15417), .Z(n15419) );
  XOR U25378 ( .A(n16037), .B(n16038), .Z(n15417) );
  ANDN U25379 ( .B(n16039), .A(n16040), .Z(n16037) );
  AND U25380 ( .A(a[75]), .B(b[29]), .Z(n16036) );
  XNOR U25381 ( .A(n16041), .B(n15422), .Z(n15424) );
  XOR U25382 ( .A(n16042), .B(n16043), .Z(n15422) );
  ANDN U25383 ( .B(n16044), .A(n16045), .Z(n16042) );
  AND U25384 ( .A(a[76]), .B(b[28]), .Z(n16041) );
  XNOR U25385 ( .A(n16046), .B(n15427), .Z(n15429) );
  XOR U25386 ( .A(n16047), .B(n16048), .Z(n15427) );
  ANDN U25387 ( .B(n16049), .A(n16050), .Z(n16047) );
  AND U25388 ( .A(a[77]), .B(b[27]), .Z(n16046) );
  XNOR U25389 ( .A(n16051), .B(n15432), .Z(n15434) );
  XOR U25390 ( .A(n16052), .B(n16053), .Z(n15432) );
  ANDN U25391 ( .B(n16054), .A(n16055), .Z(n16052) );
  AND U25392 ( .A(a[78]), .B(b[26]), .Z(n16051) );
  XNOR U25393 ( .A(n16056), .B(n15437), .Z(n15439) );
  XOR U25394 ( .A(n16057), .B(n16058), .Z(n15437) );
  ANDN U25395 ( .B(n16059), .A(n16060), .Z(n16057) );
  AND U25396 ( .A(a[79]), .B(b[25]), .Z(n16056) );
  XNOR U25397 ( .A(n16061), .B(n15442), .Z(n15444) );
  XOR U25398 ( .A(n16062), .B(n16063), .Z(n15442) );
  ANDN U25399 ( .B(n16064), .A(n16065), .Z(n16062) );
  AND U25400 ( .A(a[80]), .B(b[24]), .Z(n16061) );
  XNOR U25401 ( .A(n16066), .B(n15447), .Z(n15449) );
  XOR U25402 ( .A(n16067), .B(n16068), .Z(n15447) );
  ANDN U25403 ( .B(n16069), .A(n16070), .Z(n16067) );
  AND U25404 ( .A(a[81]), .B(b[23]), .Z(n16066) );
  XNOR U25405 ( .A(n16071), .B(n15452), .Z(n15454) );
  XOR U25406 ( .A(n16072), .B(n16073), .Z(n15452) );
  ANDN U25407 ( .B(n16074), .A(n16075), .Z(n16072) );
  AND U25408 ( .A(a[82]), .B(b[22]), .Z(n16071) );
  XNOR U25409 ( .A(n16076), .B(n15457), .Z(n15459) );
  XOR U25410 ( .A(n16077), .B(n16078), .Z(n15457) );
  ANDN U25411 ( .B(n16079), .A(n16080), .Z(n16077) );
  AND U25412 ( .A(a[83]), .B(b[21]), .Z(n16076) );
  XNOR U25413 ( .A(n16081), .B(n15462), .Z(n15464) );
  XOR U25414 ( .A(n16082), .B(n16083), .Z(n15462) );
  ANDN U25415 ( .B(n16084), .A(n16085), .Z(n16082) );
  AND U25416 ( .A(a[84]), .B(b[20]), .Z(n16081) );
  XNOR U25417 ( .A(n16086), .B(n15467), .Z(n15469) );
  XOR U25418 ( .A(n16087), .B(n16088), .Z(n15467) );
  ANDN U25419 ( .B(n16089), .A(n16090), .Z(n16087) );
  AND U25420 ( .A(a[85]), .B(b[19]), .Z(n16086) );
  XNOR U25421 ( .A(n16091), .B(n15472), .Z(n15474) );
  XOR U25422 ( .A(n16092), .B(n16093), .Z(n15472) );
  ANDN U25423 ( .B(n16094), .A(n16095), .Z(n16092) );
  AND U25424 ( .A(a[86]), .B(b[18]), .Z(n16091) );
  XNOR U25425 ( .A(n16096), .B(n15477), .Z(n15479) );
  XOR U25426 ( .A(n16097), .B(n16098), .Z(n15477) );
  ANDN U25427 ( .B(n16099), .A(n16100), .Z(n16097) );
  AND U25428 ( .A(a[87]), .B(b[17]), .Z(n16096) );
  XNOR U25429 ( .A(n16101), .B(n15482), .Z(n15484) );
  XOR U25430 ( .A(n16102), .B(n16103), .Z(n15482) );
  ANDN U25431 ( .B(n16104), .A(n16105), .Z(n16102) );
  AND U25432 ( .A(a[88]), .B(b[16]), .Z(n16101) );
  XNOR U25433 ( .A(n16106), .B(n15487), .Z(n15489) );
  XOR U25434 ( .A(n16107), .B(n16108), .Z(n15487) );
  ANDN U25435 ( .B(n16109), .A(n16110), .Z(n16107) );
  AND U25436 ( .A(a[89]), .B(b[15]), .Z(n16106) );
  XNOR U25437 ( .A(n16111), .B(n15492), .Z(n15494) );
  XOR U25438 ( .A(n16112), .B(n16113), .Z(n15492) );
  ANDN U25439 ( .B(n16114), .A(n16115), .Z(n16112) );
  AND U25440 ( .A(a[90]), .B(b[14]), .Z(n16111) );
  XNOR U25441 ( .A(n16116), .B(n15497), .Z(n15499) );
  XOR U25442 ( .A(n16117), .B(n16118), .Z(n15497) );
  ANDN U25443 ( .B(n16119), .A(n16120), .Z(n16117) );
  AND U25444 ( .A(a[91]), .B(b[13]), .Z(n16116) );
  XNOR U25445 ( .A(n16121), .B(n15502), .Z(n15504) );
  XOR U25446 ( .A(n16122), .B(n16123), .Z(n15502) );
  ANDN U25447 ( .B(n16124), .A(n16125), .Z(n16122) );
  AND U25448 ( .A(a[92]), .B(b[12]), .Z(n16121) );
  XNOR U25449 ( .A(n16126), .B(n15507), .Z(n15509) );
  XOR U25450 ( .A(n16127), .B(n16128), .Z(n15507) );
  ANDN U25451 ( .B(n16129), .A(n16130), .Z(n16127) );
  AND U25452 ( .A(a[93]), .B(b[11]), .Z(n16126) );
  XNOR U25453 ( .A(n16131), .B(n15512), .Z(n15514) );
  XOR U25454 ( .A(n16132), .B(n16133), .Z(n15512) );
  ANDN U25455 ( .B(n16134), .A(n16135), .Z(n16132) );
  AND U25456 ( .A(a[94]), .B(b[10]), .Z(n16131) );
  XNOR U25457 ( .A(n16136), .B(n15517), .Z(n15519) );
  XOR U25458 ( .A(n16137), .B(n16138), .Z(n15517) );
  ANDN U25459 ( .B(n16139), .A(n16140), .Z(n16137) );
  AND U25460 ( .A(b[9]), .B(a[95]), .Z(n16136) );
  XNOR U25461 ( .A(n16141), .B(n15522), .Z(n15524) );
  XOR U25462 ( .A(n16142), .B(n16143), .Z(n15522) );
  ANDN U25463 ( .B(n16144), .A(n16145), .Z(n16142) );
  AND U25464 ( .A(b[8]), .B(a[96]), .Z(n16141) );
  XNOR U25465 ( .A(n16146), .B(n15527), .Z(n15529) );
  XOR U25466 ( .A(n16147), .B(n16148), .Z(n15527) );
  ANDN U25467 ( .B(n16149), .A(n16150), .Z(n16147) );
  AND U25468 ( .A(b[7]), .B(a[97]), .Z(n16146) );
  XNOR U25469 ( .A(n16151), .B(n15532), .Z(n15534) );
  XOR U25470 ( .A(n16152), .B(n16153), .Z(n15532) );
  ANDN U25471 ( .B(n16154), .A(n16155), .Z(n16152) );
  AND U25472 ( .A(b[6]), .B(a[98]), .Z(n16151) );
  XNOR U25473 ( .A(n16156), .B(n15537), .Z(n15539) );
  XOR U25474 ( .A(n16157), .B(n16158), .Z(n15537) );
  ANDN U25475 ( .B(n16159), .A(n16160), .Z(n16157) );
  AND U25476 ( .A(b[5]), .B(a[99]), .Z(n16156) );
  XNOR U25477 ( .A(n16161), .B(n15542), .Z(n15544) );
  XOR U25478 ( .A(n16162), .B(n16163), .Z(n15542) );
  ANDN U25479 ( .B(n16164), .A(n16165), .Z(n16162) );
  AND U25480 ( .A(b[4]), .B(a[100]), .Z(n16161) );
  XNOR U25481 ( .A(n16166), .B(n16167), .Z(n15556) );
  NANDN U25482 ( .A(n16168), .B(n16169), .Z(n16167) );
  XNOR U25483 ( .A(n16170), .B(n15547), .Z(n15549) );
  XNOR U25484 ( .A(n16171), .B(n16172), .Z(n15547) );
  AND U25485 ( .A(n16173), .B(n16174), .Z(n16171) );
  AND U25486 ( .A(b[3]), .B(a[101]), .Z(n16170) );
  NAND U25487 ( .A(a[104]), .B(b[0]), .Z(n14940) );
  XNOR U25488 ( .A(n15562), .B(n15563), .Z(c[103]) );
  XNOR U25489 ( .A(n16168), .B(n16169), .Z(n15563) );
  XOR U25490 ( .A(n16166), .B(n16175), .Z(n16169) );
  NAND U25491 ( .A(b[1]), .B(a[102]), .Z(n16175) );
  XOR U25492 ( .A(n16174), .B(n16176), .Z(n16168) );
  XOR U25493 ( .A(n16166), .B(n16173), .Z(n16176) );
  XNOR U25494 ( .A(n16177), .B(n16172), .Z(n16173) );
  AND U25495 ( .A(b[2]), .B(a[101]), .Z(n16177) );
  NANDN U25496 ( .A(n16178), .B(n16179), .Z(n16166) );
  XOR U25497 ( .A(n16172), .B(n16164), .Z(n16180) );
  XNOR U25498 ( .A(n16163), .B(n16159), .Z(n16181) );
  XNOR U25499 ( .A(n16158), .B(n16154), .Z(n16182) );
  XNOR U25500 ( .A(n16153), .B(n16149), .Z(n16183) );
  XNOR U25501 ( .A(n16148), .B(n16144), .Z(n16184) );
  XNOR U25502 ( .A(n16143), .B(n16139), .Z(n16185) );
  XNOR U25503 ( .A(n16138), .B(n16134), .Z(n16186) );
  XNOR U25504 ( .A(n16133), .B(n16129), .Z(n16187) );
  XNOR U25505 ( .A(n16128), .B(n16124), .Z(n16188) );
  XNOR U25506 ( .A(n16123), .B(n16119), .Z(n16189) );
  XNOR U25507 ( .A(n16118), .B(n16114), .Z(n16190) );
  XNOR U25508 ( .A(n16113), .B(n16109), .Z(n16191) );
  XNOR U25509 ( .A(n16108), .B(n16104), .Z(n16192) );
  XNOR U25510 ( .A(n16103), .B(n16099), .Z(n16193) );
  XNOR U25511 ( .A(n16098), .B(n16094), .Z(n16194) );
  XNOR U25512 ( .A(n16093), .B(n16089), .Z(n16195) );
  XNOR U25513 ( .A(n16088), .B(n16084), .Z(n16196) );
  XNOR U25514 ( .A(n16083), .B(n16079), .Z(n16197) );
  XNOR U25515 ( .A(n16078), .B(n16074), .Z(n16198) );
  XNOR U25516 ( .A(n16073), .B(n16069), .Z(n16199) );
  XNOR U25517 ( .A(n16068), .B(n16064), .Z(n16200) );
  XNOR U25518 ( .A(n16063), .B(n16059), .Z(n16201) );
  XNOR U25519 ( .A(n16058), .B(n16054), .Z(n16202) );
  XNOR U25520 ( .A(n16053), .B(n16049), .Z(n16203) );
  XNOR U25521 ( .A(n16048), .B(n16044), .Z(n16204) );
  XNOR U25522 ( .A(n16043), .B(n16039), .Z(n16205) );
  XNOR U25523 ( .A(n16038), .B(n16034), .Z(n16206) );
  XNOR U25524 ( .A(n16033), .B(n16029), .Z(n16207) );
  XNOR U25525 ( .A(n16028), .B(n16024), .Z(n16208) );
  XNOR U25526 ( .A(n16023), .B(n16019), .Z(n16209) );
  XNOR U25527 ( .A(n16018), .B(n16014), .Z(n16210) );
  XNOR U25528 ( .A(n16013), .B(n16009), .Z(n16211) );
  XNOR U25529 ( .A(n16008), .B(n16004), .Z(n16212) );
  XNOR U25530 ( .A(n16003), .B(n15999), .Z(n16213) );
  XNOR U25531 ( .A(n15998), .B(n15994), .Z(n16214) );
  XNOR U25532 ( .A(n15993), .B(n15989), .Z(n16215) );
  XNOR U25533 ( .A(n15988), .B(n15984), .Z(n16216) );
  XNOR U25534 ( .A(n15983), .B(n15979), .Z(n16217) );
  XNOR U25535 ( .A(n15978), .B(n15974), .Z(n16218) );
  XNOR U25536 ( .A(n15973), .B(n15969), .Z(n16219) );
  XNOR U25537 ( .A(n15968), .B(n15964), .Z(n16220) );
  XNOR U25538 ( .A(n15963), .B(n15959), .Z(n16221) );
  XNOR U25539 ( .A(n15958), .B(n15954), .Z(n16222) );
  XNOR U25540 ( .A(n15953), .B(n15949), .Z(n16223) );
  XNOR U25541 ( .A(n15948), .B(n15944), .Z(n16224) );
  XNOR U25542 ( .A(n15943), .B(n15939), .Z(n16225) );
  XNOR U25543 ( .A(n15938), .B(n15934), .Z(n16226) );
  XNOR U25544 ( .A(n15933), .B(n15929), .Z(n16227) );
  XNOR U25545 ( .A(n15928), .B(n15924), .Z(n16228) );
  XNOR U25546 ( .A(n15923), .B(n15919), .Z(n16229) );
  XNOR U25547 ( .A(n15918), .B(n15914), .Z(n16230) );
  XNOR U25548 ( .A(n15913), .B(n15909), .Z(n16231) );
  XNOR U25549 ( .A(n15908), .B(n15904), .Z(n16232) );
  XNOR U25550 ( .A(n15903), .B(n15899), .Z(n16233) );
  XNOR U25551 ( .A(n15898), .B(n15894), .Z(n16234) );
  XNOR U25552 ( .A(n15893), .B(n15889), .Z(n16235) );
  XNOR U25553 ( .A(n15888), .B(n15884), .Z(n16236) );
  XNOR U25554 ( .A(n15883), .B(n15879), .Z(n16237) );
  XNOR U25555 ( .A(n15878), .B(n15874), .Z(n16238) );
  XNOR U25556 ( .A(n15873), .B(n15869), .Z(n16239) );
  XNOR U25557 ( .A(n15868), .B(n15864), .Z(n16240) );
  XNOR U25558 ( .A(n15863), .B(n15859), .Z(n16241) );
  XNOR U25559 ( .A(n15858), .B(n15854), .Z(n16242) );
  XNOR U25560 ( .A(n15853), .B(n15849), .Z(n16243) );
  XNOR U25561 ( .A(n15848), .B(n15844), .Z(n16244) );
  XNOR U25562 ( .A(n15843), .B(n15839), .Z(n16245) );
  XNOR U25563 ( .A(n15838), .B(n15834), .Z(n16246) );
  XNOR U25564 ( .A(n15833), .B(n15829), .Z(n16247) );
  XNOR U25565 ( .A(n15828), .B(n15824), .Z(n16248) );
  XNOR U25566 ( .A(n15823), .B(n15819), .Z(n16249) );
  XNOR U25567 ( .A(n15818), .B(n15814), .Z(n16250) );
  XNOR U25568 ( .A(n15813), .B(n15809), .Z(n16251) );
  XNOR U25569 ( .A(n15808), .B(n15804), .Z(n16252) );
  XNOR U25570 ( .A(n15803), .B(n15799), .Z(n16253) );
  XNOR U25571 ( .A(n15798), .B(n15794), .Z(n16254) );
  XNOR U25572 ( .A(n15793), .B(n15789), .Z(n16255) );
  XNOR U25573 ( .A(n15788), .B(n15784), .Z(n16256) );
  XNOR U25574 ( .A(n15783), .B(n15779), .Z(n16257) );
  XNOR U25575 ( .A(n15778), .B(n15774), .Z(n16258) );
  XNOR U25576 ( .A(n15773), .B(n15769), .Z(n16259) );
  XNOR U25577 ( .A(n15768), .B(n15764), .Z(n16260) );
  XNOR U25578 ( .A(n15763), .B(n15759), .Z(n16261) );
  XNOR U25579 ( .A(n15758), .B(n15754), .Z(n16262) );
  XNOR U25580 ( .A(n15753), .B(n15749), .Z(n16263) );
  XNOR U25581 ( .A(n15748), .B(n15744), .Z(n16264) );
  XNOR U25582 ( .A(n15743), .B(n15739), .Z(n16265) );
  XNOR U25583 ( .A(n15738), .B(n15734), .Z(n16266) );
  XNOR U25584 ( .A(n15733), .B(n15729), .Z(n16267) );
  XNOR U25585 ( .A(n15728), .B(n15724), .Z(n16268) );
  XNOR U25586 ( .A(n15723), .B(n15719), .Z(n16269) );
  XNOR U25587 ( .A(n15718), .B(n15714), .Z(n16270) );
  XNOR U25588 ( .A(n15713), .B(n15709), .Z(n16271) );
  XNOR U25589 ( .A(n15708), .B(n15704), .Z(n16272) );
  XNOR U25590 ( .A(n15703), .B(n15699), .Z(n16273) );
  XNOR U25591 ( .A(n15698), .B(n15694), .Z(n16274) );
  XNOR U25592 ( .A(n15693), .B(n15689), .Z(n16275) );
  XNOR U25593 ( .A(n15688), .B(n15684), .Z(n16276) );
  XNOR U25594 ( .A(n15683), .B(n15679), .Z(n16277) );
  XNOR U25595 ( .A(n15678), .B(n15674), .Z(n16278) );
  XNOR U25596 ( .A(n15673), .B(n15669), .Z(n16279) );
  XNOR U25597 ( .A(n16280), .B(n15668), .Z(n15669) );
  AND U25598 ( .A(a[0]), .B(b[103]), .Z(n16280) );
  XOR U25599 ( .A(n16281), .B(n15668), .Z(n15670) );
  XNOR U25600 ( .A(n16282), .B(n16283), .Z(n15668) );
  ANDN U25601 ( .B(n16284), .A(n16285), .Z(n16282) );
  AND U25602 ( .A(a[1]), .B(b[102]), .Z(n16281) );
  XNOR U25603 ( .A(n16286), .B(n15673), .Z(n15675) );
  XOR U25604 ( .A(n16287), .B(n16288), .Z(n15673) );
  ANDN U25605 ( .B(n16289), .A(n16290), .Z(n16287) );
  AND U25606 ( .A(a[2]), .B(b[101]), .Z(n16286) );
  XNOR U25607 ( .A(n16291), .B(n15678), .Z(n15680) );
  XOR U25608 ( .A(n16292), .B(n16293), .Z(n15678) );
  ANDN U25609 ( .B(n16294), .A(n16295), .Z(n16292) );
  AND U25610 ( .A(a[3]), .B(b[100]), .Z(n16291) );
  XNOR U25611 ( .A(n16296), .B(n15683), .Z(n15685) );
  XOR U25612 ( .A(n16297), .B(n16298), .Z(n15683) );
  ANDN U25613 ( .B(n16299), .A(n16300), .Z(n16297) );
  AND U25614 ( .A(a[4]), .B(b[99]), .Z(n16296) );
  XNOR U25615 ( .A(n16301), .B(n15688), .Z(n15690) );
  XOR U25616 ( .A(n16302), .B(n16303), .Z(n15688) );
  ANDN U25617 ( .B(n16304), .A(n16305), .Z(n16302) );
  AND U25618 ( .A(a[5]), .B(b[98]), .Z(n16301) );
  XNOR U25619 ( .A(n16306), .B(n15693), .Z(n15695) );
  XOR U25620 ( .A(n16307), .B(n16308), .Z(n15693) );
  ANDN U25621 ( .B(n16309), .A(n16310), .Z(n16307) );
  AND U25622 ( .A(a[6]), .B(b[97]), .Z(n16306) );
  XNOR U25623 ( .A(n16311), .B(n15698), .Z(n15700) );
  XOR U25624 ( .A(n16312), .B(n16313), .Z(n15698) );
  ANDN U25625 ( .B(n16314), .A(n16315), .Z(n16312) );
  AND U25626 ( .A(a[7]), .B(b[96]), .Z(n16311) );
  XNOR U25627 ( .A(n16316), .B(n15703), .Z(n15705) );
  XOR U25628 ( .A(n16317), .B(n16318), .Z(n15703) );
  ANDN U25629 ( .B(n16319), .A(n16320), .Z(n16317) );
  AND U25630 ( .A(a[8]), .B(b[95]), .Z(n16316) );
  XNOR U25631 ( .A(n16321), .B(n15708), .Z(n15710) );
  XOR U25632 ( .A(n16322), .B(n16323), .Z(n15708) );
  ANDN U25633 ( .B(n16324), .A(n16325), .Z(n16322) );
  AND U25634 ( .A(a[9]), .B(b[94]), .Z(n16321) );
  XNOR U25635 ( .A(n16326), .B(n15713), .Z(n15715) );
  XOR U25636 ( .A(n16327), .B(n16328), .Z(n15713) );
  ANDN U25637 ( .B(n16329), .A(n16330), .Z(n16327) );
  AND U25638 ( .A(a[10]), .B(b[93]), .Z(n16326) );
  XNOR U25639 ( .A(n16331), .B(n15718), .Z(n15720) );
  XOR U25640 ( .A(n16332), .B(n16333), .Z(n15718) );
  ANDN U25641 ( .B(n16334), .A(n16335), .Z(n16332) );
  AND U25642 ( .A(a[11]), .B(b[92]), .Z(n16331) );
  XNOR U25643 ( .A(n16336), .B(n15723), .Z(n15725) );
  XOR U25644 ( .A(n16337), .B(n16338), .Z(n15723) );
  ANDN U25645 ( .B(n16339), .A(n16340), .Z(n16337) );
  AND U25646 ( .A(a[12]), .B(b[91]), .Z(n16336) );
  XNOR U25647 ( .A(n16341), .B(n15728), .Z(n15730) );
  XOR U25648 ( .A(n16342), .B(n16343), .Z(n15728) );
  ANDN U25649 ( .B(n16344), .A(n16345), .Z(n16342) );
  AND U25650 ( .A(a[13]), .B(b[90]), .Z(n16341) );
  XNOR U25651 ( .A(n16346), .B(n15733), .Z(n15735) );
  XOR U25652 ( .A(n16347), .B(n16348), .Z(n15733) );
  ANDN U25653 ( .B(n16349), .A(n16350), .Z(n16347) );
  AND U25654 ( .A(a[14]), .B(b[89]), .Z(n16346) );
  XNOR U25655 ( .A(n16351), .B(n15738), .Z(n15740) );
  XOR U25656 ( .A(n16352), .B(n16353), .Z(n15738) );
  ANDN U25657 ( .B(n16354), .A(n16355), .Z(n16352) );
  AND U25658 ( .A(a[15]), .B(b[88]), .Z(n16351) );
  XNOR U25659 ( .A(n16356), .B(n15743), .Z(n15745) );
  XOR U25660 ( .A(n16357), .B(n16358), .Z(n15743) );
  ANDN U25661 ( .B(n16359), .A(n16360), .Z(n16357) );
  AND U25662 ( .A(a[16]), .B(b[87]), .Z(n16356) );
  XNOR U25663 ( .A(n16361), .B(n15748), .Z(n15750) );
  XOR U25664 ( .A(n16362), .B(n16363), .Z(n15748) );
  ANDN U25665 ( .B(n16364), .A(n16365), .Z(n16362) );
  AND U25666 ( .A(a[17]), .B(b[86]), .Z(n16361) );
  XNOR U25667 ( .A(n16366), .B(n15753), .Z(n15755) );
  XOR U25668 ( .A(n16367), .B(n16368), .Z(n15753) );
  ANDN U25669 ( .B(n16369), .A(n16370), .Z(n16367) );
  AND U25670 ( .A(a[18]), .B(b[85]), .Z(n16366) );
  XNOR U25671 ( .A(n16371), .B(n15758), .Z(n15760) );
  XOR U25672 ( .A(n16372), .B(n16373), .Z(n15758) );
  ANDN U25673 ( .B(n16374), .A(n16375), .Z(n16372) );
  AND U25674 ( .A(a[19]), .B(b[84]), .Z(n16371) );
  XNOR U25675 ( .A(n16376), .B(n15763), .Z(n15765) );
  XOR U25676 ( .A(n16377), .B(n16378), .Z(n15763) );
  ANDN U25677 ( .B(n16379), .A(n16380), .Z(n16377) );
  AND U25678 ( .A(a[20]), .B(b[83]), .Z(n16376) );
  XNOR U25679 ( .A(n16381), .B(n15768), .Z(n15770) );
  XOR U25680 ( .A(n16382), .B(n16383), .Z(n15768) );
  ANDN U25681 ( .B(n16384), .A(n16385), .Z(n16382) );
  AND U25682 ( .A(a[21]), .B(b[82]), .Z(n16381) );
  XNOR U25683 ( .A(n16386), .B(n15773), .Z(n15775) );
  XOR U25684 ( .A(n16387), .B(n16388), .Z(n15773) );
  ANDN U25685 ( .B(n16389), .A(n16390), .Z(n16387) );
  AND U25686 ( .A(a[22]), .B(b[81]), .Z(n16386) );
  XNOR U25687 ( .A(n16391), .B(n15778), .Z(n15780) );
  XOR U25688 ( .A(n16392), .B(n16393), .Z(n15778) );
  ANDN U25689 ( .B(n16394), .A(n16395), .Z(n16392) );
  AND U25690 ( .A(a[23]), .B(b[80]), .Z(n16391) );
  XNOR U25691 ( .A(n16396), .B(n15783), .Z(n15785) );
  XOR U25692 ( .A(n16397), .B(n16398), .Z(n15783) );
  ANDN U25693 ( .B(n16399), .A(n16400), .Z(n16397) );
  AND U25694 ( .A(a[24]), .B(b[79]), .Z(n16396) );
  XNOR U25695 ( .A(n16401), .B(n15788), .Z(n15790) );
  XOR U25696 ( .A(n16402), .B(n16403), .Z(n15788) );
  ANDN U25697 ( .B(n16404), .A(n16405), .Z(n16402) );
  AND U25698 ( .A(a[25]), .B(b[78]), .Z(n16401) );
  XNOR U25699 ( .A(n16406), .B(n15793), .Z(n15795) );
  XOR U25700 ( .A(n16407), .B(n16408), .Z(n15793) );
  ANDN U25701 ( .B(n16409), .A(n16410), .Z(n16407) );
  AND U25702 ( .A(a[26]), .B(b[77]), .Z(n16406) );
  XNOR U25703 ( .A(n16411), .B(n15798), .Z(n15800) );
  XOR U25704 ( .A(n16412), .B(n16413), .Z(n15798) );
  ANDN U25705 ( .B(n16414), .A(n16415), .Z(n16412) );
  AND U25706 ( .A(a[27]), .B(b[76]), .Z(n16411) );
  XNOR U25707 ( .A(n16416), .B(n15803), .Z(n15805) );
  XOR U25708 ( .A(n16417), .B(n16418), .Z(n15803) );
  ANDN U25709 ( .B(n16419), .A(n16420), .Z(n16417) );
  AND U25710 ( .A(a[28]), .B(b[75]), .Z(n16416) );
  XNOR U25711 ( .A(n16421), .B(n15808), .Z(n15810) );
  XOR U25712 ( .A(n16422), .B(n16423), .Z(n15808) );
  ANDN U25713 ( .B(n16424), .A(n16425), .Z(n16422) );
  AND U25714 ( .A(a[29]), .B(b[74]), .Z(n16421) );
  XNOR U25715 ( .A(n16426), .B(n15813), .Z(n15815) );
  XOR U25716 ( .A(n16427), .B(n16428), .Z(n15813) );
  ANDN U25717 ( .B(n16429), .A(n16430), .Z(n16427) );
  AND U25718 ( .A(a[30]), .B(b[73]), .Z(n16426) );
  XNOR U25719 ( .A(n16431), .B(n15818), .Z(n15820) );
  XOR U25720 ( .A(n16432), .B(n16433), .Z(n15818) );
  ANDN U25721 ( .B(n16434), .A(n16435), .Z(n16432) );
  AND U25722 ( .A(a[31]), .B(b[72]), .Z(n16431) );
  XNOR U25723 ( .A(n16436), .B(n15823), .Z(n15825) );
  XOR U25724 ( .A(n16437), .B(n16438), .Z(n15823) );
  ANDN U25725 ( .B(n16439), .A(n16440), .Z(n16437) );
  AND U25726 ( .A(a[32]), .B(b[71]), .Z(n16436) );
  XNOR U25727 ( .A(n16441), .B(n15828), .Z(n15830) );
  XOR U25728 ( .A(n16442), .B(n16443), .Z(n15828) );
  ANDN U25729 ( .B(n16444), .A(n16445), .Z(n16442) );
  AND U25730 ( .A(a[33]), .B(b[70]), .Z(n16441) );
  XNOR U25731 ( .A(n16446), .B(n15833), .Z(n15835) );
  XOR U25732 ( .A(n16447), .B(n16448), .Z(n15833) );
  ANDN U25733 ( .B(n16449), .A(n16450), .Z(n16447) );
  AND U25734 ( .A(a[34]), .B(b[69]), .Z(n16446) );
  XNOR U25735 ( .A(n16451), .B(n15838), .Z(n15840) );
  XOR U25736 ( .A(n16452), .B(n16453), .Z(n15838) );
  ANDN U25737 ( .B(n16454), .A(n16455), .Z(n16452) );
  AND U25738 ( .A(a[35]), .B(b[68]), .Z(n16451) );
  XNOR U25739 ( .A(n16456), .B(n15843), .Z(n15845) );
  XOR U25740 ( .A(n16457), .B(n16458), .Z(n15843) );
  ANDN U25741 ( .B(n16459), .A(n16460), .Z(n16457) );
  AND U25742 ( .A(a[36]), .B(b[67]), .Z(n16456) );
  XNOR U25743 ( .A(n16461), .B(n15848), .Z(n15850) );
  XOR U25744 ( .A(n16462), .B(n16463), .Z(n15848) );
  ANDN U25745 ( .B(n16464), .A(n16465), .Z(n16462) );
  AND U25746 ( .A(a[37]), .B(b[66]), .Z(n16461) );
  XNOR U25747 ( .A(n16466), .B(n15853), .Z(n15855) );
  XOR U25748 ( .A(n16467), .B(n16468), .Z(n15853) );
  ANDN U25749 ( .B(n16469), .A(n16470), .Z(n16467) );
  AND U25750 ( .A(a[38]), .B(b[65]), .Z(n16466) );
  XNOR U25751 ( .A(n16471), .B(n15858), .Z(n15860) );
  XOR U25752 ( .A(n16472), .B(n16473), .Z(n15858) );
  ANDN U25753 ( .B(n16474), .A(n16475), .Z(n16472) );
  AND U25754 ( .A(a[39]), .B(b[64]), .Z(n16471) );
  XNOR U25755 ( .A(n16476), .B(n15863), .Z(n15865) );
  XOR U25756 ( .A(n16477), .B(n16478), .Z(n15863) );
  ANDN U25757 ( .B(n16479), .A(n16480), .Z(n16477) );
  AND U25758 ( .A(a[40]), .B(b[63]), .Z(n16476) );
  XNOR U25759 ( .A(n16481), .B(n15868), .Z(n15870) );
  XOR U25760 ( .A(n16482), .B(n16483), .Z(n15868) );
  ANDN U25761 ( .B(n16484), .A(n16485), .Z(n16482) );
  AND U25762 ( .A(a[41]), .B(b[62]), .Z(n16481) );
  XNOR U25763 ( .A(n16486), .B(n15873), .Z(n15875) );
  XOR U25764 ( .A(n16487), .B(n16488), .Z(n15873) );
  ANDN U25765 ( .B(n16489), .A(n16490), .Z(n16487) );
  AND U25766 ( .A(a[42]), .B(b[61]), .Z(n16486) );
  XNOR U25767 ( .A(n16491), .B(n15878), .Z(n15880) );
  XOR U25768 ( .A(n16492), .B(n16493), .Z(n15878) );
  ANDN U25769 ( .B(n16494), .A(n16495), .Z(n16492) );
  AND U25770 ( .A(a[43]), .B(b[60]), .Z(n16491) );
  XNOR U25771 ( .A(n16496), .B(n15883), .Z(n15885) );
  XOR U25772 ( .A(n16497), .B(n16498), .Z(n15883) );
  ANDN U25773 ( .B(n16499), .A(n16500), .Z(n16497) );
  AND U25774 ( .A(a[44]), .B(b[59]), .Z(n16496) );
  XNOR U25775 ( .A(n16501), .B(n15888), .Z(n15890) );
  XOR U25776 ( .A(n16502), .B(n16503), .Z(n15888) );
  ANDN U25777 ( .B(n16504), .A(n16505), .Z(n16502) );
  AND U25778 ( .A(a[45]), .B(b[58]), .Z(n16501) );
  XNOR U25779 ( .A(n16506), .B(n15893), .Z(n15895) );
  XOR U25780 ( .A(n16507), .B(n16508), .Z(n15893) );
  ANDN U25781 ( .B(n16509), .A(n16510), .Z(n16507) );
  AND U25782 ( .A(a[46]), .B(b[57]), .Z(n16506) );
  XNOR U25783 ( .A(n16511), .B(n15898), .Z(n15900) );
  XOR U25784 ( .A(n16512), .B(n16513), .Z(n15898) );
  ANDN U25785 ( .B(n16514), .A(n16515), .Z(n16512) );
  AND U25786 ( .A(a[47]), .B(b[56]), .Z(n16511) );
  XNOR U25787 ( .A(n16516), .B(n15903), .Z(n15905) );
  XOR U25788 ( .A(n16517), .B(n16518), .Z(n15903) );
  ANDN U25789 ( .B(n16519), .A(n16520), .Z(n16517) );
  AND U25790 ( .A(a[48]), .B(b[55]), .Z(n16516) );
  XNOR U25791 ( .A(n16521), .B(n15908), .Z(n15910) );
  XOR U25792 ( .A(n16522), .B(n16523), .Z(n15908) );
  ANDN U25793 ( .B(n16524), .A(n16525), .Z(n16522) );
  AND U25794 ( .A(a[49]), .B(b[54]), .Z(n16521) );
  XNOR U25795 ( .A(n16526), .B(n15913), .Z(n15915) );
  XOR U25796 ( .A(n16527), .B(n16528), .Z(n15913) );
  ANDN U25797 ( .B(n16529), .A(n16530), .Z(n16527) );
  AND U25798 ( .A(a[50]), .B(b[53]), .Z(n16526) );
  XNOR U25799 ( .A(n16531), .B(n15918), .Z(n15920) );
  XOR U25800 ( .A(n16532), .B(n16533), .Z(n15918) );
  ANDN U25801 ( .B(n16534), .A(n16535), .Z(n16532) );
  AND U25802 ( .A(a[51]), .B(b[52]), .Z(n16531) );
  XNOR U25803 ( .A(n16536), .B(n15923), .Z(n15925) );
  XOR U25804 ( .A(n16537), .B(n16538), .Z(n15923) );
  ANDN U25805 ( .B(n16539), .A(n16540), .Z(n16537) );
  AND U25806 ( .A(a[52]), .B(b[51]), .Z(n16536) );
  XNOR U25807 ( .A(n16541), .B(n15928), .Z(n15930) );
  XOR U25808 ( .A(n16542), .B(n16543), .Z(n15928) );
  ANDN U25809 ( .B(n16544), .A(n16545), .Z(n16542) );
  AND U25810 ( .A(a[53]), .B(b[50]), .Z(n16541) );
  XNOR U25811 ( .A(n16546), .B(n15933), .Z(n15935) );
  XOR U25812 ( .A(n16547), .B(n16548), .Z(n15933) );
  ANDN U25813 ( .B(n16549), .A(n16550), .Z(n16547) );
  AND U25814 ( .A(a[54]), .B(b[49]), .Z(n16546) );
  XNOR U25815 ( .A(n16551), .B(n15938), .Z(n15940) );
  XOR U25816 ( .A(n16552), .B(n16553), .Z(n15938) );
  ANDN U25817 ( .B(n16554), .A(n16555), .Z(n16552) );
  AND U25818 ( .A(a[55]), .B(b[48]), .Z(n16551) );
  XNOR U25819 ( .A(n16556), .B(n15943), .Z(n15945) );
  XOR U25820 ( .A(n16557), .B(n16558), .Z(n15943) );
  ANDN U25821 ( .B(n16559), .A(n16560), .Z(n16557) );
  AND U25822 ( .A(a[56]), .B(b[47]), .Z(n16556) );
  XNOR U25823 ( .A(n16561), .B(n15948), .Z(n15950) );
  XOR U25824 ( .A(n16562), .B(n16563), .Z(n15948) );
  ANDN U25825 ( .B(n16564), .A(n16565), .Z(n16562) );
  AND U25826 ( .A(a[57]), .B(b[46]), .Z(n16561) );
  XNOR U25827 ( .A(n16566), .B(n15953), .Z(n15955) );
  XOR U25828 ( .A(n16567), .B(n16568), .Z(n15953) );
  ANDN U25829 ( .B(n16569), .A(n16570), .Z(n16567) );
  AND U25830 ( .A(a[58]), .B(b[45]), .Z(n16566) );
  XNOR U25831 ( .A(n16571), .B(n15958), .Z(n15960) );
  XOR U25832 ( .A(n16572), .B(n16573), .Z(n15958) );
  ANDN U25833 ( .B(n16574), .A(n16575), .Z(n16572) );
  AND U25834 ( .A(a[59]), .B(b[44]), .Z(n16571) );
  XNOR U25835 ( .A(n16576), .B(n15963), .Z(n15965) );
  XOR U25836 ( .A(n16577), .B(n16578), .Z(n15963) );
  ANDN U25837 ( .B(n16579), .A(n16580), .Z(n16577) );
  AND U25838 ( .A(a[60]), .B(b[43]), .Z(n16576) );
  XNOR U25839 ( .A(n16581), .B(n15968), .Z(n15970) );
  XOR U25840 ( .A(n16582), .B(n16583), .Z(n15968) );
  ANDN U25841 ( .B(n16584), .A(n16585), .Z(n16582) );
  AND U25842 ( .A(a[61]), .B(b[42]), .Z(n16581) );
  XNOR U25843 ( .A(n16586), .B(n15973), .Z(n15975) );
  XOR U25844 ( .A(n16587), .B(n16588), .Z(n15973) );
  ANDN U25845 ( .B(n16589), .A(n16590), .Z(n16587) );
  AND U25846 ( .A(a[62]), .B(b[41]), .Z(n16586) );
  XNOR U25847 ( .A(n16591), .B(n15978), .Z(n15980) );
  XOR U25848 ( .A(n16592), .B(n16593), .Z(n15978) );
  ANDN U25849 ( .B(n16594), .A(n16595), .Z(n16592) );
  AND U25850 ( .A(a[63]), .B(b[40]), .Z(n16591) );
  XNOR U25851 ( .A(n16596), .B(n15983), .Z(n15985) );
  XOR U25852 ( .A(n16597), .B(n16598), .Z(n15983) );
  ANDN U25853 ( .B(n16599), .A(n16600), .Z(n16597) );
  AND U25854 ( .A(a[64]), .B(b[39]), .Z(n16596) );
  XNOR U25855 ( .A(n16601), .B(n15988), .Z(n15990) );
  XOR U25856 ( .A(n16602), .B(n16603), .Z(n15988) );
  ANDN U25857 ( .B(n16604), .A(n16605), .Z(n16602) );
  AND U25858 ( .A(a[65]), .B(b[38]), .Z(n16601) );
  XNOR U25859 ( .A(n16606), .B(n15993), .Z(n15995) );
  XOR U25860 ( .A(n16607), .B(n16608), .Z(n15993) );
  ANDN U25861 ( .B(n16609), .A(n16610), .Z(n16607) );
  AND U25862 ( .A(a[66]), .B(b[37]), .Z(n16606) );
  XNOR U25863 ( .A(n16611), .B(n15998), .Z(n16000) );
  XOR U25864 ( .A(n16612), .B(n16613), .Z(n15998) );
  ANDN U25865 ( .B(n16614), .A(n16615), .Z(n16612) );
  AND U25866 ( .A(a[67]), .B(b[36]), .Z(n16611) );
  XNOR U25867 ( .A(n16616), .B(n16003), .Z(n16005) );
  XOR U25868 ( .A(n16617), .B(n16618), .Z(n16003) );
  ANDN U25869 ( .B(n16619), .A(n16620), .Z(n16617) );
  AND U25870 ( .A(a[68]), .B(b[35]), .Z(n16616) );
  XNOR U25871 ( .A(n16621), .B(n16008), .Z(n16010) );
  XOR U25872 ( .A(n16622), .B(n16623), .Z(n16008) );
  ANDN U25873 ( .B(n16624), .A(n16625), .Z(n16622) );
  AND U25874 ( .A(a[69]), .B(b[34]), .Z(n16621) );
  XNOR U25875 ( .A(n16626), .B(n16013), .Z(n16015) );
  XOR U25876 ( .A(n16627), .B(n16628), .Z(n16013) );
  ANDN U25877 ( .B(n16629), .A(n16630), .Z(n16627) );
  AND U25878 ( .A(a[70]), .B(b[33]), .Z(n16626) );
  XNOR U25879 ( .A(n16631), .B(n16018), .Z(n16020) );
  XOR U25880 ( .A(n16632), .B(n16633), .Z(n16018) );
  ANDN U25881 ( .B(n16634), .A(n16635), .Z(n16632) );
  AND U25882 ( .A(a[71]), .B(b[32]), .Z(n16631) );
  XNOR U25883 ( .A(n16636), .B(n16023), .Z(n16025) );
  XOR U25884 ( .A(n16637), .B(n16638), .Z(n16023) );
  ANDN U25885 ( .B(n16639), .A(n16640), .Z(n16637) );
  AND U25886 ( .A(a[72]), .B(b[31]), .Z(n16636) );
  XNOR U25887 ( .A(n16641), .B(n16028), .Z(n16030) );
  XOR U25888 ( .A(n16642), .B(n16643), .Z(n16028) );
  ANDN U25889 ( .B(n16644), .A(n16645), .Z(n16642) );
  AND U25890 ( .A(a[73]), .B(b[30]), .Z(n16641) );
  XNOR U25891 ( .A(n16646), .B(n16033), .Z(n16035) );
  XOR U25892 ( .A(n16647), .B(n16648), .Z(n16033) );
  ANDN U25893 ( .B(n16649), .A(n16650), .Z(n16647) );
  AND U25894 ( .A(a[74]), .B(b[29]), .Z(n16646) );
  XNOR U25895 ( .A(n16651), .B(n16038), .Z(n16040) );
  XOR U25896 ( .A(n16652), .B(n16653), .Z(n16038) );
  ANDN U25897 ( .B(n16654), .A(n16655), .Z(n16652) );
  AND U25898 ( .A(a[75]), .B(b[28]), .Z(n16651) );
  XNOR U25899 ( .A(n16656), .B(n16043), .Z(n16045) );
  XOR U25900 ( .A(n16657), .B(n16658), .Z(n16043) );
  ANDN U25901 ( .B(n16659), .A(n16660), .Z(n16657) );
  AND U25902 ( .A(a[76]), .B(b[27]), .Z(n16656) );
  XNOR U25903 ( .A(n16661), .B(n16048), .Z(n16050) );
  XOR U25904 ( .A(n16662), .B(n16663), .Z(n16048) );
  ANDN U25905 ( .B(n16664), .A(n16665), .Z(n16662) );
  AND U25906 ( .A(a[77]), .B(b[26]), .Z(n16661) );
  XNOR U25907 ( .A(n16666), .B(n16053), .Z(n16055) );
  XOR U25908 ( .A(n16667), .B(n16668), .Z(n16053) );
  ANDN U25909 ( .B(n16669), .A(n16670), .Z(n16667) );
  AND U25910 ( .A(a[78]), .B(b[25]), .Z(n16666) );
  XNOR U25911 ( .A(n16671), .B(n16058), .Z(n16060) );
  XOR U25912 ( .A(n16672), .B(n16673), .Z(n16058) );
  ANDN U25913 ( .B(n16674), .A(n16675), .Z(n16672) );
  AND U25914 ( .A(a[79]), .B(b[24]), .Z(n16671) );
  XNOR U25915 ( .A(n16676), .B(n16063), .Z(n16065) );
  XOR U25916 ( .A(n16677), .B(n16678), .Z(n16063) );
  ANDN U25917 ( .B(n16679), .A(n16680), .Z(n16677) );
  AND U25918 ( .A(a[80]), .B(b[23]), .Z(n16676) );
  XNOR U25919 ( .A(n16681), .B(n16068), .Z(n16070) );
  XOR U25920 ( .A(n16682), .B(n16683), .Z(n16068) );
  ANDN U25921 ( .B(n16684), .A(n16685), .Z(n16682) );
  AND U25922 ( .A(a[81]), .B(b[22]), .Z(n16681) );
  XNOR U25923 ( .A(n16686), .B(n16073), .Z(n16075) );
  XOR U25924 ( .A(n16687), .B(n16688), .Z(n16073) );
  ANDN U25925 ( .B(n16689), .A(n16690), .Z(n16687) );
  AND U25926 ( .A(a[82]), .B(b[21]), .Z(n16686) );
  XNOR U25927 ( .A(n16691), .B(n16078), .Z(n16080) );
  XOR U25928 ( .A(n16692), .B(n16693), .Z(n16078) );
  ANDN U25929 ( .B(n16694), .A(n16695), .Z(n16692) );
  AND U25930 ( .A(a[83]), .B(b[20]), .Z(n16691) );
  XNOR U25931 ( .A(n16696), .B(n16083), .Z(n16085) );
  XOR U25932 ( .A(n16697), .B(n16698), .Z(n16083) );
  ANDN U25933 ( .B(n16699), .A(n16700), .Z(n16697) );
  AND U25934 ( .A(a[84]), .B(b[19]), .Z(n16696) );
  XNOR U25935 ( .A(n16701), .B(n16088), .Z(n16090) );
  XOR U25936 ( .A(n16702), .B(n16703), .Z(n16088) );
  ANDN U25937 ( .B(n16704), .A(n16705), .Z(n16702) );
  AND U25938 ( .A(a[85]), .B(b[18]), .Z(n16701) );
  XNOR U25939 ( .A(n16706), .B(n16093), .Z(n16095) );
  XOR U25940 ( .A(n16707), .B(n16708), .Z(n16093) );
  ANDN U25941 ( .B(n16709), .A(n16710), .Z(n16707) );
  AND U25942 ( .A(a[86]), .B(b[17]), .Z(n16706) );
  XNOR U25943 ( .A(n16711), .B(n16098), .Z(n16100) );
  XOR U25944 ( .A(n16712), .B(n16713), .Z(n16098) );
  ANDN U25945 ( .B(n16714), .A(n16715), .Z(n16712) );
  AND U25946 ( .A(a[87]), .B(b[16]), .Z(n16711) );
  XNOR U25947 ( .A(n16716), .B(n16103), .Z(n16105) );
  XOR U25948 ( .A(n16717), .B(n16718), .Z(n16103) );
  ANDN U25949 ( .B(n16719), .A(n16720), .Z(n16717) );
  AND U25950 ( .A(a[88]), .B(b[15]), .Z(n16716) );
  XNOR U25951 ( .A(n16721), .B(n16108), .Z(n16110) );
  XOR U25952 ( .A(n16722), .B(n16723), .Z(n16108) );
  ANDN U25953 ( .B(n16724), .A(n16725), .Z(n16722) );
  AND U25954 ( .A(a[89]), .B(b[14]), .Z(n16721) );
  XNOR U25955 ( .A(n16726), .B(n16113), .Z(n16115) );
  XOR U25956 ( .A(n16727), .B(n16728), .Z(n16113) );
  ANDN U25957 ( .B(n16729), .A(n16730), .Z(n16727) );
  AND U25958 ( .A(a[90]), .B(b[13]), .Z(n16726) );
  XNOR U25959 ( .A(n16731), .B(n16118), .Z(n16120) );
  XOR U25960 ( .A(n16732), .B(n16733), .Z(n16118) );
  ANDN U25961 ( .B(n16734), .A(n16735), .Z(n16732) );
  AND U25962 ( .A(a[91]), .B(b[12]), .Z(n16731) );
  XNOR U25963 ( .A(n16736), .B(n16123), .Z(n16125) );
  XOR U25964 ( .A(n16737), .B(n16738), .Z(n16123) );
  ANDN U25965 ( .B(n16739), .A(n16740), .Z(n16737) );
  AND U25966 ( .A(a[92]), .B(b[11]), .Z(n16736) );
  XNOR U25967 ( .A(n16741), .B(n16128), .Z(n16130) );
  XOR U25968 ( .A(n16742), .B(n16743), .Z(n16128) );
  ANDN U25969 ( .B(n16744), .A(n16745), .Z(n16742) );
  AND U25970 ( .A(a[93]), .B(b[10]), .Z(n16741) );
  XNOR U25971 ( .A(n16746), .B(n16133), .Z(n16135) );
  XOR U25972 ( .A(n16747), .B(n16748), .Z(n16133) );
  ANDN U25973 ( .B(n16749), .A(n16750), .Z(n16747) );
  AND U25974 ( .A(b[9]), .B(a[94]), .Z(n16746) );
  XNOR U25975 ( .A(n16751), .B(n16138), .Z(n16140) );
  XOR U25976 ( .A(n16752), .B(n16753), .Z(n16138) );
  ANDN U25977 ( .B(n16754), .A(n16755), .Z(n16752) );
  AND U25978 ( .A(b[8]), .B(a[95]), .Z(n16751) );
  XNOR U25979 ( .A(n16756), .B(n16143), .Z(n16145) );
  XOR U25980 ( .A(n16757), .B(n16758), .Z(n16143) );
  ANDN U25981 ( .B(n16759), .A(n16760), .Z(n16757) );
  AND U25982 ( .A(b[7]), .B(a[96]), .Z(n16756) );
  XNOR U25983 ( .A(n16761), .B(n16148), .Z(n16150) );
  XOR U25984 ( .A(n16762), .B(n16763), .Z(n16148) );
  ANDN U25985 ( .B(n16764), .A(n16765), .Z(n16762) );
  AND U25986 ( .A(b[6]), .B(a[97]), .Z(n16761) );
  XNOR U25987 ( .A(n16766), .B(n16153), .Z(n16155) );
  XOR U25988 ( .A(n16767), .B(n16768), .Z(n16153) );
  ANDN U25989 ( .B(n16769), .A(n16770), .Z(n16767) );
  AND U25990 ( .A(b[5]), .B(a[98]), .Z(n16766) );
  XNOR U25991 ( .A(n16771), .B(n16158), .Z(n16160) );
  XOR U25992 ( .A(n16772), .B(n16773), .Z(n16158) );
  ANDN U25993 ( .B(n16774), .A(n16775), .Z(n16772) );
  AND U25994 ( .A(b[4]), .B(a[99]), .Z(n16771) );
  XNOR U25995 ( .A(n16776), .B(n16777), .Z(n16172) );
  NANDN U25996 ( .A(n16778), .B(n16779), .Z(n16777) );
  XNOR U25997 ( .A(n16780), .B(n16163), .Z(n16165) );
  XNOR U25998 ( .A(n16781), .B(n16782), .Z(n16163) );
  AND U25999 ( .A(n16783), .B(n16784), .Z(n16781) );
  AND U26000 ( .A(b[3]), .B(a[100]), .Z(n16780) );
  NAND U26001 ( .A(a[103]), .B(b[0]), .Z(n15562) );
  XNOR U26002 ( .A(n16178), .B(n16179), .Z(c[102]) );
  XNOR U26003 ( .A(n16778), .B(n16779), .Z(n16179) );
  XOR U26004 ( .A(n16776), .B(n16785), .Z(n16779) );
  NAND U26005 ( .A(b[1]), .B(a[101]), .Z(n16785) );
  XOR U26006 ( .A(n16784), .B(n16786), .Z(n16778) );
  XOR U26007 ( .A(n16776), .B(n16783), .Z(n16786) );
  XNOR U26008 ( .A(n16787), .B(n16782), .Z(n16783) );
  AND U26009 ( .A(b[2]), .B(a[100]), .Z(n16787) );
  NANDN U26010 ( .A(n16788), .B(n16789), .Z(n16776) );
  XOR U26011 ( .A(n16782), .B(n16774), .Z(n16790) );
  XNOR U26012 ( .A(n16773), .B(n16769), .Z(n16791) );
  XNOR U26013 ( .A(n16768), .B(n16764), .Z(n16792) );
  XNOR U26014 ( .A(n16763), .B(n16759), .Z(n16793) );
  XNOR U26015 ( .A(n16758), .B(n16754), .Z(n16794) );
  XNOR U26016 ( .A(n16753), .B(n16749), .Z(n16795) );
  XNOR U26017 ( .A(n16748), .B(n16744), .Z(n16796) );
  XNOR U26018 ( .A(n16743), .B(n16739), .Z(n16797) );
  XNOR U26019 ( .A(n16738), .B(n16734), .Z(n16798) );
  XNOR U26020 ( .A(n16733), .B(n16729), .Z(n16799) );
  XNOR U26021 ( .A(n16728), .B(n16724), .Z(n16800) );
  XNOR U26022 ( .A(n16723), .B(n16719), .Z(n16801) );
  XNOR U26023 ( .A(n16718), .B(n16714), .Z(n16802) );
  XNOR U26024 ( .A(n16713), .B(n16709), .Z(n16803) );
  XNOR U26025 ( .A(n16708), .B(n16704), .Z(n16804) );
  XNOR U26026 ( .A(n16703), .B(n16699), .Z(n16805) );
  XNOR U26027 ( .A(n16698), .B(n16694), .Z(n16806) );
  XNOR U26028 ( .A(n16693), .B(n16689), .Z(n16807) );
  XNOR U26029 ( .A(n16688), .B(n16684), .Z(n16808) );
  XNOR U26030 ( .A(n16683), .B(n16679), .Z(n16809) );
  XNOR U26031 ( .A(n16678), .B(n16674), .Z(n16810) );
  XNOR U26032 ( .A(n16673), .B(n16669), .Z(n16811) );
  XNOR U26033 ( .A(n16668), .B(n16664), .Z(n16812) );
  XNOR U26034 ( .A(n16663), .B(n16659), .Z(n16813) );
  XNOR U26035 ( .A(n16658), .B(n16654), .Z(n16814) );
  XNOR U26036 ( .A(n16653), .B(n16649), .Z(n16815) );
  XNOR U26037 ( .A(n16648), .B(n16644), .Z(n16816) );
  XNOR U26038 ( .A(n16643), .B(n16639), .Z(n16817) );
  XNOR U26039 ( .A(n16638), .B(n16634), .Z(n16818) );
  XNOR U26040 ( .A(n16633), .B(n16629), .Z(n16819) );
  XNOR U26041 ( .A(n16628), .B(n16624), .Z(n16820) );
  XNOR U26042 ( .A(n16623), .B(n16619), .Z(n16821) );
  XNOR U26043 ( .A(n16618), .B(n16614), .Z(n16822) );
  XNOR U26044 ( .A(n16613), .B(n16609), .Z(n16823) );
  XNOR U26045 ( .A(n16608), .B(n16604), .Z(n16824) );
  XNOR U26046 ( .A(n16603), .B(n16599), .Z(n16825) );
  XNOR U26047 ( .A(n16598), .B(n16594), .Z(n16826) );
  XNOR U26048 ( .A(n16593), .B(n16589), .Z(n16827) );
  XNOR U26049 ( .A(n16588), .B(n16584), .Z(n16828) );
  XNOR U26050 ( .A(n16583), .B(n16579), .Z(n16829) );
  XNOR U26051 ( .A(n16578), .B(n16574), .Z(n16830) );
  XNOR U26052 ( .A(n16573), .B(n16569), .Z(n16831) );
  XNOR U26053 ( .A(n16568), .B(n16564), .Z(n16832) );
  XNOR U26054 ( .A(n16563), .B(n16559), .Z(n16833) );
  XNOR U26055 ( .A(n16558), .B(n16554), .Z(n16834) );
  XNOR U26056 ( .A(n16553), .B(n16549), .Z(n16835) );
  XNOR U26057 ( .A(n16548), .B(n16544), .Z(n16836) );
  XNOR U26058 ( .A(n16543), .B(n16539), .Z(n16837) );
  XNOR U26059 ( .A(n16538), .B(n16534), .Z(n16838) );
  XNOR U26060 ( .A(n16533), .B(n16529), .Z(n16839) );
  XNOR U26061 ( .A(n16528), .B(n16524), .Z(n16840) );
  XNOR U26062 ( .A(n16523), .B(n16519), .Z(n16841) );
  XNOR U26063 ( .A(n16518), .B(n16514), .Z(n16842) );
  XNOR U26064 ( .A(n16513), .B(n16509), .Z(n16843) );
  XNOR U26065 ( .A(n16508), .B(n16504), .Z(n16844) );
  XNOR U26066 ( .A(n16503), .B(n16499), .Z(n16845) );
  XNOR U26067 ( .A(n16498), .B(n16494), .Z(n16846) );
  XNOR U26068 ( .A(n16493), .B(n16489), .Z(n16847) );
  XNOR U26069 ( .A(n16488), .B(n16484), .Z(n16848) );
  XNOR U26070 ( .A(n16483), .B(n16479), .Z(n16849) );
  XNOR U26071 ( .A(n16478), .B(n16474), .Z(n16850) );
  XNOR U26072 ( .A(n16473), .B(n16469), .Z(n16851) );
  XNOR U26073 ( .A(n16468), .B(n16464), .Z(n16852) );
  XNOR U26074 ( .A(n16463), .B(n16459), .Z(n16853) );
  XNOR U26075 ( .A(n16458), .B(n16454), .Z(n16854) );
  XNOR U26076 ( .A(n16453), .B(n16449), .Z(n16855) );
  XNOR U26077 ( .A(n16448), .B(n16444), .Z(n16856) );
  XNOR U26078 ( .A(n16443), .B(n16439), .Z(n16857) );
  XNOR U26079 ( .A(n16438), .B(n16434), .Z(n16858) );
  XNOR U26080 ( .A(n16433), .B(n16429), .Z(n16859) );
  XNOR U26081 ( .A(n16428), .B(n16424), .Z(n16860) );
  XNOR U26082 ( .A(n16423), .B(n16419), .Z(n16861) );
  XNOR U26083 ( .A(n16418), .B(n16414), .Z(n16862) );
  XNOR U26084 ( .A(n16413), .B(n16409), .Z(n16863) );
  XNOR U26085 ( .A(n16408), .B(n16404), .Z(n16864) );
  XNOR U26086 ( .A(n16403), .B(n16399), .Z(n16865) );
  XNOR U26087 ( .A(n16398), .B(n16394), .Z(n16866) );
  XNOR U26088 ( .A(n16393), .B(n16389), .Z(n16867) );
  XNOR U26089 ( .A(n16388), .B(n16384), .Z(n16868) );
  XNOR U26090 ( .A(n16383), .B(n16379), .Z(n16869) );
  XNOR U26091 ( .A(n16378), .B(n16374), .Z(n16870) );
  XNOR U26092 ( .A(n16373), .B(n16369), .Z(n16871) );
  XNOR U26093 ( .A(n16368), .B(n16364), .Z(n16872) );
  XNOR U26094 ( .A(n16363), .B(n16359), .Z(n16873) );
  XNOR U26095 ( .A(n16358), .B(n16354), .Z(n16874) );
  XNOR U26096 ( .A(n16353), .B(n16349), .Z(n16875) );
  XNOR U26097 ( .A(n16348), .B(n16344), .Z(n16876) );
  XNOR U26098 ( .A(n16343), .B(n16339), .Z(n16877) );
  XNOR U26099 ( .A(n16338), .B(n16334), .Z(n16878) );
  XNOR U26100 ( .A(n16333), .B(n16329), .Z(n16879) );
  XNOR U26101 ( .A(n16328), .B(n16324), .Z(n16880) );
  XNOR U26102 ( .A(n16323), .B(n16319), .Z(n16881) );
  XNOR U26103 ( .A(n16318), .B(n16314), .Z(n16882) );
  XNOR U26104 ( .A(n16313), .B(n16309), .Z(n16883) );
  XNOR U26105 ( .A(n16308), .B(n16304), .Z(n16884) );
  XNOR U26106 ( .A(n16303), .B(n16299), .Z(n16885) );
  XNOR U26107 ( .A(n16298), .B(n16294), .Z(n16886) );
  XNOR U26108 ( .A(n16293), .B(n16289), .Z(n16887) );
  XNOR U26109 ( .A(n16288), .B(n16284), .Z(n16888) );
  XOR U26110 ( .A(n16889), .B(n16283), .Z(n16284) );
  AND U26111 ( .A(a[0]), .B(b[102]), .Z(n16889) );
  XNOR U26112 ( .A(n16890), .B(n16283), .Z(n16285) );
  XNOR U26113 ( .A(n16891), .B(n16892), .Z(n16283) );
  ANDN U26114 ( .B(n16893), .A(n16894), .Z(n16891) );
  AND U26115 ( .A(a[1]), .B(b[101]), .Z(n16890) );
  XNOR U26116 ( .A(n16895), .B(n16288), .Z(n16290) );
  XOR U26117 ( .A(n16896), .B(n16897), .Z(n16288) );
  ANDN U26118 ( .B(n16898), .A(n16899), .Z(n16896) );
  AND U26119 ( .A(a[2]), .B(b[100]), .Z(n16895) );
  XNOR U26120 ( .A(n16900), .B(n16293), .Z(n16295) );
  XOR U26121 ( .A(n16901), .B(n16902), .Z(n16293) );
  ANDN U26122 ( .B(n16903), .A(n16904), .Z(n16901) );
  AND U26123 ( .A(a[3]), .B(b[99]), .Z(n16900) );
  XNOR U26124 ( .A(n16905), .B(n16298), .Z(n16300) );
  XOR U26125 ( .A(n16906), .B(n16907), .Z(n16298) );
  ANDN U26126 ( .B(n16908), .A(n16909), .Z(n16906) );
  AND U26127 ( .A(a[4]), .B(b[98]), .Z(n16905) );
  XNOR U26128 ( .A(n16910), .B(n16303), .Z(n16305) );
  XOR U26129 ( .A(n16911), .B(n16912), .Z(n16303) );
  ANDN U26130 ( .B(n16913), .A(n16914), .Z(n16911) );
  AND U26131 ( .A(a[5]), .B(b[97]), .Z(n16910) );
  XNOR U26132 ( .A(n16915), .B(n16308), .Z(n16310) );
  XOR U26133 ( .A(n16916), .B(n16917), .Z(n16308) );
  ANDN U26134 ( .B(n16918), .A(n16919), .Z(n16916) );
  AND U26135 ( .A(a[6]), .B(b[96]), .Z(n16915) );
  XNOR U26136 ( .A(n16920), .B(n16313), .Z(n16315) );
  XOR U26137 ( .A(n16921), .B(n16922), .Z(n16313) );
  ANDN U26138 ( .B(n16923), .A(n16924), .Z(n16921) );
  AND U26139 ( .A(a[7]), .B(b[95]), .Z(n16920) );
  XNOR U26140 ( .A(n16925), .B(n16318), .Z(n16320) );
  XOR U26141 ( .A(n16926), .B(n16927), .Z(n16318) );
  ANDN U26142 ( .B(n16928), .A(n16929), .Z(n16926) );
  AND U26143 ( .A(a[8]), .B(b[94]), .Z(n16925) );
  XNOR U26144 ( .A(n16930), .B(n16323), .Z(n16325) );
  XOR U26145 ( .A(n16931), .B(n16932), .Z(n16323) );
  ANDN U26146 ( .B(n16933), .A(n16934), .Z(n16931) );
  AND U26147 ( .A(a[9]), .B(b[93]), .Z(n16930) );
  XNOR U26148 ( .A(n16935), .B(n16328), .Z(n16330) );
  XOR U26149 ( .A(n16936), .B(n16937), .Z(n16328) );
  ANDN U26150 ( .B(n16938), .A(n16939), .Z(n16936) );
  AND U26151 ( .A(a[10]), .B(b[92]), .Z(n16935) );
  XNOR U26152 ( .A(n16940), .B(n16333), .Z(n16335) );
  XOR U26153 ( .A(n16941), .B(n16942), .Z(n16333) );
  ANDN U26154 ( .B(n16943), .A(n16944), .Z(n16941) );
  AND U26155 ( .A(a[11]), .B(b[91]), .Z(n16940) );
  XNOR U26156 ( .A(n16945), .B(n16338), .Z(n16340) );
  XOR U26157 ( .A(n16946), .B(n16947), .Z(n16338) );
  ANDN U26158 ( .B(n16948), .A(n16949), .Z(n16946) );
  AND U26159 ( .A(a[12]), .B(b[90]), .Z(n16945) );
  XNOR U26160 ( .A(n16950), .B(n16343), .Z(n16345) );
  XOR U26161 ( .A(n16951), .B(n16952), .Z(n16343) );
  ANDN U26162 ( .B(n16953), .A(n16954), .Z(n16951) );
  AND U26163 ( .A(a[13]), .B(b[89]), .Z(n16950) );
  XNOR U26164 ( .A(n16955), .B(n16348), .Z(n16350) );
  XOR U26165 ( .A(n16956), .B(n16957), .Z(n16348) );
  ANDN U26166 ( .B(n16958), .A(n16959), .Z(n16956) );
  AND U26167 ( .A(a[14]), .B(b[88]), .Z(n16955) );
  XNOR U26168 ( .A(n16960), .B(n16353), .Z(n16355) );
  XOR U26169 ( .A(n16961), .B(n16962), .Z(n16353) );
  ANDN U26170 ( .B(n16963), .A(n16964), .Z(n16961) );
  AND U26171 ( .A(a[15]), .B(b[87]), .Z(n16960) );
  XNOR U26172 ( .A(n16965), .B(n16358), .Z(n16360) );
  XOR U26173 ( .A(n16966), .B(n16967), .Z(n16358) );
  ANDN U26174 ( .B(n16968), .A(n16969), .Z(n16966) );
  AND U26175 ( .A(a[16]), .B(b[86]), .Z(n16965) );
  XNOR U26176 ( .A(n16970), .B(n16363), .Z(n16365) );
  XOR U26177 ( .A(n16971), .B(n16972), .Z(n16363) );
  ANDN U26178 ( .B(n16973), .A(n16974), .Z(n16971) );
  AND U26179 ( .A(a[17]), .B(b[85]), .Z(n16970) );
  XNOR U26180 ( .A(n16975), .B(n16368), .Z(n16370) );
  XOR U26181 ( .A(n16976), .B(n16977), .Z(n16368) );
  ANDN U26182 ( .B(n16978), .A(n16979), .Z(n16976) );
  AND U26183 ( .A(a[18]), .B(b[84]), .Z(n16975) );
  XNOR U26184 ( .A(n16980), .B(n16373), .Z(n16375) );
  XOR U26185 ( .A(n16981), .B(n16982), .Z(n16373) );
  ANDN U26186 ( .B(n16983), .A(n16984), .Z(n16981) );
  AND U26187 ( .A(a[19]), .B(b[83]), .Z(n16980) );
  XNOR U26188 ( .A(n16985), .B(n16378), .Z(n16380) );
  XOR U26189 ( .A(n16986), .B(n16987), .Z(n16378) );
  ANDN U26190 ( .B(n16988), .A(n16989), .Z(n16986) );
  AND U26191 ( .A(a[20]), .B(b[82]), .Z(n16985) );
  XNOR U26192 ( .A(n16990), .B(n16383), .Z(n16385) );
  XOR U26193 ( .A(n16991), .B(n16992), .Z(n16383) );
  ANDN U26194 ( .B(n16993), .A(n16994), .Z(n16991) );
  AND U26195 ( .A(a[21]), .B(b[81]), .Z(n16990) );
  XNOR U26196 ( .A(n16995), .B(n16388), .Z(n16390) );
  XOR U26197 ( .A(n16996), .B(n16997), .Z(n16388) );
  ANDN U26198 ( .B(n16998), .A(n16999), .Z(n16996) );
  AND U26199 ( .A(a[22]), .B(b[80]), .Z(n16995) );
  XNOR U26200 ( .A(n17000), .B(n16393), .Z(n16395) );
  XOR U26201 ( .A(n17001), .B(n17002), .Z(n16393) );
  ANDN U26202 ( .B(n17003), .A(n17004), .Z(n17001) );
  AND U26203 ( .A(a[23]), .B(b[79]), .Z(n17000) );
  XNOR U26204 ( .A(n17005), .B(n16398), .Z(n16400) );
  XOR U26205 ( .A(n17006), .B(n17007), .Z(n16398) );
  ANDN U26206 ( .B(n17008), .A(n17009), .Z(n17006) );
  AND U26207 ( .A(a[24]), .B(b[78]), .Z(n17005) );
  XNOR U26208 ( .A(n17010), .B(n16403), .Z(n16405) );
  XOR U26209 ( .A(n17011), .B(n17012), .Z(n16403) );
  ANDN U26210 ( .B(n17013), .A(n17014), .Z(n17011) );
  AND U26211 ( .A(a[25]), .B(b[77]), .Z(n17010) );
  XNOR U26212 ( .A(n17015), .B(n16408), .Z(n16410) );
  XOR U26213 ( .A(n17016), .B(n17017), .Z(n16408) );
  ANDN U26214 ( .B(n17018), .A(n17019), .Z(n17016) );
  AND U26215 ( .A(a[26]), .B(b[76]), .Z(n17015) );
  XNOR U26216 ( .A(n17020), .B(n16413), .Z(n16415) );
  XOR U26217 ( .A(n17021), .B(n17022), .Z(n16413) );
  ANDN U26218 ( .B(n17023), .A(n17024), .Z(n17021) );
  AND U26219 ( .A(a[27]), .B(b[75]), .Z(n17020) );
  XNOR U26220 ( .A(n17025), .B(n16418), .Z(n16420) );
  XOR U26221 ( .A(n17026), .B(n17027), .Z(n16418) );
  ANDN U26222 ( .B(n17028), .A(n17029), .Z(n17026) );
  AND U26223 ( .A(a[28]), .B(b[74]), .Z(n17025) );
  XNOR U26224 ( .A(n17030), .B(n16423), .Z(n16425) );
  XOR U26225 ( .A(n17031), .B(n17032), .Z(n16423) );
  ANDN U26226 ( .B(n17033), .A(n17034), .Z(n17031) );
  AND U26227 ( .A(a[29]), .B(b[73]), .Z(n17030) );
  XNOR U26228 ( .A(n17035), .B(n16428), .Z(n16430) );
  XOR U26229 ( .A(n17036), .B(n17037), .Z(n16428) );
  ANDN U26230 ( .B(n17038), .A(n17039), .Z(n17036) );
  AND U26231 ( .A(a[30]), .B(b[72]), .Z(n17035) );
  XNOR U26232 ( .A(n17040), .B(n16433), .Z(n16435) );
  XOR U26233 ( .A(n17041), .B(n17042), .Z(n16433) );
  ANDN U26234 ( .B(n17043), .A(n17044), .Z(n17041) );
  AND U26235 ( .A(a[31]), .B(b[71]), .Z(n17040) );
  XNOR U26236 ( .A(n17045), .B(n16438), .Z(n16440) );
  XOR U26237 ( .A(n17046), .B(n17047), .Z(n16438) );
  ANDN U26238 ( .B(n17048), .A(n17049), .Z(n17046) );
  AND U26239 ( .A(a[32]), .B(b[70]), .Z(n17045) );
  XNOR U26240 ( .A(n17050), .B(n16443), .Z(n16445) );
  XOR U26241 ( .A(n17051), .B(n17052), .Z(n16443) );
  ANDN U26242 ( .B(n17053), .A(n17054), .Z(n17051) );
  AND U26243 ( .A(a[33]), .B(b[69]), .Z(n17050) );
  XNOR U26244 ( .A(n17055), .B(n16448), .Z(n16450) );
  XOR U26245 ( .A(n17056), .B(n17057), .Z(n16448) );
  ANDN U26246 ( .B(n17058), .A(n17059), .Z(n17056) );
  AND U26247 ( .A(a[34]), .B(b[68]), .Z(n17055) );
  XNOR U26248 ( .A(n17060), .B(n16453), .Z(n16455) );
  XOR U26249 ( .A(n17061), .B(n17062), .Z(n16453) );
  ANDN U26250 ( .B(n17063), .A(n17064), .Z(n17061) );
  AND U26251 ( .A(a[35]), .B(b[67]), .Z(n17060) );
  XNOR U26252 ( .A(n17065), .B(n16458), .Z(n16460) );
  XOR U26253 ( .A(n17066), .B(n17067), .Z(n16458) );
  ANDN U26254 ( .B(n17068), .A(n17069), .Z(n17066) );
  AND U26255 ( .A(a[36]), .B(b[66]), .Z(n17065) );
  XNOR U26256 ( .A(n17070), .B(n16463), .Z(n16465) );
  XOR U26257 ( .A(n17071), .B(n17072), .Z(n16463) );
  ANDN U26258 ( .B(n17073), .A(n17074), .Z(n17071) );
  AND U26259 ( .A(a[37]), .B(b[65]), .Z(n17070) );
  XNOR U26260 ( .A(n17075), .B(n16468), .Z(n16470) );
  XOR U26261 ( .A(n17076), .B(n17077), .Z(n16468) );
  ANDN U26262 ( .B(n17078), .A(n17079), .Z(n17076) );
  AND U26263 ( .A(a[38]), .B(b[64]), .Z(n17075) );
  XNOR U26264 ( .A(n17080), .B(n16473), .Z(n16475) );
  XOR U26265 ( .A(n17081), .B(n17082), .Z(n16473) );
  ANDN U26266 ( .B(n17083), .A(n17084), .Z(n17081) );
  AND U26267 ( .A(a[39]), .B(b[63]), .Z(n17080) );
  XNOR U26268 ( .A(n17085), .B(n16478), .Z(n16480) );
  XOR U26269 ( .A(n17086), .B(n17087), .Z(n16478) );
  ANDN U26270 ( .B(n17088), .A(n17089), .Z(n17086) );
  AND U26271 ( .A(a[40]), .B(b[62]), .Z(n17085) );
  XNOR U26272 ( .A(n17090), .B(n16483), .Z(n16485) );
  XOR U26273 ( .A(n17091), .B(n17092), .Z(n16483) );
  ANDN U26274 ( .B(n17093), .A(n17094), .Z(n17091) );
  AND U26275 ( .A(a[41]), .B(b[61]), .Z(n17090) );
  XNOR U26276 ( .A(n17095), .B(n16488), .Z(n16490) );
  XOR U26277 ( .A(n17096), .B(n17097), .Z(n16488) );
  ANDN U26278 ( .B(n17098), .A(n17099), .Z(n17096) );
  AND U26279 ( .A(a[42]), .B(b[60]), .Z(n17095) );
  XNOR U26280 ( .A(n17100), .B(n16493), .Z(n16495) );
  XOR U26281 ( .A(n17101), .B(n17102), .Z(n16493) );
  ANDN U26282 ( .B(n17103), .A(n17104), .Z(n17101) );
  AND U26283 ( .A(a[43]), .B(b[59]), .Z(n17100) );
  XNOR U26284 ( .A(n17105), .B(n16498), .Z(n16500) );
  XOR U26285 ( .A(n17106), .B(n17107), .Z(n16498) );
  ANDN U26286 ( .B(n17108), .A(n17109), .Z(n17106) );
  AND U26287 ( .A(a[44]), .B(b[58]), .Z(n17105) );
  XNOR U26288 ( .A(n17110), .B(n16503), .Z(n16505) );
  XOR U26289 ( .A(n17111), .B(n17112), .Z(n16503) );
  ANDN U26290 ( .B(n17113), .A(n17114), .Z(n17111) );
  AND U26291 ( .A(a[45]), .B(b[57]), .Z(n17110) );
  XNOR U26292 ( .A(n17115), .B(n16508), .Z(n16510) );
  XOR U26293 ( .A(n17116), .B(n17117), .Z(n16508) );
  ANDN U26294 ( .B(n17118), .A(n17119), .Z(n17116) );
  AND U26295 ( .A(a[46]), .B(b[56]), .Z(n17115) );
  XNOR U26296 ( .A(n17120), .B(n16513), .Z(n16515) );
  XOR U26297 ( .A(n17121), .B(n17122), .Z(n16513) );
  ANDN U26298 ( .B(n17123), .A(n17124), .Z(n17121) );
  AND U26299 ( .A(a[47]), .B(b[55]), .Z(n17120) );
  XNOR U26300 ( .A(n17125), .B(n16518), .Z(n16520) );
  XOR U26301 ( .A(n17126), .B(n17127), .Z(n16518) );
  ANDN U26302 ( .B(n17128), .A(n17129), .Z(n17126) );
  AND U26303 ( .A(a[48]), .B(b[54]), .Z(n17125) );
  XNOR U26304 ( .A(n17130), .B(n16523), .Z(n16525) );
  XOR U26305 ( .A(n17131), .B(n17132), .Z(n16523) );
  ANDN U26306 ( .B(n17133), .A(n17134), .Z(n17131) );
  AND U26307 ( .A(a[49]), .B(b[53]), .Z(n17130) );
  XNOR U26308 ( .A(n17135), .B(n16528), .Z(n16530) );
  XOR U26309 ( .A(n17136), .B(n17137), .Z(n16528) );
  ANDN U26310 ( .B(n17138), .A(n17139), .Z(n17136) );
  AND U26311 ( .A(a[50]), .B(b[52]), .Z(n17135) );
  XNOR U26312 ( .A(n17140), .B(n16533), .Z(n16535) );
  XOR U26313 ( .A(n17141), .B(n17142), .Z(n16533) );
  ANDN U26314 ( .B(n17143), .A(n17144), .Z(n17141) );
  AND U26315 ( .A(a[51]), .B(b[51]), .Z(n17140) );
  XNOR U26316 ( .A(n17145), .B(n16538), .Z(n16540) );
  XOR U26317 ( .A(n17146), .B(n17147), .Z(n16538) );
  ANDN U26318 ( .B(n17148), .A(n17149), .Z(n17146) );
  AND U26319 ( .A(a[52]), .B(b[50]), .Z(n17145) );
  XNOR U26320 ( .A(n17150), .B(n16543), .Z(n16545) );
  XOR U26321 ( .A(n17151), .B(n17152), .Z(n16543) );
  ANDN U26322 ( .B(n17153), .A(n17154), .Z(n17151) );
  AND U26323 ( .A(a[53]), .B(b[49]), .Z(n17150) );
  XNOR U26324 ( .A(n17155), .B(n16548), .Z(n16550) );
  XOR U26325 ( .A(n17156), .B(n17157), .Z(n16548) );
  ANDN U26326 ( .B(n17158), .A(n17159), .Z(n17156) );
  AND U26327 ( .A(a[54]), .B(b[48]), .Z(n17155) );
  XNOR U26328 ( .A(n17160), .B(n16553), .Z(n16555) );
  XOR U26329 ( .A(n17161), .B(n17162), .Z(n16553) );
  ANDN U26330 ( .B(n17163), .A(n17164), .Z(n17161) );
  AND U26331 ( .A(a[55]), .B(b[47]), .Z(n17160) );
  XNOR U26332 ( .A(n17165), .B(n16558), .Z(n16560) );
  XOR U26333 ( .A(n17166), .B(n17167), .Z(n16558) );
  ANDN U26334 ( .B(n17168), .A(n17169), .Z(n17166) );
  AND U26335 ( .A(a[56]), .B(b[46]), .Z(n17165) );
  XNOR U26336 ( .A(n17170), .B(n16563), .Z(n16565) );
  XOR U26337 ( .A(n17171), .B(n17172), .Z(n16563) );
  ANDN U26338 ( .B(n17173), .A(n17174), .Z(n17171) );
  AND U26339 ( .A(a[57]), .B(b[45]), .Z(n17170) );
  XNOR U26340 ( .A(n17175), .B(n16568), .Z(n16570) );
  XOR U26341 ( .A(n17176), .B(n17177), .Z(n16568) );
  ANDN U26342 ( .B(n17178), .A(n17179), .Z(n17176) );
  AND U26343 ( .A(a[58]), .B(b[44]), .Z(n17175) );
  XNOR U26344 ( .A(n17180), .B(n16573), .Z(n16575) );
  XOR U26345 ( .A(n17181), .B(n17182), .Z(n16573) );
  ANDN U26346 ( .B(n17183), .A(n17184), .Z(n17181) );
  AND U26347 ( .A(a[59]), .B(b[43]), .Z(n17180) );
  XNOR U26348 ( .A(n17185), .B(n16578), .Z(n16580) );
  XOR U26349 ( .A(n17186), .B(n17187), .Z(n16578) );
  ANDN U26350 ( .B(n17188), .A(n17189), .Z(n17186) );
  AND U26351 ( .A(a[60]), .B(b[42]), .Z(n17185) );
  XNOR U26352 ( .A(n17190), .B(n16583), .Z(n16585) );
  XOR U26353 ( .A(n17191), .B(n17192), .Z(n16583) );
  ANDN U26354 ( .B(n17193), .A(n17194), .Z(n17191) );
  AND U26355 ( .A(a[61]), .B(b[41]), .Z(n17190) );
  XNOR U26356 ( .A(n17195), .B(n16588), .Z(n16590) );
  XOR U26357 ( .A(n17196), .B(n17197), .Z(n16588) );
  ANDN U26358 ( .B(n17198), .A(n17199), .Z(n17196) );
  AND U26359 ( .A(a[62]), .B(b[40]), .Z(n17195) );
  XNOR U26360 ( .A(n17200), .B(n16593), .Z(n16595) );
  XOR U26361 ( .A(n17201), .B(n17202), .Z(n16593) );
  ANDN U26362 ( .B(n17203), .A(n17204), .Z(n17201) );
  AND U26363 ( .A(a[63]), .B(b[39]), .Z(n17200) );
  XNOR U26364 ( .A(n17205), .B(n16598), .Z(n16600) );
  XOR U26365 ( .A(n17206), .B(n17207), .Z(n16598) );
  ANDN U26366 ( .B(n17208), .A(n17209), .Z(n17206) );
  AND U26367 ( .A(a[64]), .B(b[38]), .Z(n17205) );
  XNOR U26368 ( .A(n17210), .B(n16603), .Z(n16605) );
  XOR U26369 ( .A(n17211), .B(n17212), .Z(n16603) );
  ANDN U26370 ( .B(n17213), .A(n17214), .Z(n17211) );
  AND U26371 ( .A(a[65]), .B(b[37]), .Z(n17210) );
  XNOR U26372 ( .A(n17215), .B(n16608), .Z(n16610) );
  XOR U26373 ( .A(n17216), .B(n17217), .Z(n16608) );
  ANDN U26374 ( .B(n17218), .A(n17219), .Z(n17216) );
  AND U26375 ( .A(a[66]), .B(b[36]), .Z(n17215) );
  XNOR U26376 ( .A(n17220), .B(n16613), .Z(n16615) );
  XOR U26377 ( .A(n17221), .B(n17222), .Z(n16613) );
  ANDN U26378 ( .B(n17223), .A(n17224), .Z(n17221) );
  AND U26379 ( .A(a[67]), .B(b[35]), .Z(n17220) );
  XNOR U26380 ( .A(n17225), .B(n16618), .Z(n16620) );
  XOR U26381 ( .A(n17226), .B(n17227), .Z(n16618) );
  ANDN U26382 ( .B(n17228), .A(n17229), .Z(n17226) );
  AND U26383 ( .A(a[68]), .B(b[34]), .Z(n17225) );
  XNOR U26384 ( .A(n17230), .B(n16623), .Z(n16625) );
  XOR U26385 ( .A(n17231), .B(n17232), .Z(n16623) );
  ANDN U26386 ( .B(n17233), .A(n17234), .Z(n17231) );
  AND U26387 ( .A(a[69]), .B(b[33]), .Z(n17230) );
  XNOR U26388 ( .A(n17235), .B(n16628), .Z(n16630) );
  XOR U26389 ( .A(n17236), .B(n17237), .Z(n16628) );
  ANDN U26390 ( .B(n17238), .A(n17239), .Z(n17236) );
  AND U26391 ( .A(a[70]), .B(b[32]), .Z(n17235) );
  XNOR U26392 ( .A(n17240), .B(n16633), .Z(n16635) );
  XOR U26393 ( .A(n17241), .B(n17242), .Z(n16633) );
  ANDN U26394 ( .B(n17243), .A(n17244), .Z(n17241) );
  AND U26395 ( .A(a[71]), .B(b[31]), .Z(n17240) );
  XNOR U26396 ( .A(n17245), .B(n16638), .Z(n16640) );
  XOR U26397 ( .A(n17246), .B(n17247), .Z(n16638) );
  ANDN U26398 ( .B(n17248), .A(n17249), .Z(n17246) );
  AND U26399 ( .A(a[72]), .B(b[30]), .Z(n17245) );
  XNOR U26400 ( .A(n17250), .B(n16643), .Z(n16645) );
  XOR U26401 ( .A(n17251), .B(n17252), .Z(n16643) );
  ANDN U26402 ( .B(n17253), .A(n17254), .Z(n17251) );
  AND U26403 ( .A(a[73]), .B(b[29]), .Z(n17250) );
  XNOR U26404 ( .A(n17255), .B(n16648), .Z(n16650) );
  XOR U26405 ( .A(n17256), .B(n17257), .Z(n16648) );
  ANDN U26406 ( .B(n17258), .A(n17259), .Z(n17256) );
  AND U26407 ( .A(a[74]), .B(b[28]), .Z(n17255) );
  XNOR U26408 ( .A(n17260), .B(n16653), .Z(n16655) );
  XOR U26409 ( .A(n17261), .B(n17262), .Z(n16653) );
  ANDN U26410 ( .B(n17263), .A(n17264), .Z(n17261) );
  AND U26411 ( .A(a[75]), .B(b[27]), .Z(n17260) );
  XNOR U26412 ( .A(n17265), .B(n16658), .Z(n16660) );
  XOR U26413 ( .A(n17266), .B(n17267), .Z(n16658) );
  ANDN U26414 ( .B(n17268), .A(n17269), .Z(n17266) );
  AND U26415 ( .A(a[76]), .B(b[26]), .Z(n17265) );
  XNOR U26416 ( .A(n17270), .B(n16663), .Z(n16665) );
  XOR U26417 ( .A(n17271), .B(n17272), .Z(n16663) );
  ANDN U26418 ( .B(n17273), .A(n17274), .Z(n17271) );
  AND U26419 ( .A(a[77]), .B(b[25]), .Z(n17270) );
  XNOR U26420 ( .A(n17275), .B(n16668), .Z(n16670) );
  XOR U26421 ( .A(n17276), .B(n17277), .Z(n16668) );
  ANDN U26422 ( .B(n17278), .A(n17279), .Z(n17276) );
  AND U26423 ( .A(a[78]), .B(b[24]), .Z(n17275) );
  XNOR U26424 ( .A(n17280), .B(n16673), .Z(n16675) );
  XOR U26425 ( .A(n17281), .B(n17282), .Z(n16673) );
  ANDN U26426 ( .B(n17283), .A(n17284), .Z(n17281) );
  AND U26427 ( .A(a[79]), .B(b[23]), .Z(n17280) );
  XNOR U26428 ( .A(n17285), .B(n16678), .Z(n16680) );
  XOR U26429 ( .A(n17286), .B(n17287), .Z(n16678) );
  ANDN U26430 ( .B(n17288), .A(n17289), .Z(n17286) );
  AND U26431 ( .A(a[80]), .B(b[22]), .Z(n17285) );
  XNOR U26432 ( .A(n17290), .B(n16683), .Z(n16685) );
  XOR U26433 ( .A(n17291), .B(n17292), .Z(n16683) );
  ANDN U26434 ( .B(n17293), .A(n17294), .Z(n17291) );
  AND U26435 ( .A(a[81]), .B(b[21]), .Z(n17290) );
  XNOR U26436 ( .A(n17295), .B(n16688), .Z(n16690) );
  XOR U26437 ( .A(n17296), .B(n17297), .Z(n16688) );
  ANDN U26438 ( .B(n17298), .A(n17299), .Z(n17296) );
  AND U26439 ( .A(a[82]), .B(b[20]), .Z(n17295) );
  XNOR U26440 ( .A(n17300), .B(n16693), .Z(n16695) );
  XOR U26441 ( .A(n17301), .B(n17302), .Z(n16693) );
  ANDN U26442 ( .B(n17303), .A(n17304), .Z(n17301) );
  AND U26443 ( .A(a[83]), .B(b[19]), .Z(n17300) );
  XNOR U26444 ( .A(n17305), .B(n16698), .Z(n16700) );
  XOR U26445 ( .A(n17306), .B(n17307), .Z(n16698) );
  ANDN U26446 ( .B(n17308), .A(n17309), .Z(n17306) );
  AND U26447 ( .A(a[84]), .B(b[18]), .Z(n17305) );
  XNOR U26448 ( .A(n17310), .B(n16703), .Z(n16705) );
  XOR U26449 ( .A(n17311), .B(n17312), .Z(n16703) );
  ANDN U26450 ( .B(n17313), .A(n17314), .Z(n17311) );
  AND U26451 ( .A(a[85]), .B(b[17]), .Z(n17310) );
  XNOR U26452 ( .A(n17315), .B(n16708), .Z(n16710) );
  XOR U26453 ( .A(n17316), .B(n17317), .Z(n16708) );
  ANDN U26454 ( .B(n17318), .A(n17319), .Z(n17316) );
  AND U26455 ( .A(a[86]), .B(b[16]), .Z(n17315) );
  XNOR U26456 ( .A(n17320), .B(n16713), .Z(n16715) );
  XOR U26457 ( .A(n17321), .B(n17322), .Z(n16713) );
  ANDN U26458 ( .B(n17323), .A(n17324), .Z(n17321) );
  AND U26459 ( .A(a[87]), .B(b[15]), .Z(n17320) );
  XNOR U26460 ( .A(n17325), .B(n16718), .Z(n16720) );
  XOR U26461 ( .A(n17326), .B(n17327), .Z(n16718) );
  ANDN U26462 ( .B(n17328), .A(n17329), .Z(n17326) );
  AND U26463 ( .A(a[88]), .B(b[14]), .Z(n17325) );
  XNOR U26464 ( .A(n17330), .B(n16723), .Z(n16725) );
  XOR U26465 ( .A(n17331), .B(n17332), .Z(n16723) );
  ANDN U26466 ( .B(n17333), .A(n17334), .Z(n17331) );
  AND U26467 ( .A(a[89]), .B(b[13]), .Z(n17330) );
  XNOR U26468 ( .A(n17335), .B(n16728), .Z(n16730) );
  XOR U26469 ( .A(n17336), .B(n17337), .Z(n16728) );
  ANDN U26470 ( .B(n17338), .A(n17339), .Z(n17336) );
  AND U26471 ( .A(a[90]), .B(b[12]), .Z(n17335) );
  XNOR U26472 ( .A(n17340), .B(n16733), .Z(n16735) );
  XOR U26473 ( .A(n17341), .B(n17342), .Z(n16733) );
  ANDN U26474 ( .B(n17343), .A(n17344), .Z(n17341) );
  AND U26475 ( .A(a[91]), .B(b[11]), .Z(n17340) );
  XNOR U26476 ( .A(n17345), .B(n16738), .Z(n16740) );
  XOR U26477 ( .A(n17346), .B(n17347), .Z(n16738) );
  ANDN U26478 ( .B(n17348), .A(n17349), .Z(n17346) );
  AND U26479 ( .A(a[92]), .B(b[10]), .Z(n17345) );
  XNOR U26480 ( .A(n17350), .B(n16743), .Z(n16745) );
  XOR U26481 ( .A(n17351), .B(n17352), .Z(n16743) );
  ANDN U26482 ( .B(n17353), .A(n17354), .Z(n17351) );
  AND U26483 ( .A(b[9]), .B(a[93]), .Z(n17350) );
  XNOR U26484 ( .A(n17355), .B(n16748), .Z(n16750) );
  XOR U26485 ( .A(n17356), .B(n17357), .Z(n16748) );
  ANDN U26486 ( .B(n17358), .A(n17359), .Z(n17356) );
  AND U26487 ( .A(b[8]), .B(a[94]), .Z(n17355) );
  XNOR U26488 ( .A(n17360), .B(n16753), .Z(n16755) );
  XOR U26489 ( .A(n17361), .B(n17362), .Z(n16753) );
  ANDN U26490 ( .B(n17363), .A(n17364), .Z(n17361) );
  AND U26491 ( .A(b[7]), .B(a[95]), .Z(n17360) );
  XNOR U26492 ( .A(n17365), .B(n16758), .Z(n16760) );
  XOR U26493 ( .A(n17366), .B(n17367), .Z(n16758) );
  ANDN U26494 ( .B(n17368), .A(n17369), .Z(n17366) );
  AND U26495 ( .A(b[6]), .B(a[96]), .Z(n17365) );
  XNOR U26496 ( .A(n17370), .B(n16763), .Z(n16765) );
  XOR U26497 ( .A(n17371), .B(n17372), .Z(n16763) );
  ANDN U26498 ( .B(n17373), .A(n17374), .Z(n17371) );
  AND U26499 ( .A(b[5]), .B(a[97]), .Z(n17370) );
  XNOR U26500 ( .A(n17375), .B(n16768), .Z(n16770) );
  XOR U26501 ( .A(n17376), .B(n17377), .Z(n16768) );
  ANDN U26502 ( .B(n17378), .A(n17379), .Z(n17376) );
  AND U26503 ( .A(b[4]), .B(a[98]), .Z(n17375) );
  XNOR U26504 ( .A(n17380), .B(n17381), .Z(n16782) );
  NANDN U26505 ( .A(n17382), .B(n17383), .Z(n17381) );
  XNOR U26506 ( .A(n17384), .B(n16773), .Z(n16775) );
  XNOR U26507 ( .A(n17385), .B(n17386), .Z(n16773) );
  AND U26508 ( .A(n17387), .B(n17388), .Z(n17385) );
  AND U26509 ( .A(b[3]), .B(a[99]), .Z(n17384) );
  NAND U26510 ( .A(a[102]), .B(b[0]), .Z(n16178) );
  XNOR U26511 ( .A(n16788), .B(n16789), .Z(c[101]) );
  XNOR U26512 ( .A(n17382), .B(n17383), .Z(n16789) );
  XOR U26513 ( .A(n17380), .B(n17389), .Z(n17383) );
  NAND U26514 ( .A(b[1]), .B(a[100]), .Z(n17389) );
  XOR U26515 ( .A(n17388), .B(n17390), .Z(n17382) );
  XOR U26516 ( .A(n17380), .B(n17387), .Z(n17390) );
  XNOR U26517 ( .A(n17391), .B(n17386), .Z(n17387) );
  AND U26518 ( .A(b[2]), .B(a[99]), .Z(n17391) );
  NANDN U26519 ( .A(n17392), .B(n17393), .Z(n17380) );
  XOR U26520 ( .A(n17386), .B(n17378), .Z(n17394) );
  XNOR U26521 ( .A(n17377), .B(n17373), .Z(n17395) );
  XNOR U26522 ( .A(n17372), .B(n17368), .Z(n17396) );
  XNOR U26523 ( .A(n17367), .B(n17363), .Z(n17397) );
  XNOR U26524 ( .A(n17362), .B(n17358), .Z(n17398) );
  XNOR U26525 ( .A(n17357), .B(n17353), .Z(n17399) );
  XNOR U26526 ( .A(n17352), .B(n17348), .Z(n17400) );
  XNOR U26527 ( .A(n17347), .B(n17343), .Z(n17401) );
  XNOR U26528 ( .A(n17342), .B(n17338), .Z(n17402) );
  XNOR U26529 ( .A(n17337), .B(n17333), .Z(n17403) );
  XNOR U26530 ( .A(n17332), .B(n17328), .Z(n17404) );
  XNOR U26531 ( .A(n17327), .B(n17323), .Z(n17405) );
  XNOR U26532 ( .A(n17322), .B(n17318), .Z(n17406) );
  XNOR U26533 ( .A(n17317), .B(n17313), .Z(n17407) );
  XNOR U26534 ( .A(n17312), .B(n17308), .Z(n17408) );
  XNOR U26535 ( .A(n17307), .B(n17303), .Z(n17409) );
  XNOR U26536 ( .A(n17302), .B(n17298), .Z(n17410) );
  XNOR U26537 ( .A(n17297), .B(n17293), .Z(n17411) );
  XNOR U26538 ( .A(n17292), .B(n17288), .Z(n17412) );
  XNOR U26539 ( .A(n17287), .B(n17283), .Z(n17413) );
  XNOR U26540 ( .A(n17282), .B(n17278), .Z(n17414) );
  XNOR U26541 ( .A(n17277), .B(n17273), .Z(n17415) );
  XNOR U26542 ( .A(n17272), .B(n17268), .Z(n17416) );
  XNOR U26543 ( .A(n17267), .B(n17263), .Z(n17417) );
  XNOR U26544 ( .A(n17262), .B(n17258), .Z(n17418) );
  XNOR U26545 ( .A(n17257), .B(n17253), .Z(n17419) );
  XNOR U26546 ( .A(n17252), .B(n17248), .Z(n17420) );
  XNOR U26547 ( .A(n17247), .B(n17243), .Z(n17421) );
  XNOR U26548 ( .A(n17242), .B(n17238), .Z(n17422) );
  XNOR U26549 ( .A(n17237), .B(n17233), .Z(n17423) );
  XNOR U26550 ( .A(n17232), .B(n17228), .Z(n17424) );
  XNOR U26551 ( .A(n17227), .B(n17223), .Z(n17425) );
  XNOR U26552 ( .A(n17222), .B(n17218), .Z(n17426) );
  XNOR U26553 ( .A(n17217), .B(n17213), .Z(n17427) );
  XNOR U26554 ( .A(n17212), .B(n17208), .Z(n17428) );
  XNOR U26555 ( .A(n17207), .B(n17203), .Z(n17429) );
  XNOR U26556 ( .A(n17202), .B(n17198), .Z(n17430) );
  XNOR U26557 ( .A(n17197), .B(n17193), .Z(n17431) );
  XNOR U26558 ( .A(n17192), .B(n17188), .Z(n17432) );
  XNOR U26559 ( .A(n17187), .B(n17183), .Z(n17433) );
  XNOR U26560 ( .A(n17182), .B(n17178), .Z(n17434) );
  XNOR U26561 ( .A(n17177), .B(n17173), .Z(n17435) );
  XNOR U26562 ( .A(n17172), .B(n17168), .Z(n17436) );
  XNOR U26563 ( .A(n17167), .B(n17163), .Z(n17437) );
  XNOR U26564 ( .A(n17162), .B(n17158), .Z(n17438) );
  XNOR U26565 ( .A(n17157), .B(n17153), .Z(n17439) );
  XNOR U26566 ( .A(n17152), .B(n17148), .Z(n17440) );
  XNOR U26567 ( .A(n17147), .B(n17143), .Z(n17441) );
  XNOR U26568 ( .A(n17142), .B(n17138), .Z(n17442) );
  XNOR U26569 ( .A(n17137), .B(n17133), .Z(n17443) );
  XNOR U26570 ( .A(n17132), .B(n17128), .Z(n17444) );
  XNOR U26571 ( .A(n17127), .B(n17123), .Z(n17445) );
  XNOR U26572 ( .A(n17122), .B(n17118), .Z(n17446) );
  XNOR U26573 ( .A(n17117), .B(n17113), .Z(n17447) );
  XNOR U26574 ( .A(n17112), .B(n17108), .Z(n17448) );
  XNOR U26575 ( .A(n17107), .B(n17103), .Z(n17449) );
  XNOR U26576 ( .A(n17102), .B(n17098), .Z(n17450) );
  XNOR U26577 ( .A(n17097), .B(n17093), .Z(n17451) );
  XNOR U26578 ( .A(n17092), .B(n17088), .Z(n17452) );
  XNOR U26579 ( .A(n17087), .B(n17083), .Z(n17453) );
  XNOR U26580 ( .A(n17082), .B(n17078), .Z(n17454) );
  XNOR U26581 ( .A(n17077), .B(n17073), .Z(n17455) );
  XNOR U26582 ( .A(n17072), .B(n17068), .Z(n17456) );
  XNOR U26583 ( .A(n17067), .B(n17063), .Z(n17457) );
  XNOR U26584 ( .A(n17062), .B(n17058), .Z(n17458) );
  XNOR U26585 ( .A(n17057), .B(n17053), .Z(n17459) );
  XNOR U26586 ( .A(n17052), .B(n17048), .Z(n17460) );
  XNOR U26587 ( .A(n17047), .B(n17043), .Z(n17461) );
  XNOR U26588 ( .A(n17042), .B(n17038), .Z(n17462) );
  XNOR U26589 ( .A(n17037), .B(n17033), .Z(n17463) );
  XNOR U26590 ( .A(n17032), .B(n17028), .Z(n17464) );
  XNOR U26591 ( .A(n17027), .B(n17023), .Z(n17465) );
  XNOR U26592 ( .A(n17022), .B(n17018), .Z(n17466) );
  XNOR U26593 ( .A(n17017), .B(n17013), .Z(n17467) );
  XNOR U26594 ( .A(n17012), .B(n17008), .Z(n17468) );
  XNOR U26595 ( .A(n17007), .B(n17003), .Z(n17469) );
  XNOR U26596 ( .A(n17002), .B(n16998), .Z(n17470) );
  XNOR U26597 ( .A(n16997), .B(n16993), .Z(n17471) );
  XNOR U26598 ( .A(n16992), .B(n16988), .Z(n17472) );
  XNOR U26599 ( .A(n16987), .B(n16983), .Z(n17473) );
  XNOR U26600 ( .A(n16982), .B(n16978), .Z(n17474) );
  XNOR U26601 ( .A(n16977), .B(n16973), .Z(n17475) );
  XNOR U26602 ( .A(n16972), .B(n16968), .Z(n17476) );
  XNOR U26603 ( .A(n16967), .B(n16963), .Z(n17477) );
  XNOR U26604 ( .A(n16962), .B(n16958), .Z(n17478) );
  XNOR U26605 ( .A(n16957), .B(n16953), .Z(n17479) );
  XNOR U26606 ( .A(n16952), .B(n16948), .Z(n17480) );
  XNOR U26607 ( .A(n16947), .B(n16943), .Z(n17481) );
  XNOR U26608 ( .A(n16942), .B(n16938), .Z(n17482) );
  XNOR U26609 ( .A(n16937), .B(n16933), .Z(n17483) );
  XNOR U26610 ( .A(n16932), .B(n16928), .Z(n17484) );
  XNOR U26611 ( .A(n16927), .B(n16923), .Z(n17485) );
  XNOR U26612 ( .A(n16922), .B(n16918), .Z(n17486) );
  XNOR U26613 ( .A(n16917), .B(n16913), .Z(n17487) );
  XNOR U26614 ( .A(n16912), .B(n16908), .Z(n17488) );
  XNOR U26615 ( .A(n16907), .B(n16903), .Z(n17489) );
  XNOR U26616 ( .A(n16902), .B(n16898), .Z(n17490) );
  XNOR U26617 ( .A(n16897), .B(n16893), .Z(n17491) );
  XNOR U26618 ( .A(n17492), .B(n16892), .Z(n16893) );
  AND U26619 ( .A(a[0]), .B(b[101]), .Z(n17492) );
  XOR U26620 ( .A(n17493), .B(n16892), .Z(n16894) );
  XNOR U26621 ( .A(n17494), .B(n17495), .Z(n16892) );
  ANDN U26622 ( .B(n17496), .A(n17497), .Z(n17494) );
  AND U26623 ( .A(a[1]), .B(b[100]), .Z(n17493) );
  XNOR U26624 ( .A(n17498), .B(n16897), .Z(n16899) );
  XOR U26625 ( .A(n17499), .B(n17500), .Z(n16897) );
  ANDN U26626 ( .B(n17501), .A(n17502), .Z(n17499) );
  AND U26627 ( .A(a[2]), .B(b[99]), .Z(n17498) );
  XNOR U26628 ( .A(n17503), .B(n16902), .Z(n16904) );
  XOR U26629 ( .A(n17504), .B(n17505), .Z(n16902) );
  ANDN U26630 ( .B(n17506), .A(n17507), .Z(n17504) );
  AND U26631 ( .A(a[3]), .B(b[98]), .Z(n17503) );
  XNOR U26632 ( .A(n17508), .B(n16907), .Z(n16909) );
  XOR U26633 ( .A(n17509), .B(n17510), .Z(n16907) );
  ANDN U26634 ( .B(n17511), .A(n17512), .Z(n17509) );
  AND U26635 ( .A(a[4]), .B(b[97]), .Z(n17508) );
  XNOR U26636 ( .A(n17513), .B(n16912), .Z(n16914) );
  XOR U26637 ( .A(n17514), .B(n17515), .Z(n16912) );
  ANDN U26638 ( .B(n17516), .A(n17517), .Z(n17514) );
  AND U26639 ( .A(a[5]), .B(b[96]), .Z(n17513) );
  XNOR U26640 ( .A(n17518), .B(n16917), .Z(n16919) );
  XOR U26641 ( .A(n17519), .B(n17520), .Z(n16917) );
  ANDN U26642 ( .B(n17521), .A(n17522), .Z(n17519) );
  AND U26643 ( .A(a[6]), .B(b[95]), .Z(n17518) );
  XNOR U26644 ( .A(n17523), .B(n16922), .Z(n16924) );
  XOR U26645 ( .A(n17524), .B(n17525), .Z(n16922) );
  ANDN U26646 ( .B(n17526), .A(n17527), .Z(n17524) );
  AND U26647 ( .A(a[7]), .B(b[94]), .Z(n17523) );
  XNOR U26648 ( .A(n17528), .B(n16927), .Z(n16929) );
  XOR U26649 ( .A(n17529), .B(n17530), .Z(n16927) );
  ANDN U26650 ( .B(n17531), .A(n17532), .Z(n17529) );
  AND U26651 ( .A(a[8]), .B(b[93]), .Z(n17528) );
  XNOR U26652 ( .A(n17533), .B(n16932), .Z(n16934) );
  XOR U26653 ( .A(n17534), .B(n17535), .Z(n16932) );
  ANDN U26654 ( .B(n17536), .A(n17537), .Z(n17534) );
  AND U26655 ( .A(a[9]), .B(b[92]), .Z(n17533) );
  XNOR U26656 ( .A(n17538), .B(n16937), .Z(n16939) );
  XOR U26657 ( .A(n17539), .B(n17540), .Z(n16937) );
  ANDN U26658 ( .B(n17541), .A(n17542), .Z(n17539) );
  AND U26659 ( .A(a[10]), .B(b[91]), .Z(n17538) );
  XNOR U26660 ( .A(n17543), .B(n16942), .Z(n16944) );
  XOR U26661 ( .A(n17544), .B(n17545), .Z(n16942) );
  ANDN U26662 ( .B(n17546), .A(n17547), .Z(n17544) );
  AND U26663 ( .A(a[11]), .B(b[90]), .Z(n17543) );
  XNOR U26664 ( .A(n17548), .B(n16947), .Z(n16949) );
  XOR U26665 ( .A(n17549), .B(n17550), .Z(n16947) );
  ANDN U26666 ( .B(n17551), .A(n17552), .Z(n17549) );
  AND U26667 ( .A(a[12]), .B(b[89]), .Z(n17548) );
  XNOR U26668 ( .A(n17553), .B(n16952), .Z(n16954) );
  XOR U26669 ( .A(n17554), .B(n17555), .Z(n16952) );
  ANDN U26670 ( .B(n17556), .A(n17557), .Z(n17554) );
  AND U26671 ( .A(a[13]), .B(b[88]), .Z(n17553) );
  XNOR U26672 ( .A(n17558), .B(n16957), .Z(n16959) );
  XOR U26673 ( .A(n17559), .B(n17560), .Z(n16957) );
  ANDN U26674 ( .B(n17561), .A(n17562), .Z(n17559) );
  AND U26675 ( .A(a[14]), .B(b[87]), .Z(n17558) );
  XNOR U26676 ( .A(n17563), .B(n16962), .Z(n16964) );
  XOR U26677 ( .A(n17564), .B(n17565), .Z(n16962) );
  ANDN U26678 ( .B(n17566), .A(n17567), .Z(n17564) );
  AND U26679 ( .A(a[15]), .B(b[86]), .Z(n17563) );
  XNOR U26680 ( .A(n17568), .B(n16967), .Z(n16969) );
  XOR U26681 ( .A(n17569), .B(n17570), .Z(n16967) );
  ANDN U26682 ( .B(n17571), .A(n17572), .Z(n17569) );
  AND U26683 ( .A(a[16]), .B(b[85]), .Z(n17568) );
  XNOR U26684 ( .A(n17573), .B(n16972), .Z(n16974) );
  XOR U26685 ( .A(n17574), .B(n17575), .Z(n16972) );
  ANDN U26686 ( .B(n17576), .A(n17577), .Z(n17574) );
  AND U26687 ( .A(a[17]), .B(b[84]), .Z(n17573) );
  XNOR U26688 ( .A(n17578), .B(n16977), .Z(n16979) );
  XOR U26689 ( .A(n17579), .B(n17580), .Z(n16977) );
  ANDN U26690 ( .B(n17581), .A(n17582), .Z(n17579) );
  AND U26691 ( .A(a[18]), .B(b[83]), .Z(n17578) );
  XNOR U26692 ( .A(n17583), .B(n16982), .Z(n16984) );
  XOR U26693 ( .A(n17584), .B(n17585), .Z(n16982) );
  ANDN U26694 ( .B(n17586), .A(n17587), .Z(n17584) );
  AND U26695 ( .A(a[19]), .B(b[82]), .Z(n17583) );
  XNOR U26696 ( .A(n17588), .B(n16987), .Z(n16989) );
  XOR U26697 ( .A(n17589), .B(n17590), .Z(n16987) );
  ANDN U26698 ( .B(n17591), .A(n17592), .Z(n17589) );
  AND U26699 ( .A(a[20]), .B(b[81]), .Z(n17588) );
  XNOR U26700 ( .A(n17593), .B(n16992), .Z(n16994) );
  XOR U26701 ( .A(n17594), .B(n17595), .Z(n16992) );
  ANDN U26702 ( .B(n17596), .A(n17597), .Z(n17594) );
  AND U26703 ( .A(a[21]), .B(b[80]), .Z(n17593) );
  XNOR U26704 ( .A(n17598), .B(n16997), .Z(n16999) );
  XOR U26705 ( .A(n17599), .B(n17600), .Z(n16997) );
  ANDN U26706 ( .B(n17601), .A(n17602), .Z(n17599) );
  AND U26707 ( .A(a[22]), .B(b[79]), .Z(n17598) );
  XNOR U26708 ( .A(n17603), .B(n17002), .Z(n17004) );
  XOR U26709 ( .A(n17604), .B(n17605), .Z(n17002) );
  ANDN U26710 ( .B(n17606), .A(n17607), .Z(n17604) );
  AND U26711 ( .A(a[23]), .B(b[78]), .Z(n17603) );
  XNOR U26712 ( .A(n17608), .B(n17007), .Z(n17009) );
  XOR U26713 ( .A(n17609), .B(n17610), .Z(n17007) );
  ANDN U26714 ( .B(n17611), .A(n17612), .Z(n17609) );
  AND U26715 ( .A(a[24]), .B(b[77]), .Z(n17608) );
  XNOR U26716 ( .A(n17613), .B(n17012), .Z(n17014) );
  XOR U26717 ( .A(n17614), .B(n17615), .Z(n17012) );
  ANDN U26718 ( .B(n17616), .A(n17617), .Z(n17614) );
  AND U26719 ( .A(a[25]), .B(b[76]), .Z(n17613) );
  XNOR U26720 ( .A(n17618), .B(n17017), .Z(n17019) );
  XOR U26721 ( .A(n17619), .B(n17620), .Z(n17017) );
  ANDN U26722 ( .B(n17621), .A(n17622), .Z(n17619) );
  AND U26723 ( .A(a[26]), .B(b[75]), .Z(n17618) );
  XNOR U26724 ( .A(n17623), .B(n17022), .Z(n17024) );
  XOR U26725 ( .A(n17624), .B(n17625), .Z(n17022) );
  ANDN U26726 ( .B(n17626), .A(n17627), .Z(n17624) );
  AND U26727 ( .A(a[27]), .B(b[74]), .Z(n17623) );
  XNOR U26728 ( .A(n17628), .B(n17027), .Z(n17029) );
  XOR U26729 ( .A(n17629), .B(n17630), .Z(n17027) );
  ANDN U26730 ( .B(n17631), .A(n17632), .Z(n17629) );
  AND U26731 ( .A(a[28]), .B(b[73]), .Z(n17628) );
  XNOR U26732 ( .A(n17633), .B(n17032), .Z(n17034) );
  XOR U26733 ( .A(n17634), .B(n17635), .Z(n17032) );
  ANDN U26734 ( .B(n17636), .A(n17637), .Z(n17634) );
  AND U26735 ( .A(a[29]), .B(b[72]), .Z(n17633) );
  XNOR U26736 ( .A(n17638), .B(n17037), .Z(n17039) );
  XOR U26737 ( .A(n17639), .B(n17640), .Z(n17037) );
  ANDN U26738 ( .B(n17641), .A(n17642), .Z(n17639) );
  AND U26739 ( .A(a[30]), .B(b[71]), .Z(n17638) );
  XNOR U26740 ( .A(n17643), .B(n17042), .Z(n17044) );
  XOR U26741 ( .A(n17644), .B(n17645), .Z(n17042) );
  ANDN U26742 ( .B(n17646), .A(n17647), .Z(n17644) );
  AND U26743 ( .A(a[31]), .B(b[70]), .Z(n17643) );
  XNOR U26744 ( .A(n17648), .B(n17047), .Z(n17049) );
  XOR U26745 ( .A(n17649), .B(n17650), .Z(n17047) );
  ANDN U26746 ( .B(n17651), .A(n17652), .Z(n17649) );
  AND U26747 ( .A(a[32]), .B(b[69]), .Z(n17648) );
  XNOR U26748 ( .A(n17653), .B(n17052), .Z(n17054) );
  XOR U26749 ( .A(n17654), .B(n17655), .Z(n17052) );
  ANDN U26750 ( .B(n17656), .A(n17657), .Z(n17654) );
  AND U26751 ( .A(a[33]), .B(b[68]), .Z(n17653) );
  XNOR U26752 ( .A(n17658), .B(n17057), .Z(n17059) );
  XOR U26753 ( .A(n17659), .B(n17660), .Z(n17057) );
  ANDN U26754 ( .B(n17661), .A(n17662), .Z(n17659) );
  AND U26755 ( .A(a[34]), .B(b[67]), .Z(n17658) );
  XNOR U26756 ( .A(n17663), .B(n17062), .Z(n17064) );
  XOR U26757 ( .A(n17664), .B(n17665), .Z(n17062) );
  ANDN U26758 ( .B(n17666), .A(n17667), .Z(n17664) );
  AND U26759 ( .A(a[35]), .B(b[66]), .Z(n17663) );
  XNOR U26760 ( .A(n17668), .B(n17067), .Z(n17069) );
  XOR U26761 ( .A(n17669), .B(n17670), .Z(n17067) );
  ANDN U26762 ( .B(n17671), .A(n17672), .Z(n17669) );
  AND U26763 ( .A(a[36]), .B(b[65]), .Z(n17668) );
  XNOR U26764 ( .A(n17673), .B(n17072), .Z(n17074) );
  XOR U26765 ( .A(n17674), .B(n17675), .Z(n17072) );
  ANDN U26766 ( .B(n17676), .A(n17677), .Z(n17674) );
  AND U26767 ( .A(a[37]), .B(b[64]), .Z(n17673) );
  XNOR U26768 ( .A(n17678), .B(n17077), .Z(n17079) );
  XOR U26769 ( .A(n17679), .B(n17680), .Z(n17077) );
  ANDN U26770 ( .B(n17681), .A(n17682), .Z(n17679) );
  AND U26771 ( .A(a[38]), .B(b[63]), .Z(n17678) );
  XNOR U26772 ( .A(n17683), .B(n17082), .Z(n17084) );
  XOR U26773 ( .A(n17684), .B(n17685), .Z(n17082) );
  ANDN U26774 ( .B(n17686), .A(n17687), .Z(n17684) );
  AND U26775 ( .A(a[39]), .B(b[62]), .Z(n17683) );
  XNOR U26776 ( .A(n17688), .B(n17087), .Z(n17089) );
  XOR U26777 ( .A(n17689), .B(n17690), .Z(n17087) );
  ANDN U26778 ( .B(n17691), .A(n17692), .Z(n17689) );
  AND U26779 ( .A(a[40]), .B(b[61]), .Z(n17688) );
  XNOR U26780 ( .A(n17693), .B(n17092), .Z(n17094) );
  XOR U26781 ( .A(n17694), .B(n17695), .Z(n17092) );
  ANDN U26782 ( .B(n17696), .A(n17697), .Z(n17694) );
  AND U26783 ( .A(a[41]), .B(b[60]), .Z(n17693) );
  XNOR U26784 ( .A(n17698), .B(n17097), .Z(n17099) );
  XOR U26785 ( .A(n17699), .B(n17700), .Z(n17097) );
  ANDN U26786 ( .B(n17701), .A(n17702), .Z(n17699) );
  AND U26787 ( .A(a[42]), .B(b[59]), .Z(n17698) );
  XNOR U26788 ( .A(n17703), .B(n17102), .Z(n17104) );
  XOR U26789 ( .A(n17704), .B(n17705), .Z(n17102) );
  ANDN U26790 ( .B(n17706), .A(n17707), .Z(n17704) );
  AND U26791 ( .A(a[43]), .B(b[58]), .Z(n17703) );
  XNOR U26792 ( .A(n17708), .B(n17107), .Z(n17109) );
  XOR U26793 ( .A(n17709), .B(n17710), .Z(n17107) );
  ANDN U26794 ( .B(n17711), .A(n17712), .Z(n17709) );
  AND U26795 ( .A(a[44]), .B(b[57]), .Z(n17708) );
  XNOR U26796 ( .A(n17713), .B(n17112), .Z(n17114) );
  XOR U26797 ( .A(n17714), .B(n17715), .Z(n17112) );
  ANDN U26798 ( .B(n17716), .A(n17717), .Z(n17714) );
  AND U26799 ( .A(a[45]), .B(b[56]), .Z(n17713) );
  XNOR U26800 ( .A(n17718), .B(n17117), .Z(n17119) );
  XOR U26801 ( .A(n17719), .B(n17720), .Z(n17117) );
  ANDN U26802 ( .B(n17721), .A(n17722), .Z(n17719) );
  AND U26803 ( .A(a[46]), .B(b[55]), .Z(n17718) );
  XNOR U26804 ( .A(n17723), .B(n17122), .Z(n17124) );
  XOR U26805 ( .A(n17724), .B(n17725), .Z(n17122) );
  ANDN U26806 ( .B(n17726), .A(n17727), .Z(n17724) );
  AND U26807 ( .A(a[47]), .B(b[54]), .Z(n17723) );
  XNOR U26808 ( .A(n17728), .B(n17127), .Z(n17129) );
  XOR U26809 ( .A(n17729), .B(n17730), .Z(n17127) );
  ANDN U26810 ( .B(n17731), .A(n17732), .Z(n17729) );
  AND U26811 ( .A(a[48]), .B(b[53]), .Z(n17728) );
  XNOR U26812 ( .A(n17733), .B(n17132), .Z(n17134) );
  XOR U26813 ( .A(n17734), .B(n17735), .Z(n17132) );
  ANDN U26814 ( .B(n17736), .A(n17737), .Z(n17734) );
  AND U26815 ( .A(a[49]), .B(b[52]), .Z(n17733) );
  XNOR U26816 ( .A(n17738), .B(n17137), .Z(n17139) );
  XOR U26817 ( .A(n17739), .B(n17740), .Z(n17137) );
  ANDN U26818 ( .B(n17741), .A(n17742), .Z(n17739) );
  AND U26819 ( .A(a[50]), .B(b[51]), .Z(n17738) );
  XNOR U26820 ( .A(n17743), .B(n17142), .Z(n17144) );
  XOR U26821 ( .A(n17744), .B(n17745), .Z(n17142) );
  ANDN U26822 ( .B(n17746), .A(n17747), .Z(n17744) );
  AND U26823 ( .A(a[51]), .B(b[50]), .Z(n17743) );
  XNOR U26824 ( .A(n17748), .B(n17147), .Z(n17149) );
  XOR U26825 ( .A(n17749), .B(n17750), .Z(n17147) );
  ANDN U26826 ( .B(n17751), .A(n17752), .Z(n17749) );
  AND U26827 ( .A(a[52]), .B(b[49]), .Z(n17748) );
  XNOR U26828 ( .A(n17753), .B(n17152), .Z(n17154) );
  XOR U26829 ( .A(n17754), .B(n17755), .Z(n17152) );
  ANDN U26830 ( .B(n17756), .A(n17757), .Z(n17754) );
  AND U26831 ( .A(a[53]), .B(b[48]), .Z(n17753) );
  XNOR U26832 ( .A(n17758), .B(n17157), .Z(n17159) );
  XOR U26833 ( .A(n17759), .B(n17760), .Z(n17157) );
  ANDN U26834 ( .B(n17761), .A(n17762), .Z(n17759) );
  AND U26835 ( .A(a[54]), .B(b[47]), .Z(n17758) );
  XNOR U26836 ( .A(n17763), .B(n17162), .Z(n17164) );
  XOR U26837 ( .A(n17764), .B(n17765), .Z(n17162) );
  ANDN U26838 ( .B(n17766), .A(n17767), .Z(n17764) );
  AND U26839 ( .A(a[55]), .B(b[46]), .Z(n17763) );
  XNOR U26840 ( .A(n17768), .B(n17167), .Z(n17169) );
  XOR U26841 ( .A(n17769), .B(n17770), .Z(n17167) );
  ANDN U26842 ( .B(n17771), .A(n17772), .Z(n17769) );
  AND U26843 ( .A(a[56]), .B(b[45]), .Z(n17768) );
  XNOR U26844 ( .A(n17773), .B(n17172), .Z(n17174) );
  XOR U26845 ( .A(n17774), .B(n17775), .Z(n17172) );
  ANDN U26846 ( .B(n17776), .A(n17777), .Z(n17774) );
  AND U26847 ( .A(a[57]), .B(b[44]), .Z(n17773) );
  XNOR U26848 ( .A(n17778), .B(n17177), .Z(n17179) );
  XOR U26849 ( .A(n17779), .B(n17780), .Z(n17177) );
  ANDN U26850 ( .B(n17781), .A(n17782), .Z(n17779) );
  AND U26851 ( .A(a[58]), .B(b[43]), .Z(n17778) );
  XNOR U26852 ( .A(n17783), .B(n17182), .Z(n17184) );
  XOR U26853 ( .A(n17784), .B(n17785), .Z(n17182) );
  ANDN U26854 ( .B(n17786), .A(n17787), .Z(n17784) );
  AND U26855 ( .A(a[59]), .B(b[42]), .Z(n17783) );
  XNOR U26856 ( .A(n17788), .B(n17187), .Z(n17189) );
  XOR U26857 ( .A(n17789), .B(n17790), .Z(n17187) );
  ANDN U26858 ( .B(n17791), .A(n17792), .Z(n17789) );
  AND U26859 ( .A(a[60]), .B(b[41]), .Z(n17788) );
  XNOR U26860 ( .A(n17793), .B(n17192), .Z(n17194) );
  XOR U26861 ( .A(n17794), .B(n17795), .Z(n17192) );
  ANDN U26862 ( .B(n17796), .A(n17797), .Z(n17794) );
  AND U26863 ( .A(a[61]), .B(b[40]), .Z(n17793) );
  XNOR U26864 ( .A(n17798), .B(n17197), .Z(n17199) );
  XOR U26865 ( .A(n17799), .B(n17800), .Z(n17197) );
  ANDN U26866 ( .B(n17801), .A(n17802), .Z(n17799) );
  AND U26867 ( .A(a[62]), .B(b[39]), .Z(n17798) );
  XNOR U26868 ( .A(n17803), .B(n17202), .Z(n17204) );
  XOR U26869 ( .A(n17804), .B(n17805), .Z(n17202) );
  ANDN U26870 ( .B(n17806), .A(n17807), .Z(n17804) );
  AND U26871 ( .A(a[63]), .B(b[38]), .Z(n17803) );
  XNOR U26872 ( .A(n17808), .B(n17207), .Z(n17209) );
  XOR U26873 ( .A(n17809), .B(n17810), .Z(n17207) );
  ANDN U26874 ( .B(n17811), .A(n17812), .Z(n17809) );
  AND U26875 ( .A(a[64]), .B(b[37]), .Z(n17808) );
  XNOR U26876 ( .A(n17813), .B(n17212), .Z(n17214) );
  XOR U26877 ( .A(n17814), .B(n17815), .Z(n17212) );
  ANDN U26878 ( .B(n17816), .A(n17817), .Z(n17814) );
  AND U26879 ( .A(a[65]), .B(b[36]), .Z(n17813) );
  XNOR U26880 ( .A(n17818), .B(n17217), .Z(n17219) );
  XOR U26881 ( .A(n17819), .B(n17820), .Z(n17217) );
  ANDN U26882 ( .B(n17821), .A(n17822), .Z(n17819) );
  AND U26883 ( .A(a[66]), .B(b[35]), .Z(n17818) );
  XNOR U26884 ( .A(n17823), .B(n17222), .Z(n17224) );
  XOR U26885 ( .A(n17824), .B(n17825), .Z(n17222) );
  ANDN U26886 ( .B(n17826), .A(n17827), .Z(n17824) );
  AND U26887 ( .A(a[67]), .B(b[34]), .Z(n17823) );
  XNOR U26888 ( .A(n17828), .B(n17227), .Z(n17229) );
  XOR U26889 ( .A(n17829), .B(n17830), .Z(n17227) );
  ANDN U26890 ( .B(n17831), .A(n17832), .Z(n17829) );
  AND U26891 ( .A(a[68]), .B(b[33]), .Z(n17828) );
  XNOR U26892 ( .A(n17833), .B(n17232), .Z(n17234) );
  XOR U26893 ( .A(n17834), .B(n17835), .Z(n17232) );
  ANDN U26894 ( .B(n17836), .A(n17837), .Z(n17834) );
  AND U26895 ( .A(a[69]), .B(b[32]), .Z(n17833) );
  XNOR U26896 ( .A(n17838), .B(n17237), .Z(n17239) );
  XOR U26897 ( .A(n17839), .B(n17840), .Z(n17237) );
  ANDN U26898 ( .B(n17841), .A(n17842), .Z(n17839) );
  AND U26899 ( .A(a[70]), .B(b[31]), .Z(n17838) );
  XNOR U26900 ( .A(n17843), .B(n17242), .Z(n17244) );
  XOR U26901 ( .A(n17844), .B(n17845), .Z(n17242) );
  ANDN U26902 ( .B(n17846), .A(n17847), .Z(n17844) );
  AND U26903 ( .A(a[71]), .B(b[30]), .Z(n17843) );
  XNOR U26904 ( .A(n17848), .B(n17247), .Z(n17249) );
  XOR U26905 ( .A(n17849), .B(n17850), .Z(n17247) );
  ANDN U26906 ( .B(n17851), .A(n17852), .Z(n17849) );
  AND U26907 ( .A(a[72]), .B(b[29]), .Z(n17848) );
  XNOR U26908 ( .A(n17853), .B(n17252), .Z(n17254) );
  XOR U26909 ( .A(n17854), .B(n17855), .Z(n17252) );
  ANDN U26910 ( .B(n17856), .A(n17857), .Z(n17854) );
  AND U26911 ( .A(a[73]), .B(b[28]), .Z(n17853) );
  XNOR U26912 ( .A(n17858), .B(n17257), .Z(n17259) );
  XOR U26913 ( .A(n17859), .B(n17860), .Z(n17257) );
  ANDN U26914 ( .B(n17861), .A(n17862), .Z(n17859) );
  AND U26915 ( .A(a[74]), .B(b[27]), .Z(n17858) );
  XNOR U26916 ( .A(n17863), .B(n17262), .Z(n17264) );
  XOR U26917 ( .A(n17864), .B(n17865), .Z(n17262) );
  ANDN U26918 ( .B(n17866), .A(n17867), .Z(n17864) );
  AND U26919 ( .A(a[75]), .B(b[26]), .Z(n17863) );
  XNOR U26920 ( .A(n17868), .B(n17267), .Z(n17269) );
  XOR U26921 ( .A(n17869), .B(n17870), .Z(n17267) );
  ANDN U26922 ( .B(n17871), .A(n17872), .Z(n17869) );
  AND U26923 ( .A(a[76]), .B(b[25]), .Z(n17868) );
  XNOR U26924 ( .A(n17873), .B(n17272), .Z(n17274) );
  XOR U26925 ( .A(n17874), .B(n17875), .Z(n17272) );
  ANDN U26926 ( .B(n17876), .A(n17877), .Z(n17874) );
  AND U26927 ( .A(a[77]), .B(b[24]), .Z(n17873) );
  XNOR U26928 ( .A(n17878), .B(n17277), .Z(n17279) );
  XOR U26929 ( .A(n17879), .B(n17880), .Z(n17277) );
  ANDN U26930 ( .B(n17881), .A(n17882), .Z(n17879) );
  AND U26931 ( .A(a[78]), .B(b[23]), .Z(n17878) );
  XNOR U26932 ( .A(n17883), .B(n17282), .Z(n17284) );
  XOR U26933 ( .A(n17884), .B(n17885), .Z(n17282) );
  ANDN U26934 ( .B(n17886), .A(n17887), .Z(n17884) );
  AND U26935 ( .A(a[79]), .B(b[22]), .Z(n17883) );
  XNOR U26936 ( .A(n17888), .B(n17287), .Z(n17289) );
  XOR U26937 ( .A(n17889), .B(n17890), .Z(n17287) );
  ANDN U26938 ( .B(n17891), .A(n17892), .Z(n17889) );
  AND U26939 ( .A(a[80]), .B(b[21]), .Z(n17888) );
  XNOR U26940 ( .A(n17893), .B(n17292), .Z(n17294) );
  XOR U26941 ( .A(n17894), .B(n17895), .Z(n17292) );
  ANDN U26942 ( .B(n17896), .A(n17897), .Z(n17894) );
  AND U26943 ( .A(a[81]), .B(b[20]), .Z(n17893) );
  XNOR U26944 ( .A(n17898), .B(n17297), .Z(n17299) );
  XOR U26945 ( .A(n17899), .B(n17900), .Z(n17297) );
  ANDN U26946 ( .B(n17901), .A(n17902), .Z(n17899) );
  AND U26947 ( .A(a[82]), .B(b[19]), .Z(n17898) );
  XNOR U26948 ( .A(n17903), .B(n17302), .Z(n17304) );
  XOR U26949 ( .A(n17904), .B(n17905), .Z(n17302) );
  ANDN U26950 ( .B(n17906), .A(n17907), .Z(n17904) );
  AND U26951 ( .A(a[83]), .B(b[18]), .Z(n17903) );
  XNOR U26952 ( .A(n17908), .B(n17307), .Z(n17309) );
  XOR U26953 ( .A(n17909), .B(n17910), .Z(n17307) );
  ANDN U26954 ( .B(n17911), .A(n17912), .Z(n17909) );
  AND U26955 ( .A(a[84]), .B(b[17]), .Z(n17908) );
  XNOR U26956 ( .A(n17913), .B(n17312), .Z(n17314) );
  XOR U26957 ( .A(n17914), .B(n17915), .Z(n17312) );
  ANDN U26958 ( .B(n17916), .A(n17917), .Z(n17914) );
  AND U26959 ( .A(a[85]), .B(b[16]), .Z(n17913) );
  XNOR U26960 ( .A(n17918), .B(n17317), .Z(n17319) );
  XOR U26961 ( .A(n17919), .B(n17920), .Z(n17317) );
  ANDN U26962 ( .B(n17921), .A(n17922), .Z(n17919) );
  AND U26963 ( .A(a[86]), .B(b[15]), .Z(n17918) );
  XNOR U26964 ( .A(n17923), .B(n17322), .Z(n17324) );
  XOR U26965 ( .A(n17924), .B(n17925), .Z(n17322) );
  ANDN U26966 ( .B(n17926), .A(n17927), .Z(n17924) );
  AND U26967 ( .A(a[87]), .B(b[14]), .Z(n17923) );
  XNOR U26968 ( .A(n17928), .B(n17327), .Z(n17329) );
  XOR U26969 ( .A(n17929), .B(n17930), .Z(n17327) );
  ANDN U26970 ( .B(n17931), .A(n17932), .Z(n17929) );
  AND U26971 ( .A(a[88]), .B(b[13]), .Z(n17928) );
  XNOR U26972 ( .A(n17933), .B(n17332), .Z(n17334) );
  XOR U26973 ( .A(n17934), .B(n17935), .Z(n17332) );
  ANDN U26974 ( .B(n17936), .A(n17937), .Z(n17934) );
  AND U26975 ( .A(a[89]), .B(b[12]), .Z(n17933) );
  XNOR U26976 ( .A(n17938), .B(n17337), .Z(n17339) );
  XOR U26977 ( .A(n17939), .B(n17940), .Z(n17337) );
  ANDN U26978 ( .B(n17941), .A(n17942), .Z(n17939) );
  AND U26979 ( .A(a[90]), .B(b[11]), .Z(n17938) );
  XNOR U26980 ( .A(n17943), .B(n17342), .Z(n17344) );
  XOR U26981 ( .A(n17944), .B(n17945), .Z(n17342) );
  ANDN U26982 ( .B(n17946), .A(n17947), .Z(n17944) );
  AND U26983 ( .A(a[91]), .B(b[10]), .Z(n17943) );
  XNOR U26984 ( .A(n17948), .B(n17347), .Z(n17349) );
  XOR U26985 ( .A(n17949), .B(n17950), .Z(n17347) );
  ANDN U26986 ( .B(n17951), .A(n17952), .Z(n17949) );
  AND U26987 ( .A(b[9]), .B(a[92]), .Z(n17948) );
  XNOR U26988 ( .A(n17953), .B(n17352), .Z(n17354) );
  XOR U26989 ( .A(n17954), .B(n17955), .Z(n17352) );
  ANDN U26990 ( .B(n17956), .A(n17957), .Z(n17954) );
  AND U26991 ( .A(b[8]), .B(a[93]), .Z(n17953) );
  XNOR U26992 ( .A(n17958), .B(n17357), .Z(n17359) );
  XOR U26993 ( .A(n17959), .B(n17960), .Z(n17357) );
  ANDN U26994 ( .B(n17961), .A(n17962), .Z(n17959) );
  AND U26995 ( .A(b[7]), .B(a[94]), .Z(n17958) );
  XNOR U26996 ( .A(n17963), .B(n17362), .Z(n17364) );
  XOR U26997 ( .A(n17964), .B(n17965), .Z(n17362) );
  ANDN U26998 ( .B(n17966), .A(n17967), .Z(n17964) );
  AND U26999 ( .A(b[6]), .B(a[95]), .Z(n17963) );
  XNOR U27000 ( .A(n17968), .B(n17367), .Z(n17369) );
  XOR U27001 ( .A(n17969), .B(n17970), .Z(n17367) );
  ANDN U27002 ( .B(n17971), .A(n17972), .Z(n17969) );
  AND U27003 ( .A(b[5]), .B(a[96]), .Z(n17968) );
  XNOR U27004 ( .A(n17973), .B(n17372), .Z(n17374) );
  XOR U27005 ( .A(n17974), .B(n17975), .Z(n17372) );
  ANDN U27006 ( .B(n17976), .A(n17977), .Z(n17974) );
  AND U27007 ( .A(b[4]), .B(a[97]), .Z(n17973) );
  XNOR U27008 ( .A(n17978), .B(n17979), .Z(n17386) );
  NANDN U27009 ( .A(n17980), .B(n17981), .Z(n17979) );
  XNOR U27010 ( .A(n17982), .B(n17377), .Z(n17379) );
  XNOR U27011 ( .A(n17983), .B(n17984), .Z(n17377) );
  AND U27012 ( .A(n17985), .B(n17986), .Z(n17983) );
  AND U27013 ( .A(b[3]), .B(a[98]), .Z(n17982) );
  NAND U27014 ( .A(a[101]), .B(b[0]), .Z(n16788) );
  XNOR U27015 ( .A(n17392), .B(n17393), .Z(c[100]) );
  XNOR U27016 ( .A(n17980), .B(n17981), .Z(n17393) );
  XOR U27017 ( .A(n17978), .B(n17987), .Z(n17981) );
  NAND U27018 ( .A(b[1]), .B(a[99]), .Z(n17987) );
  XOR U27019 ( .A(n17986), .B(n17988), .Z(n17980) );
  XOR U27020 ( .A(n17978), .B(n17985), .Z(n17988) );
  XNOR U27021 ( .A(n17989), .B(n17984), .Z(n17985) );
  AND U27022 ( .A(b[2]), .B(a[98]), .Z(n17989) );
  OR U27023 ( .A(n3), .B(n4), .Z(n17978) );
  XOR U27024 ( .A(n17990), .B(n17991), .Z(n4) );
  NAND U27025 ( .A(a[99]), .B(b[0]), .Z(n3) );
  XOR U27026 ( .A(n17984), .B(n17976), .Z(n17992) );
  XNOR U27027 ( .A(n17975), .B(n17971), .Z(n17993) );
  XNOR U27028 ( .A(n17970), .B(n17966), .Z(n17994) );
  XNOR U27029 ( .A(n17965), .B(n17961), .Z(n17995) );
  XNOR U27030 ( .A(n17960), .B(n17956), .Z(n17996) );
  XNOR U27031 ( .A(n17955), .B(n17951), .Z(n17997) );
  XNOR U27032 ( .A(n17950), .B(n17946), .Z(n17998) );
  XNOR U27033 ( .A(n17945), .B(n17941), .Z(n17999) );
  XNOR U27034 ( .A(n17940), .B(n17936), .Z(n18000) );
  XNOR U27035 ( .A(n17935), .B(n17931), .Z(n18001) );
  XNOR U27036 ( .A(n17930), .B(n17926), .Z(n18002) );
  XNOR U27037 ( .A(n17925), .B(n17921), .Z(n18003) );
  XNOR U27038 ( .A(n17920), .B(n17916), .Z(n18004) );
  XNOR U27039 ( .A(n17915), .B(n17911), .Z(n18005) );
  XNOR U27040 ( .A(n17910), .B(n17906), .Z(n18006) );
  XNOR U27041 ( .A(n17905), .B(n17901), .Z(n18007) );
  XNOR U27042 ( .A(n17900), .B(n17896), .Z(n18008) );
  XNOR U27043 ( .A(n17895), .B(n17891), .Z(n18009) );
  XNOR U27044 ( .A(n17890), .B(n17886), .Z(n18010) );
  XNOR U27045 ( .A(n17885), .B(n17881), .Z(n18011) );
  XNOR U27046 ( .A(n17880), .B(n17876), .Z(n18012) );
  XNOR U27047 ( .A(n17875), .B(n17871), .Z(n18013) );
  XNOR U27048 ( .A(n17870), .B(n17866), .Z(n18014) );
  XNOR U27049 ( .A(n17865), .B(n17861), .Z(n18015) );
  XNOR U27050 ( .A(n17860), .B(n17856), .Z(n18016) );
  XNOR U27051 ( .A(n17855), .B(n17851), .Z(n18017) );
  XNOR U27052 ( .A(n17850), .B(n17846), .Z(n18018) );
  XNOR U27053 ( .A(n17845), .B(n17841), .Z(n18019) );
  XNOR U27054 ( .A(n17840), .B(n17836), .Z(n18020) );
  XNOR U27055 ( .A(n17835), .B(n17831), .Z(n18021) );
  XNOR U27056 ( .A(n17830), .B(n17826), .Z(n18022) );
  XNOR U27057 ( .A(n17825), .B(n17821), .Z(n18023) );
  XNOR U27058 ( .A(n17820), .B(n17816), .Z(n18024) );
  XNOR U27059 ( .A(n17815), .B(n17811), .Z(n18025) );
  XNOR U27060 ( .A(n17810), .B(n17806), .Z(n18026) );
  XNOR U27061 ( .A(n17805), .B(n17801), .Z(n18027) );
  XNOR U27062 ( .A(n17800), .B(n17796), .Z(n18028) );
  XNOR U27063 ( .A(n17795), .B(n17791), .Z(n18029) );
  XNOR U27064 ( .A(n17790), .B(n17786), .Z(n18030) );
  XNOR U27065 ( .A(n17785), .B(n17781), .Z(n18031) );
  XNOR U27066 ( .A(n17780), .B(n17776), .Z(n18032) );
  XNOR U27067 ( .A(n17775), .B(n17771), .Z(n18033) );
  XNOR U27068 ( .A(n17770), .B(n17766), .Z(n18034) );
  XNOR U27069 ( .A(n17765), .B(n17761), .Z(n18035) );
  XNOR U27070 ( .A(n17760), .B(n17756), .Z(n18036) );
  XNOR U27071 ( .A(n17755), .B(n17751), .Z(n18037) );
  XNOR U27072 ( .A(n17750), .B(n17746), .Z(n18038) );
  XNOR U27073 ( .A(n17745), .B(n17741), .Z(n18039) );
  XNOR U27074 ( .A(n17740), .B(n17736), .Z(n18040) );
  XNOR U27075 ( .A(n17735), .B(n17731), .Z(n18041) );
  XNOR U27076 ( .A(n17730), .B(n17726), .Z(n18042) );
  XNOR U27077 ( .A(n17725), .B(n17721), .Z(n18043) );
  XNOR U27078 ( .A(n17720), .B(n17716), .Z(n18044) );
  XNOR U27079 ( .A(n17715), .B(n17711), .Z(n18045) );
  XNOR U27080 ( .A(n17710), .B(n17706), .Z(n18046) );
  XNOR U27081 ( .A(n17705), .B(n17701), .Z(n18047) );
  XNOR U27082 ( .A(n17700), .B(n17696), .Z(n18048) );
  XNOR U27083 ( .A(n17695), .B(n17691), .Z(n18049) );
  XNOR U27084 ( .A(n17690), .B(n17686), .Z(n18050) );
  XNOR U27085 ( .A(n17685), .B(n17681), .Z(n18051) );
  XNOR U27086 ( .A(n17680), .B(n17676), .Z(n18052) );
  XNOR U27087 ( .A(n17675), .B(n17671), .Z(n18053) );
  XNOR U27088 ( .A(n17670), .B(n17666), .Z(n18054) );
  XNOR U27089 ( .A(n17665), .B(n17661), .Z(n18055) );
  XNOR U27090 ( .A(n17660), .B(n17656), .Z(n18056) );
  XNOR U27091 ( .A(n17655), .B(n17651), .Z(n18057) );
  XNOR U27092 ( .A(n17650), .B(n17646), .Z(n18058) );
  XNOR U27093 ( .A(n17645), .B(n17641), .Z(n18059) );
  XNOR U27094 ( .A(n17640), .B(n17636), .Z(n18060) );
  XNOR U27095 ( .A(n17635), .B(n17631), .Z(n18061) );
  XNOR U27096 ( .A(n17630), .B(n17626), .Z(n18062) );
  XNOR U27097 ( .A(n17625), .B(n17621), .Z(n18063) );
  XNOR U27098 ( .A(n17620), .B(n17616), .Z(n18064) );
  XNOR U27099 ( .A(n17615), .B(n17611), .Z(n18065) );
  XNOR U27100 ( .A(n17610), .B(n17606), .Z(n18066) );
  XNOR U27101 ( .A(n17605), .B(n17601), .Z(n18067) );
  XNOR U27102 ( .A(n17600), .B(n17596), .Z(n18068) );
  XNOR U27103 ( .A(n17595), .B(n17591), .Z(n18069) );
  XNOR U27104 ( .A(n17590), .B(n17586), .Z(n18070) );
  XNOR U27105 ( .A(n17585), .B(n17581), .Z(n18071) );
  XNOR U27106 ( .A(n17580), .B(n17576), .Z(n18072) );
  XNOR U27107 ( .A(n17575), .B(n17571), .Z(n18073) );
  XNOR U27108 ( .A(n17570), .B(n17566), .Z(n18074) );
  XNOR U27109 ( .A(n17565), .B(n17561), .Z(n18075) );
  XNOR U27110 ( .A(n17560), .B(n17556), .Z(n18076) );
  XNOR U27111 ( .A(n17555), .B(n17551), .Z(n18077) );
  XNOR U27112 ( .A(n17550), .B(n17546), .Z(n18078) );
  XNOR U27113 ( .A(n17545), .B(n17541), .Z(n18079) );
  XNOR U27114 ( .A(n17540), .B(n17536), .Z(n18080) );
  XNOR U27115 ( .A(n17535), .B(n17531), .Z(n18081) );
  XNOR U27116 ( .A(n17530), .B(n17526), .Z(n18082) );
  XNOR U27117 ( .A(n17525), .B(n17521), .Z(n18083) );
  XNOR U27118 ( .A(n17520), .B(n17516), .Z(n18084) );
  XNOR U27119 ( .A(n17515), .B(n17511), .Z(n18085) );
  XNOR U27120 ( .A(n17510), .B(n17506), .Z(n18086) );
  XNOR U27121 ( .A(n17505), .B(n17501), .Z(n18087) );
  XNOR U27122 ( .A(n17500), .B(n17496), .Z(n18088) );
  XOR U27123 ( .A(n18089), .B(n17495), .Z(n17496) );
  AND U27124 ( .A(a[0]), .B(b[100]), .Z(n18089) );
  XNOR U27125 ( .A(n18090), .B(n17495), .Z(n17497) );
  XNOR U27126 ( .A(n18091), .B(n18092), .Z(n17495) );
  ANDN U27127 ( .B(n18093), .A(n18094), .Z(n18091) );
  AND U27128 ( .A(a[1]), .B(b[99]), .Z(n18090) );
  XNOR U27129 ( .A(n18095), .B(n17500), .Z(n17502) );
  XNOR U27130 ( .A(n18096), .B(n18097), .Z(n17500) );
  ANDN U27131 ( .B(n18098), .A(n18099), .Z(n18096) );
  AND U27132 ( .A(a[2]), .B(b[98]), .Z(n18095) );
  XNOR U27133 ( .A(n18100), .B(n17505), .Z(n17507) );
  XNOR U27134 ( .A(n18101), .B(n18102), .Z(n17505) );
  ANDN U27135 ( .B(n18103), .A(n18104), .Z(n18101) );
  AND U27136 ( .A(a[3]), .B(b[97]), .Z(n18100) );
  XNOR U27137 ( .A(n18105), .B(n17510), .Z(n17512) );
  XNOR U27138 ( .A(n18106), .B(n18107), .Z(n17510) );
  ANDN U27139 ( .B(n18108), .A(n18109), .Z(n18106) );
  AND U27140 ( .A(a[4]), .B(b[96]), .Z(n18105) );
  XNOR U27141 ( .A(n18110), .B(n17515), .Z(n17517) );
  XNOR U27142 ( .A(n18111), .B(n18112), .Z(n17515) );
  ANDN U27143 ( .B(n18113), .A(n18114), .Z(n18111) );
  AND U27144 ( .A(a[5]), .B(b[95]), .Z(n18110) );
  XNOR U27145 ( .A(n18115), .B(n17520), .Z(n17522) );
  XNOR U27146 ( .A(n18116), .B(n18117), .Z(n17520) );
  ANDN U27147 ( .B(n18118), .A(n18119), .Z(n18116) );
  AND U27148 ( .A(a[6]), .B(b[94]), .Z(n18115) );
  XNOR U27149 ( .A(n18120), .B(n17525), .Z(n17527) );
  XNOR U27150 ( .A(n18121), .B(n18122), .Z(n17525) );
  ANDN U27151 ( .B(n18123), .A(n18124), .Z(n18121) );
  AND U27152 ( .A(a[7]), .B(b[93]), .Z(n18120) );
  XNOR U27153 ( .A(n18125), .B(n17530), .Z(n17532) );
  XNOR U27154 ( .A(n18126), .B(n18127), .Z(n17530) );
  ANDN U27155 ( .B(n18128), .A(n18129), .Z(n18126) );
  AND U27156 ( .A(a[8]), .B(b[92]), .Z(n18125) );
  XNOR U27157 ( .A(n18130), .B(n17535), .Z(n17537) );
  XNOR U27158 ( .A(n18131), .B(n18132), .Z(n17535) );
  ANDN U27159 ( .B(n18133), .A(n18134), .Z(n18131) );
  AND U27160 ( .A(a[9]), .B(b[91]), .Z(n18130) );
  XNOR U27161 ( .A(n18135), .B(n17540), .Z(n17542) );
  XNOR U27162 ( .A(n18136), .B(n18137), .Z(n17540) );
  ANDN U27163 ( .B(n18138), .A(n18139), .Z(n18136) );
  AND U27164 ( .A(a[10]), .B(b[90]), .Z(n18135) );
  XNOR U27165 ( .A(n18140), .B(n17545), .Z(n17547) );
  XNOR U27166 ( .A(n18141), .B(n18142), .Z(n17545) );
  ANDN U27167 ( .B(n18143), .A(n18144), .Z(n18141) );
  AND U27168 ( .A(a[11]), .B(b[89]), .Z(n18140) );
  XNOR U27169 ( .A(n18145), .B(n17550), .Z(n17552) );
  XNOR U27170 ( .A(n18146), .B(n18147), .Z(n17550) );
  ANDN U27171 ( .B(n18148), .A(n18149), .Z(n18146) );
  AND U27172 ( .A(a[12]), .B(b[88]), .Z(n18145) );
  XNOR U27173 ( .A(n18150), .B(n17555), .Z(n17557) );
  XNOR U27174 ( .A(n18151), .B(n18152), .Z(n17555) );
  ANDN U27175 ( .B(n18153), .A(n18154), .Z(n18151) );
  AND U27176 ( .A(a[13]), .B(b[87]), .Z(n18150) );
  XNOR U27177 ( .A(n18155), .B(n17560), .Z(n17562) );
  XNOR U27178 ( .A(n18156), .B(n18157), .Z(n17560) );
  ANDN U27179 ( .B(n18158), .A(n18159), .Z(n18156) );
  AND U27180 ( .A(a[14]), .B(b[86]), .Z(n18155) );
  XNOR U27181 ( .A(n18160), .B(n17565), .Z(n17567) );
  XNOR U27182 ( .A(n18161), .B(n18162), .Z(n17565) );
  ANDN U27183 ( .B(n18163), .A(n18164), .Z(n18161) );
  AND U27184 ( .A(a[15]), .B(b[85]), .Z(n18160) );
  XNOR U27185 ( .A(n18165), .B(n17570), .Z(n17572) );
  XNOR U27186 ( .A(n18166), .B(n18167), .Z(n17570) );
  ANDN U27187 ( .B(n18168), .A(n18169), .Z(n18166) );
  AND U27188 ( .A(a[16]), .B(b[84]), .Z(n18165) );
  XNOR U27189 ( .A(n18170), .B(n17575), .Z(n17577) );
  XNOR U27190 ( .A(n18171), .B(n18172), .Z(n17575) );
  ANDN U27191 ( .B(n18173), .A(n18174), .Z(n18171) );
  AND U27192 ( .A(a[17]), .B(b[83]), .Z(n18170) );
  XNOR U27193 ( .A(n18175), .B(n17580), .Z(n17582) );
  XNOR U27194 ( .A(n18176), .B(n18177), .Z(n17580) );
  ANDN U27195 ( .B(n18178), .A(n18179), .Z(n18176) );
  AND U27196 ( .A(a[18]), .B(b[82]), .Z(n18175) );
  XNOR U27197 ( .A(n18180), .B(n17585), .Z(n17587) );
  XNOR U27198 ( .A(n18181), .B(n18182), .Z(n17585) );
  ANDN U27199 ( .B(n18183), .A(n18184), .Z(n18181) );
  AND U27200 ( .A(a[19]), .B(b[81]), .Z(n18180) );
  XNOR U27201 ( .A(n18185), .B(n17590), .Z(n17592) );
  XNOR U27202 ( .A(n18186), .B(n18187), .Z(n17590) );
  ANDN U27203 ( .B(n18188), .A(n18189), .Z(n18186) );
  AND U27204 ( .A(a[20]), .B(b[80]), .Z(n18185) );
  XNOR U27205 ( .A(n18190), .B(n17595), .Z(n17597) );
  XNOR U27206 ( .A(n18191), .B(n18192), .Z(n17595) );
  ANDN U27207 ( .B(n18193), .A(n18194), .Z(n18191) );
  AND U27208 ( .A(a[21]), .B(b[79]), .Z(n18190) );
  XNOR U27209 ( .A(n18195), .B(n17600), .Z(n17602) );
  XNOR U27210 ( .A(n18196), .B(n18197), .Z(n17600) );
  ANDN U27211 ( .B(n18198), .A(n18199), .Z(n18196) );
  AND U27212 ( .A(a[22]), .B(b[78]), .Z(n18195) );
  XNOR U27213 ( .A(n18200), .B(n17605), .Z(n17607) );
  XNOR U27214 ( .A(n18201), .B(n18202), .Z(n17605) );
  ANDN U27215 ( .B(n18203), .A(n18204), .Z(n18201) );
  AND U27216 ( .A(a[23]), .B(b[77]), .Z(n18200) );
  XNOR U27217 ( .A(n18205), .B(n17610), .Z(n17612) );
  XNOR U27218 ( .A(n18206), .B(n18207), .Z(n17610) );
  ANDN U27219 ( .B(n18208), .A(n18209), .Z(n18206) );
  AND U27220 ( .A(a[24]), .B(b[76]), .Z(n18205) );
  XNOR U27221 ( .A(n18210), .B(n17615), .Z(n17617) );
  XNOR U27222 ( .A(n18211), .B(n18212), .Z(n17615) );
  ANDN U27223 ( .B(n18213), .A(n18214), .Z(n18211) );
  AND U27224 ( .A(a[25]), .B(b[75]), .Z(n18210) );
  XNOR U27225 ( .A(n18215), .B(n17620), .Z(n17622) );
  XNOR U27226 ( .A(n18216), .B(n18217), .Z(n17620) );
  ANDN U27227 ( .B(n18218), .A(n18219), .Z(n18216) );
  AND U27228 ( .A(a[26]), .B(b[74]), .Z(n18215) );
  XNOR U27229 ( .A(n18220), .B(n17625), .Z(n17627) );
  XNOR U27230 ( .A(n18221), .B(n18222), .Z(n17625) );
  ANDN U27231 ( .B(n18223), .A(n18224), .Z(n18221) );
  AND U27232 ( .A(a[27]), .B(b[73]), .Z(n18220) );
  XNOR U27233 ( .A(n18225), .B(n17630), .Z(n17632) );
  XNOR U27234 ( .A(n18226), .B(n18227), .Z(n17630) );
  ANDN U27235 ( .B(n18228), .A(n18229), .Z(n18226) );
  AND U27236 ( .A(a[28]), .B(b[72]), .Z(n18225) );
  XNOR U27237 ( .A(n18230), .B(n17635), .Z(n17637) );
  XNOR U27238 ( .A(n18231), .B(n18232), .Z(n17635) );
  ANDN U27239 ( .B(n18233), .A(n18234), .Z(n18231) );
  AND U27240 ( .A(a[29]), .B(b[71]), .Z(n18230) );
  XNOR U27241 ( .A(n18235), .B(n17640), .Z(n17642) );
  XNOR U27242 ( .A(n18236), .B(n18237), .Z(n17640) );
  ANDN U27243 ( .B(n18238), .A(n18239), .Z(n18236) );
  AND U27244 ( .A(a[30]), .B(b[70]), .Z(n18235) );
  XNOR U27245 ( .A(n18240), .B(n17645), .Z(n17647) );
  XNOR U27246 ( .A(n18241), .B(n18242), .Z(n17645) );
  ANDN U27247 ( .B(n18243), .A(n18244), .Z(n18241) );
  AND U27248 ( .A(a[31]), .B(b[69]), .Z(n18240) );
  XNOR U27249 ( .A(n18245), .B(n17650), .Z(n17652) );
  XNOR U27250 ( .A(n18246), .B(n18247), .Z(n17650) );
  ANDN U27251 ( .B(n18248), .A(n18249), .Z(n18246) );
  AND U27252 ( .A(a[32]), .B(b[68]), .Z(n18245) );
  XNOR U27253 ( .A(n18250), .B(n17655), .Z(n17657) );
  XNOR U27254 ( .A(n18251), .B(n18252), .Z(n17655) );
  ANDN U27255 ( .B(n18253), .A(n18254), .Z(n18251) );
  AND U27256 ( .A(a[33]), .B(b[67]), .Z(n18250) );
  XNOR U27257 ( .A(n18255), .B(n17660), .Z(n17662) );
  XNOR U27258 ( .A(n18256), .B(n18257), .Z(n17660) );
  ANDN U27259 ( .B(n18258), .A(n18259), .Z(n18256) );
  AND U27260 ( .A(a[34]), .B(b[66]), .Z(n18255) );
  XNOR U27261 ( .A(n18260), .B(n17665), .Z(n17667) );
  XNOR U27262 ( .A(n18261), .B(n18262), .Z(n17665) );
  ANDN U27263 ( .B(n18263), .A(n18264), .Z(n18261) );
  AND U27264 ( .A(a[35]), .B(b[65]), .Z(n18260) );
  XNOR U27265 ( .A(n18265), .B(n17670), .Z(n17672) );
  XNOR U27266 ( .A(n18266), .B(n18267), .Z(n17670) );
  ANDN U27267 ( .B(n18268), .A(n18269), .Z(n18266) );
  AND U27268 ( .A(a[36]), .B(b[64]), .Z(n18265) );
  XNOR U27269 ( .A(n18270), .B(n17675), .Z(n17677) );
  XNOR U27270 ( .A(n18271), .B(n18272), .Z(n17675) );
  ANDN U27271 ( .B(n18273), .A(n18274), .Z(n18271) );
  AND U27272 ( .A(a[37]), .B(b[63]), .Z(n18270) );
  XNOR U27273 ( .A(n18275), .B(n17680), .Z(n17682) );
  XNOR U27274 ( .A(n18276), .B(n18277), .Z(n17680) );
  ANDN U27275 ( .B(n18278), .A(n18279), .Z(n18276) );
  AND U27276 ( .A(a[38]), .B(b[62]), .Z(n18275) );
  XNOR U27277 ( .A(n18280), .B(n17685), .Z(n17687) );
  XNOR U27278 ( .A(n18281), .B(n18282), .Z(n17685) );
  ANDN U27279 ( .B(n18283), .A(n18284), .Z(n18281) );
  AND U27280 ( .A(a[39]), .B(b[61]), .Z(n18280) );
  XNOR U27281 ( .A(n18285), .B(n17690), .Z(n17692) );
  XNOR U27282 ( .A(n18286), .B(n18287), .Z(n17690) );
  ANDN U27283 ( .B(n18288), .A(n18289), .Z(n18286) );
  AND U27284 ( .A(a[40]), .B(b[60]), .Z(n18285) );
  XNOR U27285 ( .A(n18290), .B(n17695), .Z(n17697) );
  XNOR U27286 ( .A(n18291), .B(n18292), .Z(n17695) );
  ANDN U27287 ( .B(n18293), .A(n18294), .Z(n18291) );
  AND U27288 ( .A(a[41]), .B(b[59]), .Z(n18290) );
  XNOR U27289 ( .A(n18295), .B(n17700), .Z(n17702) );
  XNOR U27290 ( .A(n18296), .B(n18297), .Z(n17700) );
  ANDN U27291 ( .B(n18298), .A(n18299), .Z(n18296) );
  AND U27292 ( .A(a[42]), .B(b[58]), .Z(n18295) );
  XNOR U27293 ( .A(n18300), .B(n17705), .Z(n17707) );
  XNOR U27294 ( .A(n18301), .B(n18302), .Z(n17705) );
  ANDN U27295 ( .B(n18303), .A(n18304), .Z(n18301) );
  AND U27296 ( .A(a[43]), .B(b[57]), .Z(n18300) );
  XNOR U27297 ( .A(n18305), .B(n17710), .Z(n17712) );
  XNOR U27298 ( .A(n18306), .B(n18307), .Z(n17710) );
  ANDN U27299 ( .B(n18308), .A(n18309), .Z(n18306) );
  AND U27300 ( .A(a[44]), .B(b[56]), .Z(n18305) );
  XNOR U27301 ( .A(n18310), .B(n17715), .Z(n17717) );
  XNOR U27302 ( .A(n18311), .B(n18312), .Z(n17715) );
  ANDN U27303 ( .B(n18313), .A(n18314), .Z(n18311) );
  AND U27304 ( .A(a[45]), .B(b[55]), .Z(n18310) );
  XNOR U27305 ( .A(n18315), .B(n17720), .Z(n17722) );
  XNOR U27306 ( .A(n18316), .B(n18317), .Z(n17720) );
  ANDN U27307 ( .B(n18318), .A(n18319), .Z(n18316) );
  AND U27308 ( .A(a[46]), .B(b[54]), .Z(n18315) );
  XNOR U27309 ( .A(n18320), .B(n17725), .Z(n17727) );
  XNOR U27310 ( .A(n18321), .B(n18322), .Z(n17725) );
  ANDN U27311 ( .B(n18323), .A(n18324), .Z(n18321) );
  AND U27312 ( .A(a[47]), .B(b[53]), .Z(n18320) );
  XNOR U27313 ( .A(n18325), .B(n17730), .Z(n17732) );
  XNOR U27314 ( .A(n18326), .B(n18327), .Z(n17730) );
  ANDN U27315 ( .B(n18328), .A(n18329), .Z(n18326) );
  AND U27316 ( .A(a[48]), .B(b[52]), .Z(n18325) );
  XNOR U27317 ( .A(n18330), .B(n17735), .Z(n17737) );
  XNOR U27318 ( .A(n18331), .B(n18332), .Z(n17735) );
  ANDN U27319 ( .B(n18333), .A(n18334), .Z(n18331) );
  AND U27320 ( .A(a[49]), .B(b[51]), .Z(n18330) );
  XNOR U27321 ( .A(n18335), .B(n17740), .Z(n17742) );
  XNOR U27322 ( .A(n18336), .B(n18337), .Z(n17740) );
  ANDN U27323 ( .B(n18338), .A(n18339), .Z(n18336) );
  AND U27324 ( .A(a[50]), .B(b[50]), .Z(n18335) );
  XNOR U27325 ( .A(n18340), .B(n17745), .Z(n17747) );
  XNOR U27326 ( .A(n18341), .B(n18342), .Z(n17745) );
  ANDN U27327 ( .B(n18343), .A(n18344), .Z(n18341) );
  AND U27328 ( .A(a[51]), .B(b[49]), .Z(n18340) );
  XNOR U27329 ( .A(n18345), .B(n17750), .Z(n17752) );
  XNOR U27330 ( .A(n18346), .B(n18347), .Z(n17750) );
  ANDN U27331 ( .B(n18348), .A(n18349), .Z(n18346) );
  AND U27332 ( .A(a[52]), .B(b[48]), .Z(n18345) );
  XNOR U27333 ( .A(n18350), .B(n17755), .Z(n17757) );
  XNOR U27334 ( .A(n18351), .B(n18352), .Z(n17755) );
  ANDN U27335 ( .B(n18353), .A(n18354), .Z(n18351) );
  AND U27336 ( .A(a[53]), .B(b[47]), .Z(n18350) );
  XNOR U27337 ( .A(n18355), .B(n17760), .Z(n17762) );
  XNOR U27338 ( .A(n18356), .B(n18357), .Z(n17760) );
  ANDN U27339 ( .B(n18358), .A(n18359), .Z(n18356) );
  AND U27340 ( .A(a[54]), .B(b[46]), .Z(n18355) );
  XNOR U27341 ( .A(n18360), .B(n17765), .Z(n17767) );
  XNOR U27342 ( .A(n18361), .B(n18362), .Z(n17765) );
  ANDN U27343 ( .B(n18363), .A(n18364), .Z(n18361) );
  AND U27344 ( .A(a[55]), .B(b[45]), .Z(n18360) );
  XNOR U27345 ( .A(n18365), .B(n17770), .Z(n17772) );
  XNOR U27346 ( .A(n18366), .B(n18367), .Z(n17770) );
  ANDN U27347 ( .B(n18368), .A(n18369), .Z(n18366) );
  AND U27348 ( .A(a[56]), .B(b[44]), .Z(n18365) );
  XNOR U27349 ( .A(n18370), .B(n17775), .Z(n17777) );
  XNOR U27350 ( .A(n18371), .B(n18372), .Z(n17775) );
  ANDN U27351 ( .B(n18373), .A(n18374), .Z(n18371) );
  AND U27352 ( .A(a[57]), .B(b[43]), .Z(n18370) );
  XNOR U27353 ( .A(n18375), .B(n17780), .Z(n17782) );
  XNOR U27354 ( .A(n18376), .B(n18377), .Z(n17780) );
  ANDN U27355 ( .B(n18378), .A(n18379), .Z(n18376) );
  AND U27356 ( .A(a[58]), .B(b[42]), .Z(n18375) );
  XNOR U27357 ( .A(n18380), .B(n17785), .Z(n17787) );
  XNOR U27358 ( .A(n18381), .B(n18382), .Z(n17785) );
  ANDN U27359 ( .B(n18383), .A(n18384), .Z(n18381) );
  AND U27360 ( .A(a[59]), .B(b[41]), .Z(n18380) );
  XNOR U27361 ( .A(n18385), .B(n17790), .Z(n17792) );
  XNOR U27362 ( .A(n18386), .B(n18387), .Z(n17790) );
  ANDN U27363 ( .B(n18388), .A(n18389), .Z(n18386) );
  AND U27364 ( .A(a[60]), .B(b[40]), .Z(n18385) );
  XNOR U27365 ( .A(n18390), .B(n17795), .Z(n17797) );
  XNOR U27366 ( .A(n18391), .B(n18392), .Z(n17795) );
  ANDN U27367 ( .B(n18393), .A(n18394), .Z(n18391) );
  AND U27368 ( .A(a[61]), .B(b[39]), .Z(n18390) );
  XNOR U27369 ( .A(n18395), .B(n17800), .Z(n17802) );
  XNOR U27370 ( .A(n18396), .B(n18397), .Z(n17800) );
  ANDN U27371 ( .B(n18398), .A(n18399), .Z(n18396) );
  AND U27372 ( .A(a[62]), .B(b[38]), .Z(n18395) );
  XNOR U27373 ( .A(n18400), .B(n17805), .Z(n17807) );
  XNOR U27374 ( .A(n18401), .B(n18402), .Z(n17805) );
  ANDN U27375 ( .B(n18403), .A(n18404), .Z(n18401) );
  AND U27376 ( .A(a[63]), .B(b[37]), .Z(n18400) );
  XNOR U27377 ( .A(n18405), .B(n17810), .Z(n17812) );
  XNOR U27378 ( .A(n18406), .B(n18407), .Z(n17810) );
  ANDN U27379 ( .B(n18408), .A(n18409), .Z(n18406) );
  AND U27380 ( .A(a[64]), .B(b[36]), .Z(n18405) );
  XNOR U27381 ( .A(n18410), .B(n17815), .Z(n17817) );
  XNOR U27382 ( .A(n18411), .B(n18412), .Z(n17815) );
  ANDN U27383 ( .B(n18413), .A(n18414), .Z(n18411) );
  AND U27384 ( .A(a[65]), .B(b[35]), .Z(n18410) );
  XNOR U27385 ( .A(n18415), .B(n17820), .Z(n17822) );
  XNOR U27386 ( .A(n18416), .B(n18417), .Z(n17820) );
  ANDN U27387 ( .B(n18418), .A(n18419), .Z(n18416) );
  AND U27388 ( .A(a[66]), .B(b[34]), .Z(n18415) );
  XNOR U27389 ( .A(n18420), .B(n17825), .Z(n17827) );
  XNOR U27390 ( .A(n18421), .B(n18422), .Z(n17825) );
  ANDN U27391 ( .B(n18423), .A(n18424), .Z(n18421) );
  AND U27392 ( .A(a[67]), .B(b[33]), .Z(n18420) );
  XNOR U27393 ( .A(n18425), .B(n17830), .Z(n17832) );
  XNOR U27394 ( .A(n18426), .B(n18427), .Z(n17830) );
  ANDN U27395 ( .B(n18428), .A(n18429), .Z(n18426) );
  AND U27396 ( .A(a[68]), .B(b[32]), .Z(n18425) );
  XNOR U27397 ( .A(n18430), .B(n17835), .Z(n17837) );
  XNOR U27398 ( .A(n18431), .B(n18432), .Z(n17835) );
  ANDN U27399 ( .B(n18433), .A(n18434), .Z(n18431) );
  AND U27400 ( .A(a[69]), .B(b[31]), .Z(n18430) );
  XNOR U27401 ( .A(n18435), .B(n17840), .Z(n17842) );
  XNOR U27402 ( .A(n18436), .B(n18437), .Z(n17840) );
  ANDN U27403 ( .B(n18438), .A(n18439), .Z(n18436) );
  AND U27404 ( .A(a[70]), .B(b[30]), .Z(n18435) );
  XNOR U27405 ( .A(n18440), .B(n17845), .Z(n17847) );
  XNOR U27406 ( .A(n18441), .B(n18442), .Z(n17845) );
  ANDN U27407 ( .B(n18443), .A(n18444), .Z(n18441) );
  AND U27408 ( .A(a[71]), .B(b[29]), .Z(n18440) );
  XNOR U27409 ( .A(n18445), .B(n17850), .Z(n17852) );
  XNOR U27410 ( .A(n18446), .B(n18447), .Z(n17850) );
  ANDN U27411 ( .B(n18448), .A(n18449), .Z(n18446) );
  AND U27412 ( .A(a[72]), .B(b[28]), .Z(n18445) );
  XNOR U27413 ( .A(n18450), .B(n17855), .Z(n17857) );
  XNOR U27414 ( .A(n18451), .B(n18452), .Z(n17855) );
  ANDN U27415 ( .B(n18453), .A(n18454), .Z(n18451) );
  AND U27416 ( .A(a[73]), .B(b[27]), .Z(n18450) );
  XNOR U27417 ( .A(n18455), .B(n17860), .Z(n17862) );
  XNOR U27418 ( .A(n18456), .B(n18457), .Z(n17860) );
  ANDN U27419 ( .B(n18458), .A(n18459), .Z(n18456) );
  AND U27420 ( .A(a[74]), .B(b[26]), .Z(n18455) );
  XNOR U27421 ( .A(n18460), .B(n17865), .Z(n17867) );
  XNOR U27422 ( .A(n18461), .B(n18462), .Z(n17865) );
  ANDN U27423 ( .B(n18463), .A(n18464), .Z(n18461) );
  AND U27424 ( .A(a[75]), .B(b[25]), .Z(n18460) );
  XNOR U27425 ( .A(n18465), .B(n17870), .Z(n17872) );
  XNOR U27426 ( .A(n18466), .B(n18467), .Z(n17870) );
  ANDN U27427 ( .B(n18468), .A(n18469), .Z(n18466) );
  AND U27428 ( .A(a[76]), .B(b[24]), .Z(n18465) );
  XNOR U27429 ( .A(n18470), .B(n17875), .Z(n17877) );
  XNOR U27430 ( .A(n18471), .B(n18472), .Z(n17875) );
  ANDN U27431 ( .B(n18473), .A(n18474), .Z(n18471) );
  AND U27432 ( .A(a[77]), .B(b[23]), .Z(n18470) );
  XNOR U27433 ( .A(n18475), .B(n17880), .Z(n17882) );
  XNOR U27434 ( .A(n18476), .B(n18477), .Z(n17880) );
  ANDN U27435 ( .B(n18478), .A(n18479), .Z(n18476) );
  AND U27436 ( .A(a[78]), .B(b[22]), .Z(n18475) );
  XNOR U27437 ( .A(n18480), .B(n17885), .Z(n17887) );
  XNOR U27438 ( .A(n18481), .B(n18482), .Z(n17885) );
  ANDN U27439 ( .B(n18483), .A(n18484), .Z(n18481) );
  AND U27440 ( .A(a[79]), .B(b[21]), .Z(n18480) );
  XNOR U27441 ( .A(n18485), .B(n17890), .Z(n17892) );
  XNOR U27442 ( .A(n18486), .B(n18487), .Z(n17890) );
  ANDN U27443 ( .B(n18488), .A(n18489), .Z(n18486) );
  AND U27444 ( .A(a[80]), .B(b[20]), .Z(n18485) );
  XNOR U27445 ( .A(n18490), .B(n17895), .Z(n17897) );
  XNOR U27446 ( .A(n18491), .B(n18492), .Z(n17895) );
  ANDN U27447 ( .B(n18493), .A(n18494), .Z(n18491) );
  AND U27448 ( .A(a[81]), .B(b[19]), .Z(n18490) );
  XNOR U27449 ( .A(n18495), .B(n17900), .Z(n17902) );
  XNOR U27450 ( .A(n18496), .B(n18497), .Z(n17900) );
  ANDN U27451 ( .B(n18498), .A(n18499), .Z(n18496) );
  AND U27452 ( .A(a[82]), .B(b[18]), .Z(n18495) );
  XNOR U27453 ( .A(n18500), .B(n17905), .Z(n17907) );
  XNOR U27454 ( .A(n18501), .B(n18502), .Z(n17905) );
  ANDN U27455 ( .B(n18503), .A(n18504), .Z(n18501) );
  AND U27456 ( .A(a[83]), .B(b[17]), .Z(n18500) );
  XNOR U27457 ( .A(n18505), .B(n17910), .Z(n17912) );
  XNOR U27458 ( .A(n18506), .B(n18507), .Z(n17910) );
  ANDN U27459 ( .B(n18508), .A(n18509), .Z(n18506) );
  AND U27460 ( .A(a[84]), .B(b[16]), .Z(n18505) );
  XNOR U27461 ( .A(n18510), .B(n17915), .Z(n17917) );
  XNOR U27462 ( .A(n18511), .B(n18512), .Z(n17915) );
  ANDN U27463 ( .B(n18513), .A(n18514), .Z(n18511) );
  AND U27464 ( .A(a[85]), .B(b[15]), .Z(n18510) );
  XNOR U27465 ( .A(n18515), .B(n17920), .Z(n17922) );
  XNOR U27466 ( .A(n18516), .B(n18517), .Z(n17920) );
  ANDN U27467 ( .B(n18518), .A(n18519), .Z(n18516) );
  AND U27468 ( .A(a[86]), .B(b[14]), .Z(n18515) );
  XNOR U27469 ( .A(n18520), .B(n17925), .Z(n17927) );
  XNOR U27470 ( .A(n18521), .B(n18522), .Z(n17925) );
  ANDN U27471 ( .B(n18523), .A(n18524), .Z(n18521) );
  AND U27472 ( .A(a[87]), .B(b[13]), .Z(n18520) );
  XNOR U27473 ( .A(n18525), .B(n17930), .Z(n17932) );
  XNOR U27474 ( .A(n18526), .B(n18527), .Z(n17930) );
  ANDN U27475 ( .B(n18528), .A(n18529), .Z(n18526) );
  AND U27476 ( .A(a[88]), .B(b[12]), .Z(n18525) );
  XNOR U27477 ( .A(n18530), .B(n17935), .Z(n17937) );
  XNOR U27478 ( .A(n18531), .B(n18532), .Z(n17935) );
  ANDN U27479 ( .B(n18533), .A(n18534), .Z(n18531) );
  AND U27480 ( .A(a[89]), .B(b[11]), .Z(n18530) );
  XNOR U27481 ( .A(n18535), .B(n17940), .Z(n17942) );
  XNOR U27482 ( .A(n18536), .B(n18537), .Z(n17940) );
  ANDN U27483 ( .B(n18538), .A(n18539), .Z(n18536) );
  AND U27484 ( .A(a[90]), .B(b[10]), .Z(n18535) );
  XNOR U27485 ( .A(n18540), .B(n17945), .Z(n17947) );
  XNOR U27486 ( .A(n18541), .B(n18542), .Z(n17945) );
  ANDN U27487 ( .B(n18543), .A(n18544), .Z(n18541) );
  AND U27488 ( .A(b[9]), .B(a[91]), .Z(n18540) );
  XNOR U27489 ( .A(n18545), .B(n17950), .Z(n17952) );
  XNOR U27490 ( .A(n18546), .B(n18547), .Z(n17950) );
  ANDN U27491 ( .B(n18548), .A(n18549), .Z(n18546) );
  AND U27492 ( .A(b[8]), .B(a[92]), .Z(n18545) );
  XNOR U27493 ( .A(n18550), .B(n17955), .Z(n17957) );
  XNOR U27494 ( .A(n18551), .B(n18552), .Z(n17955) );
  ANDN U27495 ( .B(n18553), .A(n18554), .Z(n18551) );
  AND U27496 ( .A(b[7]), .B(a[93]), .Z(n18550) );
  XNOR U27497 ( .A(n18555), .B(n17960), .Z(n17962) );
  XNOR U27498 ( .A(n18556), .B(n18557), .Z(n17960) );
  ANDN U27499 ( .B(n18558), .A(n18559), .Z(n18556) );
  AND U27500 ( .A(b[6]), .B(a[94]), .Z(n18555) );
  XNOR U27501 ( .A(n18560), .B(n17965), .Z(n17967) );
  XNOR U27502 ( .A(n18561), .B(n18562), .Z(n17965) );
  ANDN U27503 ( .B(n18563), .A(n18564), .Z(n18561) );
  AND U27504 ( .A(b[5]), .B(a[95]), .Z(n18560) );
  XNOR U27505 ( .A(n18565), .B(n17970), .Z(n17972) );
  XNOR U27506 ( .A(n18566), .B(n18567), .Z(n17970) );
  ANDN U27507 ( .B(n18568), .A(n18569), .Z(n18566) );
  AND U27508 ( .A(b[4]), .B(a[96]), .Z(n18565) );
  XNOR U27509 ( .A(n18570), .B(n18571), .Z(n17984) );
  NANDN U27510 ( .A(n17991), .B(n17990), .Z(n18571) );
  XOR U27511 ( .A(n18570), .B(n18572), .Z(n17990) );
  NAND U27512 ( .A(b[1]), .B(a[98]), .Z(n18572) );
  XOR U27513 ( .A(n18570), .B(n18574), .Z(n18573) );
  NANDN U27514 ( .A(n5), .B(n6), .Z(n18570) );
  XOR U27515 ( .A(n18576), .B(n18577), .Z(n6) );
  NAND U27516 ( .A(a[98]), .B(b[0]), .Z(n5) );
  XNOR U27517 ( .A(n18578), .B(n17975), .Z(n17977) );
  XNOR U27518 ( .A(n18579), .B(n18580), .Z(n17975) );
  ANDN U27519 ( .B(n18574), .A(n18575), .Z(n18579) );
  XOR U27520 ( .A(n18581), .B(n18580), .Z(n18575) );
  IV U27521 ( .A(n18582), .Z(n18580) );
  AND U27522 ( .A(b[2]), .B(a[97]), .Z(n18581) );
  XNOR U27523 ( .A(n18568), .B(n18582), .Z(n18583) );
  XOR U27524 ( .A(n18584), .B(n18585), .Z(n18582) );
  OR U27525 ( .A(n18576), .B(n18577), .Z(n18585) );
  XNOR U27526 ( .A(n18587), .B(n18588), .Z(n18586) );
  XOR U27527 ( .A(n18587), .B(n18590), .Z(n18576) );
  NAND U27528 ( .A(b[1]), .B(a[97]), .Z(n18590) );
  IV U27529 ( .A(n18584), .Z(n18587) );
  NANDN U27530 ( .A(n7), .B(n8), .Z(n18584) );
  XOR U27531 ( .A(n18591), .B(n18592), .Z(n8) );
  NAND U27532 ( .A(a[97]), .B(b[0]), .Z(n7) );
  XNOR U27533 ( .A(n18563), .B(n18594), .Z(n18593) );
  XNOR U27534 ( .A(n18558), .B(n18596), .Z(n18595) );
  XNOR U27535 ( .A(n18553), .B(n18598), .Z(n18597) );
  XNOR U27536 ( .A(n18548), .B(n18600), .Z(n18599) );
  XNOR U27537 ( .A(n18543), .B(n18602), .Z(n18601) );
  XNOR U27538 ( .A(n18538), .B(n18604), .Z(n18603) );
  XNOR U27539 ( .A(n18533), .B(n18606), .Z(n18605) );
  XNOR U27540 ( .A(n18528), .B(n18608), .Z(n18607) );
  XNOR U27541 ( .A(n18523), .B(n18610), .Z(n18609) );
  XNOR U27542 ( .A(n18518), .B(n18612), .Z(n18611) );
  XNOR U27543 ( .A(n18513), .B(n18614), .Z(n18613) );
  XNOR U27544 ( .A(n18508), .B(n18616), .Z(n18615) );
  XNOR U27545 ( .A(n18503), .B(n18618), .Z(n18617) );
  XNOR U27546 ( .A(n18498), .B(n18620), .Z(n18619) );
  XNOR U27547 ( .A(n18493), .B(n18622), .Z(n18621) );
  XNOR U27548 ( .A(n18488), .B(n18624), .Z(n18623) );
  XNOR U27549 ( .A(n18483), .B(n18626), .Z(n18625) );
  XNOR U27550 ( .A(n18478), .B(n18628), .Z(n18627) );
  XNOR U27551 ( .A(n18473), .B(n18630), .Z(n18629) );
  XNOR U27552 ( .A(n18468), .B(n18632), .Z(n18631) );
  XNOR U27553 ( .A(n18463), .B(n18634), .Z(n18633) );
  XNOR U27554 ( .A(n18458), .B(n18636), .Z(n18635) );
  XNOR U27555 ( .A(n18453), .B(n18638), .Z(n18637) );
  XNOR U27556 ( .A(n18448), .B(n18640), .Z(n18639) );
  XNOR U27557 ( .A(n18443), .B(n18642), .Z(n18641) );
  XNOR U27558 ( .A(n18438), .B(n18644), .Z(n18643) );
  XNOR U27559 ( .A(n18433), .B(n18646), .Z(n18645) );
  XNOR U27560 ( .A(n18428), .B(n18648), .Z(n18647) );
  XNOR U27561 ( .A(n18423), .B(n18650), .Z(n18649) );
  XNOR U27562 ( .A(n18418), .B(n18652), .Z(n18651) );
  XNOR U27563 ( .A(n18413), .B(n18654), .Z(n18653) );
  XNOR U27564 ( .A(n18408), .B(n18656), .Z(n18655) );
  XNOR U27565 ( .A(n18403), .B(n18658), .Z(n18657) );
  XNOR U27566 ( .A(n18398), .B(n18660), .Z(n18659) );
  XNOR U27567 ( .A(n18393), .B(n18662), .Z(n18661) );
  XNOR U27568 ( .A(n18388), .B(n18664), .Z(n18663) );
  XNOR U27569 ( .A(n18383), .B(n18666), .Z(n18665) );
  XNOR U27570 ( .A(n18378), .B(n18668), .Z(n18667) );
  XNOR U27571 ( .A(n18373), .B(n18670), .Z(n18669) );
  XNOR U27572 ( .A(n18368), .B(n18672), .Z(n18671) );
  XNOR U27573 ( .A(n18363), .B(n18674), .Z(n18673) );
  XNOR U27574 ( .A(n18358), .B(n18676), .Z(n18675) );
  XNOR U27575 ( .A(n18353), .B(n18678), .Z(n18677) );
  XNOR U27576 ( .A(n18348), .B(n18680), .Z(n18679) );
  XNOR U27577 ( .A(n18343), .B(n18682), .Z(n18681) );
  XNOR U27578 ( .A(n18338), .B(n18684), .Z(n18683) );
  XNOR U27579 ( .A(n18333), .B(n18686), .Z(n18685) );
  XNOR U27580 ( .A(n18328), .B(n18688), .Z(n18687) );
  XNOR U27581 ( .A(n18323), .B(n18690), .Z(n18689) );
  XNOR U27582 ( .A(n18318), .B(n18692), .Z(n18691) );
  XNOR U27583 ( .A(n18313), .B(n18694), .Z(n18693) );
  XNOR U27584 ( .A(n18308), .B(n18696), .Z(n18695) );
  XNOR U27585 ( .A(n18303), .B(n18698), .Z(n18697) );
  XNOR U27586 ( .A(n18298), .B(n18700), .Z(n18699) );
  XNOR U27587 ( .A(n18293), .B(n18702), .Z(n18701) );
  XNOR U27588 ( .A(n18288), .B(n18704), .Z(n18703) );
  XNOR U27589 ( .A(n18283), .B(n18706), .Z(n18705) );
  XNOR U27590 ( .A(n18278), .B(n18708), .Z(n18707) );
  XNOR U27591 ( .A(n18273), .B(n18710), .Z(n18709) );
  XNOR U27592 ( .A(n18268), .B(n18712), .Z(n18711) );
  XNOR U27593 ( .A(n18263), .B(n18714), .Z(n18713) );
  XNOR U27594 ( .A(n18258), .B(n18716), .Z(n18715) );
  XNOR U27595 ( .A(n18253), .B(n18718), .Z(n18717) );
  XNOR U27596 ( .A(n18248), .B(n18720), .Z(n18719) );
  XNOR U27597 ( .A(n18243), .B(n18722), .Z(n18721) );
  XNOR U27598 ( .A(n18238), .B(n18724), .Z(n18723) );
  XNOR U27599 ( .A(n18233), .B(n18726), .Z(n18725) );
  XNOR U27600 ( .A(n18228), .B(n18728), .Z(n18727) );
  XNOR U27601 ( .A(n18223), .B(n18730), .Z(n18729) );
  XNOR U27602 ( .A(n18218), .B(n18732), .Z(n18731) );
  XNOR U27603 ( .A(n18213), .B(n18734), .Z(n18733) );
  XNOR U27604 ( .A(n18208), .B(n18736), .Z(n18735) );
  XNOR U27605 ( .A(n18203), .B(n18738), .Z(n18737) );
  XNOR U27606 ( .A(n18198), .B(n18740), .Z(n18739) );
  XNOR U27607 ( .A(n18193), .B(n18742), .Z(n18741) );
  XNOR U27608 ( .A(n18188), .B(n18744), .Z(n18743) );
  XNOR U27609 ( .A(n18183), .B(n18746), .Z(n18745) );
  XNOR U27610 ( .A(n18178), .B(n18748), .Z(n18747) );
  XNOR U27611 ( .A(n18173), .B(n18750), .Z(n18749) );
  XNOR U27612 ( .A(n18168), .B(n18752), .Z(n18751) );
  XNOR U27613 ( .A(n18163), .B(n18754), .Z(n18753) );
  XNOR U27614 ( .A(n18158), .B(n18756), .Z(n18755) );
  XNOR U27615 ( .A(n18153), .B(n18758), .Z(n18757) );
  XNOR U27616 ( .A(n18148), .B(n18760), .Z(n18759) );
  XNOR U27617 ( .A(n18143), .B(n18762), .Z(n18761) );
  XNOR U27618 ( .A(n18138), .B(n18764), .Z(n18763) );
  XNOR U27619 ( .A(n18133), .B(n18766), .Z(n18765) );
  XNOR U27620 ( .A(n18128), .B(n18768), .Z(n18767) );
  XNOR U27621 ( .A(n18123), .B(n18770), .Z(n18769) );
  XNOR U27622 ( .A(n18118), .B(n18772), .Z(n18771) );
  XNOR U27623 ( .A(n18113), .B(n18774), .Z(n18773) );
  XNOR U27624 ( .A(n18108), .B(n18776), .Z(n18775) );
  XNOR U27625 ( .A(n18103), .B(n18778), .Z(n18777) );
  XNOR U27626 ( .A(n18098), .B(n18780), .Z(n18779) );
  XNOR U27627 ( .A(n18093), .B(n18782), .Z(n18781) );
  XNOR U27628 ( .A(n18783), .B(n18092), .Z(n18093) );
  AND U27629 ( .A(a[0]), .B(b[99]), .Z(n18783) );
  XOR U27630 ( .A(n18784), .B(n18092), .Z(n18094) );
  XNOR U27631 ( .A(n18785), .B(n18786), .Z(n18092) );
  ANDN U27632 ( .B(n18787), .A(n18788), .Z(n18785) );
  AND U27633 ( .A(a[1]), .B(b[98]), .Z(n18784) );
  XOR U27634 ( .A(n18789), .B(n18097), .Z(n18099) );
  IV U27635 ( .A(n18782), .Z(n18097) );
  XOR U27636 ( .A(n18790), .B(n18791), .Z(n18782) );
  ANDN U27637 ( .B(n18792), .A(n18793), .Z(n18790) );
  AND U27638 ( .A(a[2]), .B(b[97]), .Z(n18789) );
  XOR U27639 ( .A(n18794), .B(n18102), .Z(n18104) );
  IV U27640 ( .A(n18780), .Z(n18102) );
  XOR U27641 ( .A(n18795), .B(n18796), .Z(n18780) );
  ANDN U27642 ( .B(n18797), .A(n18798), .Z(n18795) );
  AND U27643 ( .A(a[3]), .B(b[96]), .Z(n18794) );
  XOR U27644 ( .A(n18799), .B(n18107), .Z(n18109) );
  IV U27645 ( .A(n18778), .Z(n18107) );
  XOR U27646 ( .A(n18800), .B(n18801), .Z(n18778) );
  ANDN U27647 ( .B(n18802), .A(n18803), .Z(n18800) );
  AND U27648 ( .A(a[4]), .B(b[95]), .Z(n18799) );
  XOR U27649 ( .A(n18804), .B(n18112), .Z(n18114) );
  IV U27650 ( .A(n18776), .Z(n18112) );
  XOR U27651 ( .A(n18805), .B(n18806), .Z(n18776) );
  ANDN U27652 ( .B(n18807), .A(n18808), .Z(n18805) );
  AND U27653 ( .A(a[5]), .B(b[94]), .Z(n18804) );
  XOR U27654 ( .A(n18809), .B(n18117), .Z(n18119) );
  IV U27655 ( .A(n18774), .Z(n18117) );
  XOR U27656 ( .A(n18810), .B(n18811), .Z(n18774) );
  ANDN U27657 ( .B(n18812), .A(n18813), .Z(n18810) );
  AND U27658 ( .A(a[6]), .B(b[93]), .Z(n18809) );
  XOR U27659 ( .A(n18814), .B(n18122), .Z(n18124) );
  IV U27660 ( .A(n18772), .Z(n18122) );
  XOR U27661 ( .A(n18815), .B(n18816), .Z(n18772) );
  ANDN U27662 ( .B(n18817), .A(n18818), .Z(n18815) );
  AND U27663 ( .A(a[7]), .B(b[92]), .Z(n18814) );
  XOR U27664 ( .A(n18819), .B(n18127), .Z(n18129) );
  IV U27665 ( .A(n18770), .Z(n18127) );
  XOR U27666 ( .A(n18820), .B(n18821), .Z(n18770) );
  ANDN U27667 ( .B(n18822), .A(n18823), .Z(n18820) );
  AND U27668 ( .A(a[8]), .B(b[91]), .Z(n18819) );
  XOR U27669 ( .A(n18824), .B(n18132), .Z(n18134) );
  IV U27670 ( .A(n18768), .Z(n18132) );
  XOR U27671 ( .A(n18825), .B(n18826), .Z(n18768) );
  ANDN U27672 ( .B(n18827), .A(n18828), .Z(n18825) );
  AND U27673 ( .A(a[9]), .B(b[90]), .Z(n18824) );
  XOR U27674 ( .A(n18829), .B(n18137), .Z(n18139) );
  IV U27675 ( .A(n18766), .Z(n18137) );
  XOR U27676 ( .A(n18830), .B(n18831), .Z(n18766) );
  ANDN U27677 ( .B(n18832), .A(n18833), .Z(n18830) );
  AND U27678 ( .A(a[10]), .B(b[89]), .Z(n18829) );
  XOR U27679 ( .A(n18834), .B(n18142), .Z(n18144) );
  IV U27680 ( .A(n18764), .Z(n18142) );
  XOR U27681 ( .A(n18835), .B(n18836), .Z(n18764) );
  ANDN U27682 ( .B(n18837), .A(n18838), .Z(n18835) );
  AND U27683 ( .A(a[11]), .B(b[88]), .Z(n18834) );
  XOR U27684 ( .A(n18839), .B(n18147), .Z(n18149) );
  IV U27685 ( .A(n18762), .Z(n18147) );
  XOR U27686 ( .A(n18840), .B(n18841), .Z(n18762) );
  ANDN U27687 ( .B(n18842), .A(n18843), .Z(n18840) );
  AND U27688 ( .A(a[12]), .B(b[87]), .Z(n18839) );
  XOR U27689 ( .A(n18844), .B(n18152), .Z(n18154) );
  IV U27690 ( .A(n18760), .Z(n18152) );
  XOR U27691 ( .A(n18845), .B(n18846), .Z(n18760) );
  ANDN U27692 ( .B(n18847), .A(n18848), .Z(n18845) );
  AND U27693 ( .A(a[13]), .B(b[86]), .Z(n18844) );
  XOR U27694 ( .A(n18849), .B(n18157), .Z(n18159) );
  IV U27695 ( .A(n18758), .Z(n18157) );
  XOR U27696 ( .A(n18850), .B(n18851), .Z(n18758) );
  ANDN U27697 ( .B(n18852), .A(n18853), .Z(n18850) );
  AND U27698 ( .A(a[14]), .B(b[85]), .Z(n18849) );
  XOR U27699 ( .A(n18854), .B(n18162), .Z(n18164) );
  IV U27700 ( .A(n18756), .Z(n18162) );
  XOR U27701 ( .A(n18855), .B(n18856), .Z(n18756) );
  ANDN U27702 ( .B(n18857), .A(n18858), .Z(n18855) );
  AND U27703 ( .A(a[15]), .B(b[84]), .Z(n18854) );
  XOR U27704 ( .A(n18859), .B(n18167), .Z(n18169) );
  IV U27705 ( .A(n18754), .Z(n18167) );
  XOR U27706 ( .A(n18860), .B(n18861), .Z(n18754) );
  ANDN U27707 ( .B(n18862), .A(n18863), .Z(n18860) );
  AND U27708 ( .A(a[16]), .B(b[83]), .Z(n18859) );
  XOR U27709 ( .A(n18864), .B(n18172), .Z(n18174) );
  IV U27710 ( .A(n18752), .Z(n18172) );
  XOR U27711 ( .A(n18865), .B(n18866), .Z(n18752) );
  ANDN U27712 ( .B(n18867), .A(n18868), .Z(n18865) );
  AND U27713 ( .A(a[17]), .B(b[82]), .Z(n18864) );
  XOR U27714 ( .A(n18869), .B(n18177), .Z(n18179) );
  IV U27715 ( .A(n18750), .Z(n18177) );
  XOR U27716 ( .A(n18870), .B(n18871), .Z(n18750) );
  ANDN U27717 ( .B(n18872), .A(n18873), .Z(n18870) );
  AND U27718 ( .A(a[18]), .B(b[81]), .Z(n18869) );
  XOR U27719 ( .A(n18874), .B(n18182), .Z(n18184) );
  IV U27720 ( .A(n18748), .Z(n18182) );
  XOR U27721 ( .A(n18875), .B(n18876), .Z(n18748) );
  ANDN U27722 ( .B(n18877), .A(n18878), .Z(n18875) );
  AND U27723 ( .A(a[19]), .B(b[80]), .Z(n18874) );
  XOR U27724 ( .A(n18879), .B(n18187), .Z(n18189) );
  IV U27725 ( .A(n18746), .Z(n18187) );
  XOR U27726 ( .A(n18880), .B(n18881), .Z(n18746) );
  ANDN U27727 ( .B(n18882), .A(n18883), .Z(n18880) );
  AND U27728 ( .A(a[20]), .B(b[79]), .Z(n18879) );
  XOR U27729 ( .A(n18884), .B(n18192), .Z(n18194) );
  IV U27730 ( .A(n18744), .Z(n18192) );
  XOR U27731 ( .A(n18885), .B(n18886), .Z(n18744) );
  ANDN U27732 ( .B(n18887), .A(n18888), .Z(n18885) );
  AND U27733 ( .A(a[21]), .B(b[78]), .Z(n18884) );
  XOR U27734 ( .A(n18889), .B(n18197), .Z(n18199) );
  IV U27735 ( .A(n18742), .Z(n18197) );
  XOR U27736 ( .A(n18890), .B(n18891), .Z(n18742) );
  ANDN U27737 ( .B(n18892), .A(n18893), .Z(n18890) );
  AND U27738 ( .A(a[22]), .B(b[77]), .Z(n18889) );
  XOR U27739 ( .A(n18894), .B(n18202), .Z(n18204) );
  IV U27740 ( .A(n18740), .Z(n18202) );
  XOR U27741 ( .A(n18895), .B(n18896), .Z(n18740) );
  ANDN U27742 ( .B(n18897), .A(n18898), .Z(n18895) );
  AND U27743 ( .A(a[23]), .B(b[76]), .Z(n18894) );
  XOR U27744 ( .A(n18899), .B(n18207), .Z(n18209) );
  IV U27745 ( .A(n18738), .Z(n18207) );
  XOR U27746 ( .A(n18900), .B(n18901), .Z(n18738) );
  ANDN U27747 ( .B(n18902), .A(n18903), .Z(n18900) );
  AND U27748 ( .A(a[24]), .B(b[75]), .Z(n18899) );
  XOR U27749 ( .A(n18904), .B(n18212), .Z(n18214) );
  IV U27750 ( .A(n18736), .Z(n18212) );
  XOR U27751 ( .A(n18905), .B(n18906), .Z(n18736) );
  ANDN U27752 ( .B(n18907), .A(n18908), .Z(n18905) );
  AND U27753 ( .A(a[25]), .B(b[74]), .Z(n18904) );
  XOR U27754 ( .A(n18909), .B(n18217), .Z(n18219) );
  IV U27755 ( .A(n18734), .Z(n18217) );
  XOR U27756 ( .A(n18910), .B(n18911), .Z(n18734) );
  ANDN U27757 ( .B(n18912), .A(n18913), .Z(n18910) );
  AND U27758 ( .A(a[26]), .B(b[73]), .Z(n18909) );
  XOR U27759 ( .A(n18914), .B(n18222), .Z(n18224) );
  IV U27760 ( .A(n18732), .Z(n18222) );
  XOR U27761 ( .A(n18915), .B(n18916), .Z(n18732) );
  ANDN U27762 ( .B(n18917), .A(n18918), .Z(n18915) );
  AND U27763 ( .A(a[27]), .B(b[72]), .Z(n18914) );
  XOR U27764 ( .A(n18919), .B(n18227), .Z(n18229) );
  IV U27765 ( .A(n18730), .Z(n18227) );
  XOR U27766 ( .A(n18920), .B(n18921), .Z(n18730) );
  ANDN U27767 ( .B(n18922), .A(n18923), .Z(n18920) );
  AND U27768 ( .A(a[28]), .B(b[71]), .Z(n18919) );
  XOR U27769 ( .A(n18924), .B(n18232), .Z(n18234) );
  IV U27770 ( .A(n18728), .Z(n18232) );
  XOR U27771 ( .A(n18925), .B(n18926), .Z(n18728) );
  ANDN U27772 ( .B(n18927), .A(n18928), .Z(n18925) );
  AND U27773 ( .A(a[29]), .B(b[70]), .Z(n18924) );
  XOR U27774 ( .A(n18929), .B(n18237), .Z(n18239) );
  IV U27775 ( .A(n18726), .Z(n18237) );
  XOR U27776 ( .A(n18930), .B(n18931), .Z(n18726) );
  ANDN U27777 ( .B(n18932), .A(n18933), .Z(n18930) );
  AND U27778 ( .A(a[30]), .B(b[69]), .Z(n18929) );
  XOR U27779 ( .A(n18934), .B(n18242), .Z(n18244) );
  IV U27780 ( .A(n18724), .Z(n18242) );
  XOR U27781 ( .A(n18935), .B(n18936), .Z(n18724) );
  ANDN U27782 ( .B(n18937), .A(n18938), .Z(n18935) );
  AND U27783 ( .A(a[31]), .B(b[68]), .Z(n18934) );
  XOR U27784 ( .A(n18939), .B(n18247), .Z(n18249) );
  IV U27785 ( .A(n18722), .Z(n18247) );
  XOR U27786 ( .A(n18940), .B(n18941), .Z(n18722) );
  ANDN U27787 ( .B(n18942), .A(n18943), .Z(n18940) );
  AND U27788 ( .A(a[32]), .B(b[67]), .Z(n18939) );
  XOR U27789 ( .A(n18944), .B(n18252), .Z(n18254) );
  IV U27790 ( .A(n18720), .Z(n18252) );
  XOR U27791 ( .A(n18945), .B(n18946), .Z(n18720) );
  ANDN U27792 ( .B(n18947), .A(n18948), .Z(n18945) );
  AND U27793 ( .A(a[33]), .B(b[66]), .Z(n18944) );
  XOR U27794 ( .A(n18949), .B(n18257), .Z(n18259) );
  IV U27795 ( .A(n18718), .Z(n18257) );
  XOR U27796 ( .A(n18950), .B(n18951), .Z(n18718) );
  ANDN U27797 ( .B(n18952), .A(n18953), .Z(n18950) );
  AND U27798 ( .A(a[34]), .B(b[65]), .Z(n18949) );
  XOR U27799 ( .A(n18954), .B(n18262), .Z(n18264) );
  IV U27800 ( .A(n18716), .Z(n18262) );
  XOR U27801 ( .A(n18955), .B(n18956), .Z(n18716) );
  ANDN U27802 ( .B(n18957), .A(n18958), .Z(n18955) );
  AND U27803 ( .A(a[35]), .B(b[64]), .Z(n18954) );
  XOR U27804 ( .A(n18959), .B(n18267), .Z(n18269) );
  IV U27805 ( .A(n18714), .Z(n18267) );
  XOR U27806 ( .A(n18960), .B(n18961), .Z(n18714) );
  ANDN U27807 ( .B(n18962), .A(n18963), .Z(n18960) );
  AND U27808 ( .A(a[36]), .B(b[63]), .Z(n18959) );
  XOR U27809 ( .A(n18964), .B(n18272), .Z(n18274) );
  IV U27810 ( .A(n18712), .Z(n18272) );
  XOR U27811 ( .A(n18965), .B(n18966), .Z(n18712) );
  ANDN U27812 ( .B(n18967), .A(n18968), .Z(n18965) );
  AND U27813 ( .A(a[37]), .B(b[62]), .Z(n18964) );
  XOR U27814 ( .A(n18969), .B(n18277), .Z(n18279) );
  IV U27815 ( .A(n18710), .Z(n18277) );
  XOR U27816 ( .A(n18970), .B(n18971), .Z(n18710) );
  ANDN U27817 ( .B(n18972), .A(n18973), .Z(n18970) );
  AND U27818 ( .A(a[38]), .B(b[61]), .Z(n18969) );
  XOR U27819 ( .A(n18974), .B(n18282), .Z(n18284) );
  IV U27820 ( .A(n18708), .Z(n18282) );
  XOR U27821 ( .A(n18975), .B(n18976), .Z(n18708) );
  ANDN U27822 ( .B(n18977), .A(n18978), .Z(n18975) );
  AND U27823 ( .A(a[39]), .B(b[60]), .Z(n18974) );
  XOR U27824 ( .A(n18979), .B(n18287), .Z(n18289) );
  IV U27825 ( .A(n18706), .Z(n18287) );
  XOR U27826 ( .A(n18980), .B(n18981), .Z(n18706) );
  ANDN U27827 ( .B(n18982), .A(n18983), .Z(n18980) );
  AND U27828 ( .A(a[40]), .B(b[59]), .Z(n18979) );
  XOR U27829 ( .A(n18984), .B(n18292), .Z(n18294) );
  IV U27830 ( .A(n18704), .Z(n18292) );
  XOR U27831 ( .A(n18985), .B(n18986), .Z(n18704) );
  ANDN U27832 ( .B(n18987), .A(n18988), .Z(n18985) );
  AND U27833 ( .A(a[41]), .B(b[58]), .Z(n18984) );
  XOR U27834 ( .A(n18989), .B(n18297), .Z(n18299) );
  IV U27835 ( .A(n18702), .Z(n18297) );
  XOR U27836 ( .A(n18990), .B(n18991), .Z(n18702) );
  ANDN U27837 ( .B(n18992), .A(n18993), .Z(n18990) );
  AND U27838 ( .A(a[42]), .B(b[57]), .Z(n18989) );
  XOR U27839 ( .A(n18994), .B(n18302), .Z(n18304) );
  IV U27840 ( .A(n18700), .Z(n18302) );
  XOR U27841 ( .A(n18995), .B(n18996), .Z(n18700) );
  ANDN U27842 ( .B(n18997), .A(n18998), .Z(n18995) );
  AND U27843 ( .A(a[43]), .B(b[56]), .Z(n18994) );
  XOR U27844 ( .A(n18999), .B(n18307), .Z(n18309) );
  IV U27845 ( .A(n18698), .Z(n18307) );
  XOR U27846 ( .A(n19000), .B(n19001), .Z(n18698) );
  ANDN U27847 ( .B(n19002), .A(n19003), .Z(n19000) );
  AND U27848 ( .A(a[44]), .B(b[55]), .Z(n18999) );
  XOR U27849 ( .A(n19004), .B(n18312), .Z(n18314) );
  IV U27850 ( .A(n18696), .Z(n18312) );
  XOR U27851 ( .A(n19005), .B(n19006), .Z(n18696) );
  ANDN U27852 ( .B(n19007), .A(n19008), .Z(n19005) );
  AND U27853 ( .A(a[45]), .B(b[54]), .Z(n19004) );
  XOR U27854 ( .A(n19009), .B(n18317), .Z(n18319) );
  IV U27855 ( .A(n18694), .Z(n18317) );
  XOR U27856 ( .A(n19010), .B(n19011), .Z(n18694) );
  ANDN U27857 ( .B(n19012), .A(n19013), .Z(n19010) );
  AND U27858 ( .A(a[46]), .B(b[53]), .Z(n19009) );
  XOR U27859 ( .A(n19014), .B(n18322), .Z(n18324) );
  IV U27860 ( .A(n18692), .Z(n18322) );
  XOR U27861 ( .A(n19015), .B(n19016), .Z(n18692) );
  ANDN U27862 ( .B(n19017), .A(n19018), .Z(n19015) );
  AND U27863 ( .A(a[47]), .B(b[52]), .Z(n19014) );
  XOR U27864 ( .A(n19019), .B(n18327), .Z(n18329) );
  IV U27865 ( .A(n18690), .Z(n18327) );
  XOR U27866 ( .A(n19020), .B(n19021), .Z(n18690) );
  ANDN U27867 ( .B(n19022), .A(n19023), .Z(n19020) );
  AND U27868 ( .A(a[48]), .B(b[51]), .Z(n19019) );
  XOR U27869 ( .A(n19024), .B(n18332), .Z(n18334) );
  IV U27870 ( .A(n18688), .Z(n18332) );
  XOR U27871 ( .A(n19025), .B(n19026), .Z(n18688) );
  ANDN U27872 ( .B(n19027), .A(n19028), .Z(n19025) );
  AND U27873 ( .A(a[49]), .B(b[50]), .Z(n19024) );
  XOR U27874 ( .A(n19029), .B(n18337), .Z(n18339) );
  IV U27875 ( .A(n18686), .Z(n18337) );
  XOR U27876 ( .A(n19030), .B(n19031), .Z(n18686) );
  ANDN U27877 ( .B(n19032), .A(n19033), .Z(n19030) );
  AND U27878 ( .A(a[50]), .B(b[49]), .Z(n19029) );
  XOR U27879 ( .A(n19034), .B(n18342), .Z(n18344) );
  IV U27880 ( .A(n18684), .Z(n18342) );
  XOR U27881 ( .A(n19035), .B(n19036), .Z(n18684) );
  ANDN U27882 ( .B(n19037), .A(n19038), .Z(n19035) );
  AND U27883 ( .A(a[51]), .B(b[48]), .Z(n19034) );
  XOR U27884 ( .A(n19039), .B(n18347), .Z(n18349) );
  IV U27885 ( .A(n18682), .Z(n18347) );
  XOR U27886 ( .A(n19040), .B(n19041), .Z(n18682) );
  ANDN U27887 ( .B(n19042), .A(n19043), .Z(n19040) );
  AND U27888 ( .A(a[52]), .B(b[47]), .Z(n19039) );
  XOR U27889 ( .A(n19044), .B(n18352), .Z(n18354) );
  IV U27890 ( .A(n18680), .Z(n18352) );
  XOR U27891 ( .A(n19045), .B(n19046), .Z(n18680) );
  ANDN U27892 ( .B(n19047), .A(n19048), .Z(n19045) );
  AND U27893 ( .A(a[53]), .B(b[46]), .Z(n19044) );
  XOR U27894 ( .A(n19049), .B(n18357), .Z(n18359) );
  IV U27895 ( .A(n18678), .Z(n18357) );
  XOR U27896 ( .A(n19050), .B(n19051), .Z(n18678) );
  ANDN U27897 ( .B(n19052), .A(n19053), .Z(n19050) );
  AND U27898 ( .A(a[54]), .B(b[45]), .Z(n19049) );
  XOR U27899 ( .A(n19054), .B(n18362), .Z(n18364) );
  IV U27900 ( .A(n18676), .Z(n18362) );
  XOR U27901 ( .A(n19055), .B(n19056), .Z(n18676) );
  ANDN U27902 ( .B(n19057), .A(n19058), .Z(n19055) );
  AND U27903 ( .A(a[55]), .B(b[44]), .Z(n19054) );
  XOR U27904 ( .A(n19059), .B(n18367), .Z(n18369) );
  IV U27905 ( .A(n18674), .Z(n18367) );
  XOR U27906 ( .A(n19060), .B(n19061), .Z(n18674) );
  ANDN U27907 ( .B(n19062), .A(n19063), .Z(n19060) );
  AND U27908 ( .A(a[56]), .B(b[43]), .Z(n19059) );
  XOR U27909 ( .A(n19064), .B(n18372), .Z(n18374) );
  IV U27910 ( .A(n18672), .Z(n18372) );
  XOR U27911 ( .A(n19065), .B(n19066), .Z(n18672) );
  ANDN U27912 ( .B(n19067), .A(n19068), .Z(n19065) );
  AND U27913 ( .A(a[57]), .B(b[42]), .Z(n19064) );
  XOR U27914 ( .A(n19069), .B(n18377), .Z(n18379) );
  IV U27915 ( .A(n18670), .Z(n18377) );
  XOR U27916 ( .A(n19070), .B(n19071), .Z(n18670) );
  ANDN U27917 ( .B(n19072), .A(n19073), .Z(n19070) );
  AND U27918 ( .A(a[58]), .B(b[41]), .Z(n19069) );
  XOR U27919 ( .A(n19074), .B(n18382), .Z(n18384) );
  IV U27920 ( .A(n18668), .Z(n18382) );
  XOR U27921 ( .A(n19075), .B(n19076), .Z(n18668) );
  ANDN U27922 ( .B(n19077), .A(n19078), .Z(n19075) );
  AND U27923 ( .A(a[59]), .B(b[40]), .Z(n19074) );
  XOR U27924 ( .A(n19079), .B(n18387), .Z(n18389) );
  IV U27925 ( .A(n18666), .Z(n18387) );
  XOR U27926 ( .A(n19080), .B(n19081), .Z(n18666) );
  ANDN U27927 ( .B(n19082), .A(n19083), .Z(n19080) );
  AND U27928 ( .A(a[60]), .B(b[39]), .Z(n19079) );
  XOR U27929 ( .A(n19084), .B(n18392), .Z(n18394) );
  IV U27930 ( .A(n18664), .Z(n18392) );
  XOR U27931 ( .A(n19085), .B(n19086), .Z(n18664) );
  ANDN U27932 ( .B(n19087), .A(n19088), .Z(n19085) );
  AND U27933 ( .A(a[61]), .B(b[38]), .Z(n19084) );
  XOR U27934 ( .A(n19089), .B(n18397), .Z(n18399) );
  IV U27935 ( .A(n18662), .Z(n18397) );
  XOR U27936 ( .A(n19090), .B(n19091), .Z(n18662) );
  ANDN U27937 ( .B(n19092), .A(n19093), .Z(n19090) );
  AND U27938 ( .A(a[62]), .B(b[37]), .Z(n19089) );
  XOR U27939 ( .A(n19094), .B(n18402), .Z(n18404) );
  IV U27940 ( .A(n18660), .Z(n18402) );
  XOR U27941 ( .A(n19095), .B(n19096), .Z(n18660) );
  ANDN U27942 ( .B(n19097), .A(n19098), .Z(n19095) );
  AND U27943 ( .A(a[63]), .B(b[36]), .Z(n19094) );
  XOR U27944 ( .A(n19099), .B(n18407), .Z(n18409) );
  IV U27945 ( .A(n18658), .Z(n18407) );
  XOR U27946 ( .A(n19100), .B(n19101), .Z(n18658) );
  ANDN U27947 ( .B(n19102), .A(n19103), .Z(n19100) );
  AND U27948 ( .A(a[64]), .B(b[35]), .Z(n19099) );
  XOR U27949 ( .A(n19104), .B(n18412), .Z(n18414) );
  IV U27950 ( .A(n18656), .Z(n18412) );
  XOR U27951 ( .A(n19105), .B(n19106), .Z(n18656) );
  ANDN U27952 ( .B(n19107), .A(n19108), .Z(n19105) );
  AND U27953 ( .A(a[65]), .B(b[34]), .Z(n19104) );
  XOR U27954 ( .A(n19109), .B(n18417), .Z(n18419) );
  IV U27955 ( .A(n18654), .Z(n18417) );
  XOR U27956 ( .A(n19110), .B(n19111), .Z(n18654) );
  ANDN U27957 ( .B(n19112), .A(n19113), .Z(n19110) );
  AND U27958 ( .A(a[66]), .B(b[33]), .Z(n19109) );
  XOR U27959 ( .A(n19114), .B(n18422), .Z(n18424) );
  IV U27960 ( .A(n18652), .Z(n18422) );
  XOR U27961 ( .A(n19115), .B(n19116), .Z(n18652) );
  ANDN U27962 ( .B(n19117), .A(n19118), .Z(n19115) );
  AND U27963 ( .A(a[67]), .B(b[32]), .Z(n19114) );
  XOR U27964 ( .A(n19119), .B(n18427), .Z(n18429) );
  IV U27965 ( .A(n18650), .Z(n18427) );
  XOR U27966 ( .A(n19120), .B(n19121), .Z(n18650) );
  ANDN U27967 ( .B(n19122), .A(n19123), .Z(n19120) );
  AND U27968 ( .A(a[68]), .B(b[31]), .Z(n19119) );
  XOR U27969 ( .A(n19124), .B(n18432), .Z(n18434) );
  IV U27970 ( .A(n18648), .Z(n18432) );
  XOR U27971 ( .A(n19125), .B(n19126), .Z(n18648) );
  ANDN U27972 ( .B(n19127), .A(n19128), .Z(n19125) );
  AND U27973 ( .A(a[69]), .B(b[30]), .Z(n19124) );
  XOR U27974 ( .A(n19129), .B(n18437), .Z(n18439) );
  IV U27975 ( .A(n18646), .Z(n18437) );
  XOR U27976 ( .A(n19130), .B(n19131), .Z(n18646) );
  ANDN U27977 ( .B(n19132), .A(n19133), .Z(n19130) );
  AND U27978 ( .A(a[70]), .B(b[29]), .Z(n19129) );
  XOR U27979 ( .A(n19134), .B(n18442), .Z(n18444) );
  IV U27980 ( .A(n18644), .Z(n18442) );
  XOR U27981 ( .A(n19135), .B(n19136), .Z(n18644) );
  ANDN U27982 ( .B(n19137), .A(n19138), .Z(n19135) );
  AND U27983 ( .A(a[71]), .B(b[28]), .Z(n19134) );
  XOR U27984 ( .A(n19139), .B(n18447), .Z(n18449) );
  IV U27985 ( .A(n18642), .Z(n18447) );
  XOR U27986 ( .A(n19140), .B(n19141), .Z(n18642) );
  ANDN U27987 ( .B(n19142), .A(n19143), .Z(n19140) );
  AND U27988 ( .A(a[72]), .B(b[27]), .Z(n19139) );
  XOR U27989 ( .A(n19144), .B(n18452), .Z(n18454) );
  IV U27990 ( .A(n18640), .Z(n18452) );
  XOR U27991 ( .A(n19145), .B(n19146), .Z(n18640) );
  ANDN U27992 ( .B(n19147), .A(n19148), .Z(n19145) );
  AND U27993 ( .A(a[73]), .B(b[26]), .Z(n19144) );
  XOR U27994 ( .A(n19149), .B(n18457), .Z(n18459) );
  IV U27995 ( .A(n18638), .Z(n18457) );
  XOR U27996 ( .A(n19150), .B(n19151), .Z(n18638) );
  ANDN U27997 ( .B(n19152), .A(n19153), .Z(n19150) );
  AND U27998 ( .A(a[74]), .B(b[25]), .Z(n19149) );
  XOR U27999 ( .A(n19154), .B(n18462), .Z(n18464) );
  IV U28000 ( .A(n18636), .Z(n18462) );
  XOR U28001 ( .A(n19155), .B(n19156), .Z(n18636) );
  ANDN U28002 ( .B(n19157), .A(n19158), .Z(n19155) );
  AND U28003 ( .A(a[75]), .B(b[24]), .Z(n19154) );
  XOR U28004 ( .A(n19159), .B(n18467), .Z(n18469) );
  IV U28005 ( .A(n18634), .Z(n18467) );
  XOR U28006 ( .A(n19160), .B(n19161), .Z(n18634) );
  ANDN U28007 ( .B(n19162), .A(n19163), .Z(n19160) );
  AND U28008 ( .A(a[76]), .B(b[23]), .Z(n19159) );
  XOR U28009 ( .A(n19164), .B(n18472), .Z(n18474) );
  IV U28010 ( .A(n18632), .Z(n18472) );
  XOR U28011 ( .A(n19165), .B(n19166), .Z(n18632) );
  ANDN U28012 ( .B(n19167), .A(n19168), .Z(n19165) );
  AND U28013 ( .A(a[77]), .B(b[22]), .Z(n19164) );
  XOR U28014 ( .A(n19169), .B(n18477), .Z(n18479) );
  IV U28015 ( .A(n18630), .Z(n18477) );
  XOR U28016 ( .A(n19170), .B(n19171), .Z(n18630) );
  ANDN U28017 ( .B(n19172), .A(n19173), .Z(n19170) );
  AND U28018 ( .A(a[78]), .B(b[21]), .Z(n19169) );
  XOR U28019 ( .A(n19174), .B(n18482), .Z(n18484) );
  IV U28020 ( .A(n18628), .Z(n18482) );
  XOR U28021 ( .A(n19175), .B(n19176), .Z(n18628) );
  ANDN U28022 ( .B(n19177), .A(n19178), .Z(n19175) );
  AND U28023 ( .A(a[79]), .B(b[20]), .Z(n19174) );
  XOR U28024 ( .A(n19179), .B(n18487), .Z(n18489) );
  IV U28025 ( .A(n18626), .Z(n18487) );
  XOR U28026 ( .A(n19180), .B(n19181), .Z(n18626) );
  ANDN U28027 ( .B(n19182), .A(n19183), .Z(n19180) );
  AND U28028 ( .A(a[80]), .B(b[19]), .Z(n19179) );
  XOR U28029 ( .A(n19184), .B(n18492), .Z(n18494) );
  IV U28030 ( .A(n18624), .Z(n18492) );
  XOR U28031 ( .A(n19185), .B(n19186), .Z(n18624) );
  ANDN U28032 ( .B(n19187), .A(n19188), .Z(n19185) );
  AND U28033 ( .A(a[81]), .B(b[18]), .Z(n19184) );
  XOR U28034 ( .A(n19189), .B(n18497), .Z(n18499) );
  IV U28035 ( .A(n18622), .Z(n18497) );
  XOR U28036 ( .A(n19190), .B(n19191), .Z(n18622) );
  ANDN U28037 ( .B(n19192), .A(n19193), .Z(n19190) );
  AND U28038 ( .A(a[82]), .B(b[17]), .Z(n19189) );
  XOR U28039 ( .A(n19194), .B(n18502), .Z(n18504) );
  IV U28040 ( .A(n18620), .Z(n18502) );
  XOR U28041 ( .A(n19195), .B(n19196), .Z(n18620) );
  ANDN U28042 ( .B(n19197), .A(n19198), .Z(n19195) );
  AND U28043 ( .A(a[83]), .B(b[16]), .Z(n19194) );
  XOR U28044 ( .A(n19199), .B(n18507), .Z(n18509) );
  IV U28045 ( .A(n18618), .Z(n18507) );
  XOR U28046 ( .A(n19200), .B(n19201), .Z(n18618) );
  ANDN U28047 ( .B(n19202), .A(n19203), .Z(n19200) );
  AND U28048 ( .A(a[84]), .B(b[15]), .Z(n19199) );
  XOR U28049 ( .A(n19204), .B(n18512), .Z(n18514) );
  IV U28050 ( .A(n18616), .Z(n18512) );
  XOR U28051 ( .A(n19205), .B(n19206), .Z(n18616) );
  ANDN U28052 ( .B(n19207), .A(n19208), .Z(n19205) );
  AND U28053 ( .A(a[85]), .B(b[14]), .Z(n19204) );
  XOR U28054 ( .A(n19209), .B(n18517), .Z(n18519) );
  IV U28055 ( .A(n18614), .Z(n18517) );
  XOR U28056 ( .A(n19210), .B(n19211), .Z(n18614) );
  ANDN U28057 ( .B(n19212), .A(n19213), .Z(n19210) );
  AND U28058 ( .A(a[86]), .B(b[13]), .Z(n19209) );
  XOR U28059 ( .A(n19214), .B(n18522), .Z(n18524) );
  IV U28060 ( .A(n18612), .Z(n18522) );
  XOR U28061 ( .A(n19215), .B(n19216), .Z(n18612) );
  ANDN U28062 ( .B(n19217), .A(n19218), .Z(n19215) );
  AND U28063 ( .A(a[87]), .B(b[12]), .Z(n19214) );
  XOR U28064 ( .A(n19219), .B(n18527), .Z(n18529) );
  IV U28065 ( .A(n18610), .Z(n18527) );
  XOR U28066 ( .A(n19220), .B(n19221), .Z(n18610) );
  ANDN U28067 ( .B(n19222), .A(n19223), .Z(n19220) );
  AND U28068 ( .A(a[88]), .B(b[11]), .Z(n19219) );
  XOR U28069 ( .A(n19224), .B(n18532), .Z(n18534) );
  IV U28070 ( .A(n18608), .Z(n18532) );
  XOR U28071 ( .A(n19225), .B(n19226), .Z(n18608) );
  ANDN U28072 ( .B(n19227), .A(n19228), .Z(n19225) );
  AND U28073 ( .A(a[89]), .B(b[10]), .Z(n19224) );
  XOR U28074 ( .A(n19229), .B(n18537), .Z(n18539) );
  IV U28075 ( .A(n18606), .Z(n18537) );
  XOR U28076 ( .A(n19230), .B(n19231), .Z(n18606) );
  ANDN U28077 ( .B(n19232), .A(n19233), .Z(n19230) );
  AND U28078 ( .A(b[9]), .B(a[90]), .Z(n19229) );
  XOR U28079 ( .A(n19234), .B(n18542), .Z(n18544) );
  IV U28080 ( .A(n18604), .Z(n18542) );
  XOR U28081 ( .A(n19235), .B(n19236), .Z(n18604) );
  ANDN U28082 ( .B(n19237), .A(n19238), .Z(n19235) );
  AND U28083 ( .A(b[8]), .B(a[91]), .Z(n19234) );
  XOR U28084 ( .A(n19239), .B(n18547), .Z(n18549) );
  IV U28085 ( .A(n18602), .Z(n18547) );
  XOR U28086 ( .A(n19240), .B(n19241), .Z(n18602) );
  ANDN U28087 ( .B(n19242), .A(n19243), .Z(n19240) );
  AND U28088 ( .A(b[7]), .B(a[92]), .Z(n19239) );
  XOR U28089 ( .A(n19244), .B(n18552), .Z(n18554) );
  IV U28090 ( .A(n18600), .Z(n18552) );
  XOR U28091 ( .A(n19245), .B(n19246), .Z(n18600) );
  ANDN U28092 ( .B(n19247), .A(n19248), .Z(n19245) );
  AND U28093 ( .A(b[6]), .B(a[93]), .Z(n19244) );
  XOR U28094 ( .A(n19249), .B(n18557), .Z(n18559) );
  IV U28095 ( .A(n18598), .Z(n18557) );
  XOR U28096 ( .A(n19250), .B(n19251), .Z(n18598) );
  ANDN U28097 ( .B(n19252), .A(n19253), .Z(n19250) );
  AND U28098 ( .A(b[5]), .B(a[94]), .Z(n19249) );
  XOR U28099 ( .A(n19254), .B(n18562), .Z(n18564) );
  IV U28100 ( .A(n18596), .Z(n18562) );
  XOR U28101 ( .A(n19255), .B(n19256), .Z(n18596) );
  ANDN U28102 ( .B(n19257), .A(n19258), .Z(n19255) );
  AND U28103 ( .A(b[4]), .B(a[95]), .Z(n19254) );
  XOR U28104 ( .A(n19259), .B(n18567), .Z(n18569) );
  IV U28105 ( .A(n18594), .Z(n18567) );
  XOR U28106 ( .A(n19260), .B(n19261), .Z(n18594) );
  ANDN U28107 ( .B(n18588), .A(n18589), .Z(n19260) );
  AND U28108 ( .A(b[2]), .B(a[96]), .Z(n19262) );
  XNOR U28109 ( .A(n19257), .B(n19261), .Z(n19263) );
  XOR U28110 ( .A(n19264), .B(n19265), .Z(n19261) );
  OR U28111 ( .A(n18591), .B(n18592), .Z(n19265) );
  XNOR U28112 ( .A(n19267), .B(n19268), .Z(n19266) );
  XOR U28113 ( .A(n19267), .B(n19270), .Z(n18591) );
  NAND U28114 ( .A(b[1]), .B(a[96]), .Z(n19270) );
  IV U28115 ( .A(n19264), .Z(n19267) );
  NANDN U28116 ( .A(n9), .B(n10), .Z(n19264) );
  XOR U28117 ( .A(n19271), .B(n19272), .Z(n10) );
  NAND U28118 ( .A(a[96]), .B(b[0]), .Z(n9) );
  XNOR U28119 ( .A(n19252), .B(n19256), .Z(n19273) );
  XNOR U28120 ( .A(n19247), .B(n19251), .Z(n19274) );
  XNOR U28121 ( .A(n19242), .B(n19246), .Z(n19275) );
  XNOR U28122 ( .A(n19237), .B(n19241), .Z(n19276) );
  XNOR U28123 ( .A(n19232), .B(n19236), .Z(n19277) );
  XNOR U28124 ( .A(n19227), .B(n19231), .Z(n19278) );
  XNOR U28125 ( .A(n19222), .B(n19226), .Z(n19279) );
  XNOR U28126 ( .A(n19217), .B(n19221), .Z(n19280) );
  XNOR U28127 ( .A(n19212), .B(n19216), .Z(n19281) );
  XNOR U28128 ( .A(n19207), .B(n19211), .Z(n19282) );
  XNOR U28129 ( .A(n19202), .B(n19206), .Z(n19283) );
  XNOR U28130 ( .A(n19197), .B(n19201), .Z(n19284) );
  XNOR U28131 ( .A(n19192), .B(n19196), .Z(n19285) );
  XNOR U28132 ( .A(n19187), .B(n19191), .Z(n19286) );
  XNOR U28133 ( .A(n19182), .B(n19186), .Z(n19287) );
  XNOR U28134 ( .A(n19177), .B(n19181), .Z(n19288) );
  XNOR U28135 ( .A(n19172), .B(n19176), .Z(n19289) );
  XNOR U28136 ( .A(n19167), .B(n19171), .Z(n19290) );
  XNOR U28137 ( .A(n19162), .B(n19166), .Z(n19291) );
  XNOR U28138 ( .A(n19157), .B(n19161), .Z(n19292) );
  XNOR U28139 ( .A(n19152), .B(n19156), .Z(n19293) );
  XNOR U28140 ( .A(n19147), .B(n19151), .Z(n19294) );
  XNOR U28141 ( .A(n19142), .B(n19146), .Z(n19295) );
  XNOR U28142 ( .A(n19137), .B(n19141), .Z(n19296) );
  XNOR U28143 ( .A(n19132), .B(n19136), .Z(n19297) );
  XNOR U28144 ( .A(n19127), .B(n19131), .Z(n19298) );
  XNOR U28145 ( .A(n19122), .B(n19126), .Z(n19299) );
  XNOR U28146 ( .A(n19117), .B(n19121), .Z(n19300) );
  XNOR U28147 ( .A(n19112), .B(n19116), .Z(n19301) );
  XNOR U28148 ( .A(n19107), .B(n19111), .Z(n19302) );
  XNOR U28149 ( .A(n19102), .B(n19106), .Z(n19303) );
  XNOR U28150 ( .A(n19097), .B(n19101), .Z(n19304) );
  XNOR U28151 ( .A(n19092), .B(n19096), .Z(n19305) );
  XNOR U28152 ( .A(n19087), .B(n19091), .Z(n19306) );
  XNOR U28153 ( .A(n19082), .B(n19086), .Z(n19307) );
  XNOR U28154 ( .A(n19077), .B(n19081), .Z(n19308) );
  XNOR U28155 ( .A(n19072), .B(n19076), .Z(n19309) );
  XNOR U28156 ( .A(n19067), .B(n19071), .Z(n19310) );
  XNOR U28157 ( .A(n19062), .B(n19066), .Z(n19311) );
  XNOR U28158 ( .A(n19057), .B(n19061), .Z(n19312) );
  XNOR U28159 ( .A(n19052), .B(n19056), .Z(n19313) );
  XNOR U28160 ( .A(n19047), .B(n19051), .Z(n19314) );
  XNOR U28161 ( .A(n19042), .B(n19046), .Z(n19315) );
  XNOR U28162 ( .A(n19037), .B(n19041), .Z(n19316) );
  XNOR U28163 ( .A(n19032), .B(n19036), .Z(n19317) );
  XNOR U28164 ( .A(n19027), .B(n19031), .Z(n19318) );
  XNOR U28165 ( .A(n19022), .B(n19026), .Z(n19319) );
  XNOR U28166 ( .A(n19017), .B(n19021), .Z(n19320) );
  XNOR U28167 ( .A(n19012), .B(n19016), .Z(n19321) );
  XNOR U28168 ( .A(n19007), .B(n19011), .Z(n19322) );
  XNOR U28169 ( .A(n19002), .B(n19006), .Z(n19323) );
  XNOR U28170 ( .A(n18997), .B(n19001), .Z(n19324) );
  XNOR U28171 ( .A(n18992), .B(n18996), .Z(n19325) );
  XNOR U28172 ( .A(n18987), .B(n18991), .Z(n19326) );
  XNOR U28173 ( .A(n18982), .B(n18986), .Z(n19327) );
  XNOR U28174 ( .A(n18977), .B(n18981), .Z(n19328) );
  XNOR U28175 ( .A(n18972), .B(n18976), .Z(n19329) );
  XNOR U28176 ( .A(n18967), .B(n18971), .Z(n19330) );
  XNOR U28177 ( .A(n18962), .B(n18966), .Z(n19331) );
  XNOR U28178 ( .A(n18957), .B(n18961), .Z(n19332) );
  XNOR U28179 ( .A(n18952), .B(n18956), .Z(n19333) );
  XNOR U28180 ( .A(n18947), .B(n18951), .Z(n19334) );
  XNOR U28181 ( .A(n18942), .B(n18946), .Z(n19335) );
  XNOR U28182 ( .A(n18937), .B(n18941), .Z(n19336) );
  XNOR U28183 ( .A(n18932), .B(n18936), .Z(n19337) );
  XNOR U28184 ( .A(n18927), .B(n18931), .Z(n19338) );
  XNOR U28185 ( .A(n18922), .B(n18926), .Z(n19339) );
  XNOR U28186 ( .A(n18917), .B(n18921), .Z(n19340) );
  XNOR U28187 ( .A(n18912), .B(n18916), .Z(n19341) );
  XNOR U28188 ( .A(n18907), .B(n18911), .Z(n19342) );
  XNOR U28189 ( .A(n18902), .B(n18906), .Z(n19343) );
  XNOR U28190 ( .A(n18897), .B(n18901), .Z(n19344) );
  XNOR U28191 ( .A(n18892), .B(n18896), .Z(n19345) );
  XNOR U28192 ( .A(n18887), .B(n18891), .Z(n19346) );
  XNOR U28193 ( .A(n18882), .B(n18886), .Z(n19347) );
  XNOR U28194 ( .A(n18877), .B(n18881), .Z(n19348) );
  XNOR U28195 ( .A(n18872), .B(n18876), .Z(n19349) );
  XNOR U28196 ( .A(n18867), .B(n18871), .Z(n19350) );
  XNOR U28197 ( .A(n18862), .B(n18866), .Z(n19351) );
  XNOR U28198 ( .A(n18857), .B(n18861), .Z(n19352) );
  XNOR U28199 ( .A(n18852), .B(n18856), .Z(n19353) );
  XNOR U28200 ( .A(n18847), .B(n18851), .Z(n19354) );
  XNOR U28201 ( .A(n18842), .B(n18846), .Z(n19355) );
  XNOR U28202 ( .A(n18837), .B(n18841), .Z(n19356) );
  XNOR U28203 ( .A(n18832), .B(n18836), .Z(n19357) );
  XNOR U28204 ( .A(n18827), .B(n18831), .Z(n19358) );
  XNOR U28205 ( .A(n18822), .B(n18826), .Z(n19359) );
  XNOR U28206 ( .A(n18817), .B(n18821), .Z(n19360) );
  XNOR U28207 ( .A(n18812), .B(n18816), .Z(n19361) );
  XNOR U28208 ( .A(n18807), .B(n18811), .Z(n19362) );
  XNOR U28209 ( .A(n18802), .B(n18806), .Z(n19363) );
  XNOR U28210 ( .A(n18797), .B(n18801), .Z(n19364) );
  XNOR U28211 ( .A(n18792), .B(n18796), .Z(n19365) );
  XNOR U28212 ( .A(n18787), .B(n18791), .Z(n19366) );
  XOR U28213 ( .A(n19367), .B(n18786), .Z(n18787) );
  AND U28214 ( .A(a[0]), .B(b[98]), .Z(n19367) );
  XNOR U28215 ( .A(n19368), .B(n18786), .Z(n18788) );
  XNOR U28216 ( .A(n19369), .B(n19370), .Z(n18786) );
  ANDN U28217 ( .B(n19371), .A(n19372), .Z(n19369) );
  AND U28218 ( .A(a[1]), .B(b[97]), .Z(n19368) );
  XOR U28219 ( .A(n19374), .B(n19375), .Z(n18791) );
  ANDN U28220 ( .B(n19376), .A(n19377), .Z(n19374) );
  AND U28221 ( .A(a[2]), .B(b[96]), .Z(n19373) );
  XOR U28222 ( .A(n19379), .B(n19380), .Z(n18796) );
  ANDN U28223 ( .B(n19381), .A(n19382), .Z(n19379) );
  AND U28224 ( .A(a[3]), .B(b[95]), .Z(n19378) );
  XOR U28225 ( .A(n19384), .B(n19385), .Z(n18801) );
  ANDN U28226 ( .B(n19386), .A(n19387), .Z(n19384) );
  AND U28227 ( .A(a[4]), .B(b[94]), .Z(n19383) );
  XOR U28228 ( .A(n19389), .B(n19390), .Z(n18806) );
  ANDN U28229 ( .B(n19391), .A(n19392), .Z(n19389) );
  AND U28230 ( .A(a[5]), .B(b[93]), .Z(n19388) );
  XOR U28231 ( .A(n19394), .B(n19395), .Z(n18811) );
  ANDN U28232 ( .B(n19396), .A(n19397), .Z(n19394) );
  AND U28233 ( .A(a[6]), .B(b[92]), .Z(n19393) );
  XOR U28234 ( .A(n19399), .B(n19400), .Z(n18816) );
  ANDN U28235 ( .B(n19401), .A(n19402), .Z(n19399) );
  AND U28236 ( .A(a[7]), .B(b[91]), .Z(n19398) );
  XOR U28237 ( .A(n19404), .B(n19405), .Z(n18821) );
  ANDN U28238 ( .B(n19406), .A(n19407), .Z(n19404) );
  AND U28239 ( .A(a[8]), .B(b[90]), .Z(n19403) );
  XOR U28240 ( .A(n19409), .B(n19410), .Z(n18826) );
  ANDN U28241 ( .B(n19411), .A(n19412), .Z(n19409) );
  AND U28242 ( .A(a[9]), .B(b[89]), .Z(n19408) );
  XOR U28243 ( .A(n19414), .B(n19415), .Z(n18831) );
  ANDN U28244 ( .B(n19416), .A(n19417), .Z(n19414) );
  AND U28245 ( .A(a[10]), .B(b[88]), .Z(n19413) );
  XOR U28246 ( .A(n19419), .B(n19420), .Z(n18836) );
  ANDN U28247 ( .B(n19421), .A(n19422), .Z(n19419) );
  AND U28248 ( .A(a[11]), .B(b[87]), .Z(n19418) );
  XOR U28249 ( .A(n19424), .B(n19425), .Z(n18841) );
  ANDN U28250 ( .B(n19426), .A(n19427), .Z(n19424) );
  AND U28251 ( .A(a[12]), .B(b[86]), .Z(n19423) );
  XOR U28252 ( .A(n19429), .B(n19430), .Z(n18846) );
  ANDN U28253 ( .B(n19431), .A(n19432), .Z(n19429) );
  AND U28254 ( .A(a[13]), .B(b[85]), .Z(n19428) );
  XOR U28255 ( .A(n19434), .B(n19435), .Z(n18851) );
  ANDN U28256 ( .B(n19436), .A(n19437), .Z(n19434) );
  AND U28257 ( .A(a[14]), .B(b[84]), .Z(n19433) );
  XOR U28258 ( .A(n19439), .B(n19440), .Z(n18856) );
  ANDN U28259 ( .B(n19441), .A(n19442), .Z(n19439) );
  AND U28260 ( .A(a[15]), .B(b[83]), .Z(n19438) );
  XOR U28261 ( .A(n19444), .B(n19445), .Z(n18861) );
  ANDN U28262 ( .B(n19446), .A(n19447), .Z(n19444) );
  AND U28263 ( .A(a[16]), .B(b[82]), .Z(n19443) );
  XOR U28264 ( .A(n19449), .B(n19450), .Z(n18866) );
  ANDN U28265 ( .B(n19451), .A(n19452), .Z(n19449) );
  AND U28266 ( .A(a[17]), .B(b[81]), .Z(n19448) );
  XOR U28267 ( .A(n19454), .B(n19455), .Z(n18871) );
  ANDN U28268 ( .B(n19456), .A(n19457), .Z(n19454) );
  AND U28269 ( .A(a[18]), .B(b[80]), .Z(n19453) );
  XOR U28270 ( .A(n19459), .B(n19460), .Z(n18876) );
  ANDN U28271 ( .B(n19461), .A(n19462), .Z(n19459) );
  AND U28272 ( .A(a[19]), .B(b[79]), .Z(n19458) );
  XOR U28273 ( .A(n19464), .B(n19465), .Z(n18881) );
  ANDN U28274 ( .B(n19466), .A(n19467), .Z(n19464) );
  AND U28275 ( .A(a[20]), .B(b[78]), .Z(n19463) );
  XOR U28276 ( .A(n19469), .B(n19470), .Z(n18886) );
  ANDN U28277 ( .B(n19471), .A(n19472), .Z(n19469) );
  AND U28278 ( .A(a[21]), .B(b[77]), .Z(n19468) );
  XOR U28279 ( .A(n19474), .B(n19475), .Z(n18891) );
  ANDN U28280 ( .B(n19476), .A(n19477), .Z(n19474) );
  AND U28281 ( .A(a[22]), .B(b[76]), .Z(n19473) );
  XOR U28282 ( .A(n19479), .B(n19480), .Z(n18896) );
  ANDN U28283 ( .B(n19481), .A(n19482), .Z(n19479) );
  AND U28284 ( .A(a[23]), .B(b[75]), .Z(n19478) );
  XOR U28285 ( .A(n19484), .B(n19485), .Z(n18901) );
  ANDN U28286 ( .B(n19486), .A(n19487), .Z(n19484) );
  AND U28287 ( .A(a[24]), .B(b[74]), .Z(n19483) );
  XOR U28288 ( .A(n19489), .B(n19490), .Z(n18906) );
  ANDN U28289 ( .B(n19491), .A(n19492), .Z(n19489) );
  AND U28290 ( .A(a[25]), .B(b[73]), .Z(n19488) );
  XOR U28291 ( .A(n19494), .B(n19495), .Z(n18911) );
  ANDN U28292 ( .B(n19496), .A(n19497), .Z(n19494) );
  AND U28293 ( .A(a[26]), .B(b[72]), .Z(n19493) );
  XOR U28294 ( .A(n19499), .B(n19500), .Z(n18916) );
  ANDN U28295 ( .B(n19501), .A(n19502), .Z(n19499) );
  AND U28296 ( .A(a[27]), .B(b[71]), .Z(n19498) );
  XOR U28297 ( .A(n19504), .B(n19505), .Z(n18921) );
  ANDN U28298 ( .B(n19506), .A(n19507), .Z(n19504) );
  AND U28299 ( .A(a[28]), .B(b[70]), .Z(n19503) );
  XOR U28300 ( .A(n19509), .B(n19510), .Z(n18926) );
  ANDN U28301 ( .B(n19511), .A(n19512), .Z(n19509) );
  AND U28302 ( .A(a[29]), .B(b[69]), .Z(n19508) );
  XOR U28303 ( .A(n19514), .B(n19515), .Z(n18931) );
  ANDN U28304 ( .B(n19516), .A(n19517), .Z(n19514) );
  AND U28305 ( .A(a[30]), .B(b[68]), .Z(n19513) );
  XOR U28306 ( .A(n19519), .B(n19520), .Z(n18936) );
  ANDN U28307 ( .B(n19521), .A(n19522), .Z(n19519) );
  AND U28308 ( .A(a[31]), .B(b[67]), .Z(n19518) );
  XOR U28309 ( .A(n19524), .B(n19525), .Z(n18941) );
  ANDN U28310 ( .B(n19526), .A(n19527), .Z(n19524) );
  AND U28311 ( .A(a[32]), .B(b[66]), .Z(n19523) );
  XOR U28312 ( .A(n19529), .B(n19530), .Z(n18946) );
  ANDN U28313 ( .B(n19531), .A(n19532), .Z(n19529) );
  AND U28314 ( .A(a[33]), .B(b[65]), .Z(n19528) );
  XOR U28315 ( .A(n19534), .B(n19535), .Z(n18951) );
  ANDN U28316 ( .B(n19536), .A(n19537), .Z(n19534) );
  AND U28317 ( .A(a[34]), .B(b[64]), .Z(n19533) );
  XOR U28318 ( .A(n19539), .B(n19540), .Z(n18956) );
  ANDN U28319 ( .B(n19541), .A(n19542), .Z(n19539) );
  AND U28320 ( .A(a[35]), .B(b[63]), .Z(n19538) );
  XOR U28321 ( .A(n19544), .B(n19545), .Z(n18961) );
  ANDN U28322 ( .B(n19546), .A(n19547), .Z(n19544) );
  AND U28323 ( .A(a[36]), .B(b[62]), .Z(n19543) );
  XOR U28324 ( .A(n19549), .B(n19550), .Z(n18966) );
  ANDN U28325 ( .B(n19551), .A(n19552), .Z(n19549) );
  AND U28326 ( .A(a[37]), .B(b[61]), .Z(n19548) );
  XOR U28327 ( .A(n19554), .B(n19555), .Z(n18971) );
  ANDN U28328 ( .B(n19556), .A(n19557), .Z(n19554) );
  AND U28329 ( .A(a[38]), .B(b[60]), .Z(n19553) );
  XOR U28330 ( .A(n19559), .B(n19560), .Z(n18976) );
  ANDN U28331 ( .B(n19561), .A(n19562), .Z(n19559) );
  AND U28332 ( .A(a[39]), .B(b[59]), .Z(n19558) );
  XOR U28333 ( .A(n19564), .B(n19565), .Z(n18981) );
  ANDN U28334 ( .B(n19566), .A(n19567), .Z(n19564) );
  AND U28335 ( .A(a[40]), .B(b[58]), .Z(n19563) );
  XOR U28336 ( .A(n19569), .B(n19570), .Z(n18986) );
  ANDN U28337 ( .B(n19571), .A(n19572), .Z(n19569) );
  AND U28338 ( .A(a[41]), .B(b[57]), .Z(n19568) );
  XOR U28339 ( .A(n19574), .B(n19575), .Z(n18991) );
  ANDN U28340 ( .B(n19576), .A(n19577), .Z(n19574) );
  AND U28341 ( .A(a[42]), .B(b[56]), .Z(n19573) );
  XOR U28342 ( .A(n19579), .B(n19580), .Z(n18996) );
  ANDN U28343 ( .B(n19581), .A(n19582), .Z(n19579) );
  AND U28344 ( .A(a[43]), .B(b[55]), .Z(n19578) );
  XOR U28345 ( .A(n19584), .B(n19585), .Z(n19001) );
  ANDN U28346 ( .B(n19586), .A(n19587), .Z(n19584) );
  AND U28347 ( .A(a[44]), .B(b[54]), .Z(n19583) );
  XOR U28348 ( .A(n19589), .B(n19590), .Z(n19006) );
  ANDN U28349 ( .B(n19591), .A(n19592), .Z(n19589) );
  AND U28350 ( .A(a[45]), .B(b[53]), .Z(n19588) );
  XOR U28351 ( .A(n19594), .B(n19595), .Z(n19011) );
  ANDN U28352 ( .B(n19596), .A(n19597), .Z(n19594) );
  AND U28353 ( .A(a[46]), .B(b[52]), .Z(n19593) );
  XOR U28354 ( .A(n19599), .B(n19600), .Z(n19016) );
  ANDN U28355 ( .B(n19601), .A(n19602), .Z(n19599) );
  AND U28356 ( .A(a[47]), .B(b[51]), .Z(n19598) );
  XOR U28357 ( .A(n19604), .B(n19605), .Z(n19021) );
  ANDN U28358 ( .B(n19606), .A(n19607), .Z(n19604) );
  AND U28359 ( .A(a[48]), .B(b[50]), .Z(n19603) );
  XOR U28360 ( .A(n19609), .B(n19610), .Z(n19026) );
  ANDN U28361 ( .B(n19611), .A(n19612), .Z(n19609) );
  AND U28362 ( .A(a[49]), .B(b[49]), .Z(n19608) );
  XOR U28363 ( .A(n19614), .B(n19615), .Z(n19031) );
  ANDN U28364 ( .B(n19616), .A(n19617), .Z(n19614) );
  AND U28365 ( .A(a[50]), .B(b[48]), .Z(n19613) );
  XOR U28366 ( .A(n19619), .B(n19620), .Z(n19036) );
  ANDN U28367 ( .B(n19621), .A(n19622), .Z(n19619) );
  AND U28368 ( .A(a[51]), .B(b[47]), .Z(n19618) );
  XOR U28369 ( .A(n19624), .B(n19625), .Z(n19041) );
  ANDN U28370 ( .B(n19626), .A(n19627), .Z(n19624) );
  AND U28371 ( .A(a[52]), .B(b[46]), .Z(n19623) );
  XOR U28372 ( .A(n19629), .B(n19630), .Z(n19046) );
  ANDN U28373 ( .B(n19631), .A(n19632), .Z(n19629) );
  AND U28374 ( .A(a[53]), .B(b[45]), .Z(n19628) );
  XOR U28375 ( .A(n19634), .B(n19635), .Z(n19051) );
  ANDN U28376 ( .B(n19636), .A(n19637), .Z(n19634) );
  AND U28377 ( .A(a[54]), .B(b[44]), .Z(n19633) );
  XOR U28378 ( .A(n19639), .B(n19640), .Z(n19056) );
  ANDN U28379 ( .B(n19641), .A(n19642), .Z(n19639) );
  AND U28380 ( .A(a[55]), .B(b[43]), .Z(n19638) );
  XOR U28381 ( .A(n19644), .B(n19645), .Z(n19061) );
  ANDN U28382 ( .B(n19646), .A(n19647), .Z(n19644) );
  AND U28383 ( .A(a[56]), .B(b[42]), .Z(n19643) );
  XOR U28384 ( .A(n19649), .B(n19650), .Z(n19066) );
  ANDN U28385 ( .B(n19651), .A(n19652), .Z(n19649) );
  AND U28386 ( .A(a[57]), .B(b[41]), .Z(n19648) );
  XOR U28387 ( .A(n19654), .B(n19655), .Z(n19071) );
  ANDN U28388 ( .B(n19656), .A(n19657), .Z(n19654) );
  AND U28389 ( .A(a[58]), .B(b[40]), .Z(n19653) );
  XOR U28390 ( .A(n19659), .B(n19660), .Z(n19076) );
  ANDN U28391 ( .B(n19661), .A(n19662), .Z(n19659) );
  AND U28392 ( .A(a[59]), .B(b[39]), .Z(n19658) );
  XOR U28393 ( .A(n19664), .B(n19665), .Z(n19081) );
  ANDN U28394 ( .B(n19666), .A(n19667), .Z(n19664) );
  AND U28395 ( .A(a[60]), .B(b[38]), .Z(n19663) );
  XOR U28396 ( .A(n19669), .B(n19670), .Z(n19086) );
  ANDN U28397 ( .B(n19671), .A(n19672), .Z(n19669) );
  AND U28398 ( .A(a[61]), .B(b[37]), .Z(n19668) );
  XOR U28399 ( .A(n19674), .B(n19675), .Z(n19091) );
  ANDN U28400 ( .B(n19676), .A(n19677), .Z(n19674) );
  AND U28401 ( .A(a[62]), .B(b[36]), .Z(n19673) );
  XOR U28402 ( .A(n19679), .B(n19680), .Z(n19096) );
  ANDN U28403 ( .B(n19681), .A(n19682), .Z(n19679) );
  AND U28404 ( .A(a[63]), .B(b[35]), .Z(n19678) );
  XOR U28405 ( .A(n19684), .B(n19685), .Z(n19101) );
  ANDN U28406 ( .B(n19686), .A(n19687), .Z(n19684) );
  AND U28407 ( .A(a[64]), .B(b[34]), .Z(n19683) );
  XOR U28408 ( .A(n19689), .B(n19690), .Z(n19106) );
  ANDN U28409 ( .B(n19691), .A(n19692), .Z(n19689) );
  AND U28410 ( .A(a[65]), .B(b[33]), .Z(n19688) );
  XOR U28411 ( .A(n19694), .B(n19695), .Z(n19111) );
  ANDN U28412 ( .B(n19696), .A(n19697), .Z(n19694) );
  AND U28413 ( .A(a[66]), .B(b[32]), .Z(n19693) );
  XOR U28414 ( .A(n19699), .B(n19700), .Z(n19116) );
  ANDN U28415 ( .B(n19701), .A(n19702), .Z(n19699) );
  AND U28416 ( .A(a[67]), .B(b[31]), .Z(n19698) );
  XOR U28417 ( .A(n19704), .B(n19705), .Z(n19121) );
  ANDN U28418 ( .B(n19706), .A(n19707), .Z(n19704) );
  AND U28419 ( .A(a[68]), .B(b[30]), .Z(n19703) );
  XOR U28420 ( .A(n19709), .B(n19710), .Z(n19126) );
  ANDN U28421 ( .B(n19711), .A(n19712), .Z(n19709) );
  AND U28422 ( .A(a[69]), .B(b[29]), .Z(n19708) );
  XOR U28423 ( .A(n19714), .B(n19715), .Z(n19131) );
  ANDN U28424 ( .B(n19716), .A(n19717), .Z(n19714) );
  AND U28425 ( .A(a[70]), .B(b[28]), .Z(n19713) );
  XOR U28426 ( .A(n19719), .B(n19720), .Z(n19136) );
  ANDN U28427 ( .B(n19721), .A(n19722), .Z(n19719) );
  AND U28428 ( .A(a[71]), .B(b[27]), .Z(n19718) );
  XOR U28429 ( .A(n19724), .B(n19725), .Z(n19141) );
  ANDN U28430 ( .B(n19726), .A(n19727), .Z(n19724) );
  AND U28431 ( .A(a[72]), .B(b[26]), .Z(n19723) );
  XOR U28432 ( .A(n19729), .B(n19730), .Z(n19146) );
  ANDN U28433 ( .B(n19731), .A(n19732), .Z(n19729) );
  AND U28434 ( .A(a[73]), .B(b[25]), .Z(n19728) );
  XOR U28435 ( .A(n19734), .B(n19735), .Z(n19151) );
  ANDN U28436 ( .B(n19736), .A(n19737), .Z(n19734) );
  AND U28437 ( .A(a[74]), .B(b[24]), .Z(n19733) );
  XOR U28438 ( .A(n19739), .B(n19740), .Z(n19156) );
  ANDN U28439 ( .B(n19741), .A(n19742), .Z(n19739) );
  AND U28440 ( .A(a[75]), .B(b[23]), .Z(n19738) );
  XOR U28441 ( .A(n19744), .B(n19745), .Z(n19161) );
  ANDN U28442 ( .B(n19746), .A(n19747), .Z(n19744) );
  AND U28443 ( .A(a[76]), .B(b[22]), .Z(n19743) );
  XOR U28444 ( .A(n19749), .B(n19750), .Z(n19166) );
  ANDN U28445 ( .B(n19751), .A(n19752), .Z(n19749) );
  AND U28446 ( .A(a[77]), .B(b[21]), .Z(n19748) );
  XOR U28447 ( .A(n19754), .B(n19755), .Z(n19171) );
  ANDN U28448 ( .B(n19756), .A(n19757), .Z(n19754) );
  AND U28449 ( .A(a[78]), .B(b[20]), .Z(n19753) );
  XOR U28450 ( .A(n19759), .B(n19760), .Z(n19176) );
  ANDN U28451 ( .B(n19761), .A(n19762), .Z(n19759) );
  AND U28452 ( .A(a[79]), .B(b[19]), .Z(n19758) );
  XOR U28453 ( .A(n19764), .B(n19765), .Z(n19181) );
  ANDN U28454 ( .B(n19766), .A(n19767), .Z(n19764) );
  AND U28455 ( .A(a[80]), .B(b[18]), .Z(n19763) );
  XOR U28456 ( .A(n19769), .B(n19770), .Z(n19186) );
  ANDN U28457 ( .B(n19771), .A(n19772), .Z(n19769) );
  AND U28458 ( .A(a[81]), .B(b[17]), .Z(n19768) );
  XOR U28459 ( .A(n19774), .B(n19775), .Z(n19191) );
  ANDN U28460 ( .B(n19776), .A(n19777), .Z(n19774) );
  AND U28461 ( .A(a[82]), .B(b[16]), .Z(n19773) );
  XOR U28462 ( .A(n19779), .B(n19780), .Z(n19196) );
  ANDN U28463 ( .B(n19781), .A(n19782), .Z(n19779) );
  AND U28464 ( .A(a[83]), .B(b[15]), .Z(n19778) );
  XOR U28465 ( .A(n19784), .B(n19785), .Z(n19201) );
  ANDN U28466 ( .B(n19786), .A(n19787), .Z(n19784) );
  AND U28467 ( .A(a[84]), .B(b[14]), .Z(n19783) );
  XOR U28468 ( .A(n19789), .B(n19790), .Z(n19206) );
  ANDN U28469 ( .B(n19791), .A(n19792), .Z(n19789) );
  AND U28470 ( .A(a[85]), .B(b[13]), .Z(n19788) );
  XOR U28471 ( .A(n19794), .B(n19795), .Z(n19211) );
  ANDN U28472 ( .B(n19796), .A(n19797), .Z(n19794) );
  AND U28473 ( .A(a[86]), .B(b[12]), .Z(n19793) );
  XOR U28474 ( .A(n19799), .B(n19800), .Z(n19216) );
  ANDN U28475 ( .B(n19801), .A(n19802), .Z(n19799) );
  AND U28476 ( .A(a[87]), .B(b[11]), .Z(n19798) );
  XOR U28477 ( .A(n19804), .B(n19805), .Z(n19221) );
  ANDN U28478 ( .B(n19806), .A(n19807), .Z(n19804) );
  AND U28479 ( .A(a[88]), .B(b[10]), .Z(n19803) );
  XOR U28480 ( .A(n19809), .B(n19810), .Z(n19226) );
  ANDN U28481 ( .B(n19811), .A(n19812), .Z(n19809) );
  AND U28482 ( .A(b[9]), .B(a[89]), .Z(n19808) );
  XOR U28483 ( .A(n19814), .B(n19815), .Z(n19231) );
  ANDN U28484 ( .B(n19816), .A(n19817), .Z(n19814) );
  AND U28485 ( .A(b[8]), .B(a[90]), .Z(n19813) );
  XOR U28486 ( .A(n19819), .B(n19820), .Z(n19236) );
  ANDN U28487 ( .B(n19821), .A(n19822), .Z(n19819) );
  AND U28488 ( .A(b[7]), .B(a[91]), .Z(n19818) );
  XOR U28489 ( .A(n19824), .B(n19825), .Z(n19241) );
  ANDN U28490 ( .B(n19826), .A(n19827), .Z(n19824) );
  AND U28491 ( .A(b[6]), .B(a[92]), .Z(n19823) );
  XOR U28492 ( .A(n19829), .B(n19830), .Z(n19246) );
  ANDN U28493 ( .B(n19831), .A(n19832), .Z(n19829) );
  AND U28494 ( .A(b[5]), .B(a[93]), .Z(n19828) );
  XOR U28495 ( .A(n19834), .B(n19835), .Z(n19251) );
  ANDN U28496 ( .B(n19836), .A(n19837), .Z(n19834) );
  AND U28497 ( .A(b[4]), .B(a[94]), .Z(n19833) );
  XOR U28498 ( .A(n19839), .B(n19840), .Z(n19256) );
  ANDN U28499 ( .B(n19268), .A(n19269), .Z(n19839) );
  AND U28500 ( .A(b[2]), .B(a[95]), .Z(n19841) );
  XNOR U28501 ( .A(n19836), .B(n19840), .Z(n19842) );
  XOR U28502 ( .A(n19843), .B(n19844), .Z(n19840) );
  OR U28503 ( .A(n19271), .B(n19272), .Z(n19844) );
  XNOR U28504 ( .A(n19846), .B(n19847), .Z(n19845) );
  XOR U28505 ( .A(n19846), .B(n19849), .Z(n19271) );
  NAND U28506 ( .A(b[1]), .B(a[95]), .Z(n19849) );
  IV U28507 ( .A(n19843), .Z(n19846) );
  NANDN U28508 ( .A(n11), .B(n12), .Z(n19843) );
  XOR U28509 ( .A(n19850), .B(n19851), .Z(n12) );
  NAND U28510 ( .A(a[95]), .B(b[0]), .Z(n11) );
  XNOR U28511 ( .A(n19831), .B(n19835), .Z(n19852) );
  XNOR U28512 ( .A(n19826), .B(n19830), .Z(n19853) );
  XNOR U28513 ( .A(n19821), .B(n19825), .Z(n19854) );
  XNOR U28514 ( .A(n19816), .B(n19820), .Z(n19855) );
  XNOR U28515 ( .A(n19811), .B(n19815), .Z(n19856) );
  XNOR U28516 ( .A(n19806), .B(n19810), .Z(n19857) );
  XNOR U28517 ( .A(n19801), .B(n19805), .Z(n19858) );
  XNOR U28518 ( .A(n19796), .B(n19800), .Z(n19859) );
  XNOR U28519 ( .A(n19791), .B(n19795), .Z(n19860) );
  XNOR U28520 ( .A(n19786), .B(n19790), .Z(n19861) );
  XNOR U28521 ( .A(n19781), .B(n19785), .Z(n19862) );
  XNOR U28522 ( .A(n19776), .B(n19780), .Z(n19863) );
  XNOR U28523 ( .A(n19771), .B(n19775), .Z(n19864) );
  XNOR U28524 ( .A(n19766), .B(n19770), .Z(n19865) );
  XNOR U28525 ( .A(n19761), .B(n19765), .Z(n19866) );
  XNOR U28526 ( .A(n19756), .B(n19760), .Z(n19867) );
  XNOR U28527 ( .A(n19751), .B(n19755), .Z(n19868) );
  XNOR U28528 ( .A(n19746), .B(n19750), .Z(n19869) );
  XNOR U28529 ( .A(n19741), .B(n19745), .Z(n19870) );
  XNOR U28530 ( .A(n19736), .B(n19740), .Z(n19871) );
  XNOR U28531 ( .A(n19731), .B(n19735), .Z(n19872) );
  XNOR U28532 ( .A(n19726), .B(n19730), .Z(n19873) );
  XNOR U28533 ( .A(n19721), .B(n19725), .Z(n19874) );
  XNOR U28534 ( .A(n19716), .B(n19720), .Z(n19875) );
  XNOR U28535 ( .A(n19711), .B(n19715), .Z(n19876) );
  XNOR U28536 ( .A(n19706), .B(n19710), .Z(n19877) );
  XNOR U28537 ( .A(n19701), .B(n19705), .Z(n19878) );
  XNOR U28538 ( .A(n19696), .B(n19700), .Z(n19879) );
  XNOR U28539 ( .A(n19691), .B(n19695), .Z(n19880) );
  XNOR U28540 ( .A(n19686), .B(n19690), .Z(n19881) );
  XNOR U28541 ( .A(n19681), .B(n19685), .Z(n19882) );
  XNOR U28542 ( .A(n19676), .B(n19680), .Z(n19883) );
  XNOR U28543 ( .A(n19671), .B(n19675), .Z(n19884) );
  XNOR U28544 ( .A(n19666), .B(n19670), .Z(n19885) );
  XNOR U28545 ( .A(n19661), .B(n19665), .Z(n19886) );
  XNOR U28546 ( .A(n19656), .B(n19660), .Z(n19887) );
  XNOR U28547 ( .A(n19651), .B(n19655), .Z(n19888) );
  XNOR U28548 ( .A(n19646), .B(n19650), .Z(n19889) );
  XNOR U28549 ( .A(n19641), .B(n19645), .Z(n19890) );
  XNOR U28550 ( .A(n19636), .B(n19640), .Z(n19891) );
  XNOR U28551 ( .A(n19631), .B(n19635), .Z(n19892) );
  XNOR U28552 ( .A(n19626), .B(n19630), .Z(n19893) );
  XNOR U28553 ( .A(n19621), .B(n19625), .Z(n19894) );
  XNOR U28554 ( .A(n19616), .B(n19620), .Z(n19895) );
  XNOR U28555 ( .A(n19611), .B(n19615), .Z(n19896) );
  XNOR U28556 ( .A(n19606), .B(n19610), .Z(n19897) );
  XNOR U28557 ( .A(n19601), .B(n19605), .Z(n19898) );
  XNOR U28558 ( .A(n19596), .B(n19600), .Z(n19899) );
  XNOR U28559 ( .A(n19591), .B(n19595), .Z(n19900) );
  XNOR U28560 ( .A(n19586), .B(n19590), .Z(n19901) );
  XNOR U28561 ( .A(n19581), .B(n19585), .Z(n19902) );
  XNOR U28562 ( .A(n19576), .B(n19580), .Z(n19903) );
  XNOR U28563 ( .A(n19571), .B(n19575), .Z(n19904) );
  XNOR U28564 ( .A(n19566), .B(n19570), .Z(n19905) );
  XNOR U28565 ( .A(n19561), .B(n19565), .Z(n19906) );
  XNOR U28566 ( .A(n19556), .B(n19560), .Z(n19907) );
  XNOR U28567 ( .A(n19551), .B(n19555), .Z(n19908) );
  XNOR U28568 ( .A(n19546), .B(n19550), .Z(n19909) );
  XNOR U28569 ( .A(n19541), .B(n19545), .Z(n19910) );
  XNOR U28570 ( .A(n19536), .B(n19540), .Z(n19911) );
  XNOR U28571 ( .A(n19531), .B(n19535), .Z(n19912) );
  XNOR U28572 ( .A(n19526), .B(n19530), .Z(n19913) );
  XNOR U28573 ( .A(n19521), .B(n19525), .Z(n19914) );
  XNOR U28574 ( .A(n19516), .B(n19520), .Z(n19915) );
  XNOR U28575 ( .A(n19511), .B(n19515), .Z(n19916) );
  XNOR U28576 ( .A(n19506), .B(n19510), .Z(n19917) );
  XNOR U28577 ( .A(n19501), .B(n19505), .Z(n19918) );
  XNOR U28578 ( .A(n19496), .B(n19500), .Z(n19919) );
  XNOR U28579 ( .A(n19491), .B(n19495), .Z(n19920) );
  XNOR U28580 ( .A(n19486), .B(n19490), .Z(n19921) );
  XNOR U28581 ( .A(n19481), .B(n19485), .Z(n19922) );
  XNOR U28582 ( .A(n19476), .B(n19480), .Z(n19923) );
  XNOR U28583 ( .A(n19471), .B(n19475), .Z(n19924) );
  XNOR U28584 ( .A(n19466), .B(n19470), .Z(n19925) );
  XNOR U28585 ( .A(n19461), .B(n19465), .Z(n19926) );
  XNOR U28586 ( .A(n19456), .B(n19460), .Z(n19927) );
  XNOR U28587 ( .A(n19451), .B(n19455), .Z(n19928) );
  XNOR U28588 ( .A(n19446), .B(n19450), .Z(n19929) );
  XNOR U28589 ( .A(n19441), .B(n19445), .Z(n19930) );
  XNOR U28590 ( .A(n19436), .B(n19440), .Z(n19931) );
  XNOR U28591 ( .A(n19431), .B(n19435), .Z(n19932) );
  XNOR U28592 ( .A(n19426), .B(n19430), .Z(n19933) );
  XNOR U28593 ( .A(n19421), .B(n19425), .Z(n19934) );
  XNOR U28594 ( .A(n19416), .B(n19420), .Z(n19935) );
  XNOR U28595 ( .A(n19411), .B(n19415), .Z(n19936) );
  XNOR U28596 ( .A(n19406), .B(n19410), .Z(n19937) );
  XNOR U28597 ( .A(n19401), .B(n19405), .Z(n19938) );
  XNOR U28598 ( .A(n19396), .B(n19400), .Z(n19939) );
  XNOR U28599 ( .A(n19391), .B(n19395), .Z(n19940) );
  XNOR U28600 ( .A(n19386), .B(n19390), .Z(n19941) );
  XNOR U28601 ( .A(n19381), .B(n19385), .Z(n19942) );
  XNOR U28602 ( .A(n19376), .B(n19380), .Z(n19943) );
  XNOR U28603 ( .A(n19371), .B(n19375), .Z(n19944) );
  XNOR U28604 ( .A(n19945), .B(n19370), .Z(n19371) );
  AND U28605 ( .A(a[0]), .B(b[97]), .Z(n19945) );
  XOR U28606 ( .A(n19946), .B(n19370), .Z(n19372) );
  XNOR U28607 ( .A(n19947), .B(n19948), .Z(n19370) );
  ANDN U28608 ( .B(n19949), .A(n19950), .Z(n19947) );
  AND U28609 ( .A(a[1]), .B(b[96]), .Z(n19946) );
  XOR U28610 ( .A(n19952), .B(n19953), .Z(n19375) );
  ANDN U28611 ( .B(n19954), .A(n19955), .Z(n19952) );
  AND U28612 ( .A(a[2]), .B(b[95]), .Z(n19951) );
  XOR U28613 ( .A(n19957), .B(n19958), .Z(n19380) );
  ANDN U28614 ( .B(n19959), .A(n19960), .Z(n19957) );
  AND U28615 ( .A(a[3]), .B(b[94]), .Z(n19956) );
  XOR U28616 ( .A(n19962), .B(n19963), .Z(n19385) );
  ANDN U28617 ( .B(n19964), .A(n19965), .Z(n19962) );
  AND U28618 ( .A(a[4]), .B(b[93]), .Z(n19961) );
  XOR U28619 ( .A(n19967), .B(n19968), .Z(n19390) );
  ANDN U28620 ( .B(n19969), .A(n19970), .Z(n19967) );
  AND U28621 ( .A(a[5]), .B(b[92]), .Z(n19966) );
  XOR U28622 ( .A(n19972), .B(n19973), .Z(n19395) );
  ANDN U28623 ( .B(n19974), .A(n19975), .Z(n19972) );
  AND U28624 ( .A(a[6]), .B(b[91]), .Z(n19971) );
  XOR U28625 ( .A(n19977), .B(n19978), .Z(n19400) );
  ANDN U28626 ( .B(n19979), .A(n19980), .Z(n19977) );
  AND U28627 ( .A(a[7]), .B(b[90]), .Z(n19976) );
  XOR U28628 ( .A(n19982), .B(n19983), .Z(n19405) );
  ANDN U28629 ( .B(n19984), .A(n19985), .Z(n19982) );
  AND U28630 ( .A(a[8]), .B(b[89]), .Z(n19981) );
  XOR U28631 ( .A(n19987), .B(n19988), .Z(n19410) );
  ANDN U28632 ( .B(n19989), .A(n19990), .Z(n19987) );
  AND U28633 ( .A(a[9]), .B(b[88]), .Z(n19986) );
  XOR U28634 ( .A(n19992), .B(n19993), .Z(n19415) );
  ANDN U28635 ( .B(n19994), .A(n19995), .Z(n19992) );
  AND U28636 ( .A(a[10]), .B(b[87]), .Z(n19991) );
  XOR U28637 ( .A(n19997), .B(n19998), .Z(n19420) );
  ANDN U28638 ( .B(n19999), .A(n20000), .Z(n19997) );
  AND U28639 ( .A(a[11]), .B(b[86]), .Z(n19996) );
  XOR U28640 ( .A(n20002), .B(n20003), .Z(n19425) );
  ANDN U28641 ( .B(n20004), .A(n20005), .Z(n20002) );
  AND U28642 ( .A(a[12]), .B(b[85]), .Z(n20001) );
  XOR U28643 ( .A(n20007), .B(n20008), .Z(n19430) );
  ANDN U28644 ( .B(n20009), .A(n20010), .Z(n20007) );
  AND U28645 ( .A(a[13]), .B(b[84]), .Z(n20006) );
  XOR U28646 ( .A(n20012), .B(n20013), .Z(n19435) );
  ANDN U28647 ( .B(n20014), .A(n20015), .Z(n20012) );
  AND U28648 ( .A(a[14]), .B(b[83]), .Z(n20011) );
  XOR U28649 ( .A(n20017), .B(n20018), .Z(n19440) );
  ANDN U28650 ( .B(n20019), .A(n20020), .Z(n20017) );
  AND U28651 ( .A(a[15]), .B(b[82]), .Z(n20016) );
  XOR U28652 ( .A(n20022), .B(n20023), .Z(n19445) );
  ANDN U28653 ( .B(n20024), .A(n20025), .Z(n20022) );
  AND U28654 ( .A(a[16]), .B(b[81]), .Z(n20021) );
  XOR U28655 ( .A(n20027), .B(n20028), .Z(n19450) );
  ANDN U28656 ( .B(n20029), .A(n20030), .Z(n20027) );
  AND U28657 ( .A(a[17]), .B(b[80]), .Z(n20026) );
  XOR U28658 ( .A(n20032), .B(n20033), .Z(n19455) );
  ANDN U28659 ( .B(n20034), .A(n20035), .Z(n20032) );
  AND U28660 ( .A(a[18]), .B(b[79]), .Z(n20031) );
  XOR U28661 ( .A(n20037), .B(n20038), .Z(n19460) );
  ANDN U28662 ( .B(n20039), .A(n20040), .Z(n20037) );
  AND U28663 ( .A(a[19]), .B(b[78]), .Z(n20036) );
  XOR U28664 ( .A(n20042), .B(n20043), .Z(n19465) );
  ANDN U28665 ( .B(n20044), .A(n20045), .Z(n20042) );
  AND U28666 ( .A(a[20]), .B(b[77]), .Z(n20041) );
  XOR U28667 ( .A(n20047), .B(n20048), .Z(n19470) );
  ANDN U28668 ( .B(n20049), .A(n20050), .Z(n20047) );
  AND U28669 ( .A(a[21]), .B(b[76]), .Z(n20046) );
  XOR U28670 ( .A(n20052), .B(n20053), .Z(n19475) );
  ANDN U28671 ( .B(n20054), .A(n20055), .Z(n20052) );
  AND U28672 ( .A(a[22]), .B(b[75]), .Z(n20051) );
  XOR U28673 ( .A(n20057), .B(n20058), .Z(n19480) );
  ANDN U28674 ( .B(n20059), .A(n20060), .Z(n20057) );
  AND U28675 ( .A(a[23]), .B(b[74]), .Z(n20056) );
  XOR U28676 ( .A(n20062), .B(n20063), .Z(n19485) );
  ANDN U28677 ( .B(n20064), .A(n20065), .Z(n20062) );
  AND U28678 ( .A(a[24]), .B(b[73]), .Z(n20061) );
  XOR U28679 ( .A(n20067), .B(n20068), .Z(n19490) );
  ANDN U28680 ( .B(n20069), .A(n20070), .Z(n20067) );
  AND U28681 ( .A(a[25]), .B(b[72]), .Z(n20066) );
  XOR U28682 ( .A(n20072), .B(n20073), .Z(n19495) );
  ANDN U28683 ( .B(n20074), .A(n20075), .Z(n20072) );
  AND U28684 ( .A(a[26]), .B(b[71]), .Z(n20071) );
  XOR U28685 ( .A(n20077), .B(n20078), .Z(n19500) );
  ANDN U28686 ( .B(n20079), .A(n20080), .Z(n20077) );
  AND U28687 ( .A(a[27]), .B(b[70]), .Z(n20076) );
  XOR U28688 ( .A(n20082), .B(n20083), .Z(n19505) );
  ANDN U28689 ( .B(n20084), .A(n20085), .Z(n20082) );
  AND U28690 ( .A(a[28]), .B(b[69]), .Z(n20081) );
  XOR U28691 ( .A(n20087), .B(n20088), .Z(n19510) );
  ANDN U28692 ( .B(n20089), .A(n20090), .Z(n20087) );
  AND U28693 ( .A(a[29]), .B(b[68]), .Z(n20086) );
  XOR U28694 ( .A(n20092), .B(n20093), .Z(n19515) );
  ANDN U28695 ( .B(n20094), .A(n20095), .Z(n20092) );
  AND U28696 ( .A(a[30]), .B(b[67]), .Z(n20091) );
  XOR U28697 ( .A(n20097), .B(n20098), .Z(n19520) );
  ANDN U28698 ( .B(n20099), .A(n20100), .Z(n20097) );
  AND U28699 ( .A(a[31]), .B(b[66]), .Z(n20096) );
  XOR U28700 ( .A(n20102), .B(n20103), .Z(n19525) );
  ANDN U28701 ( .B(n20104), .A(n20105), .Z(n20102) );
  AND U28702 ( .A(a[32]), .B(b[65]), .Z(n20101) );
  XOR U28703 ( .A(n20107), .B(n20108), .Z(n19530) );
  ANDN U28704 ( .B(n20109), .A(n20110), .Z(n20107) );
  AND U28705 ( .A(a[33]), .B(b[64]), .Z(n20106) );
  XOR U28706 ( .A(n20112), .B(n20113), .Z(n19535) );
  ANDN U28707 ( .B(n20114), .A(n20115), .Z(n20112) );
  AND U28708 ( .A(a[34]), .B(b[63]), .Z(n20111) );
  XOR U28709 ( .A(n20117), .B(n20118), .Z(n19540) );
  ANDN U28710 ( .B(n20119), .A(n20120), .Z(n20117) );
  AND U28711 ( .A(a[35]), .B(b[62]), .Z(n20116) );
  XOR U28712 ( .A(n20122), .B(n20123), .Z(n19545) );
  ANDN U28713 ( .B(n20124), .A(n20125), .Z(n20122) );
  AND U28714 ( .A(a[36]), .B(b[61]), .Z(n20121) );
  XOR U28715 ( .A(n20127), .B(n20128), .Z(n19550) );
  ANDN U28716 ( .B(n20129), .A(n20130), .Z(n20127) );
  AND U28717 ( .A(a[37]), .B(b[60]), .Z(n20126) );
  XOR U28718 ( .A(n20132), .B(n20133), .Z(n19555) );
  ANDN U28719 ( .B(n20134), .A(n20135), .Z(n20132) );
  AND U28720 ( .A(a[38]), .B(b[59]), .Z(n20131) );
  XOR U28721 ( .A(n20137), .B(n20138), .Z(n19560) );
  ANDN U28722 ( .B(n20139), .A(n20140), .Z(n20137) );
  AND U28723 ( .A(a[39]), .B(b[58]), .Z(n20136) );
  XOR U28724 ( .A(n20142), .B(n20143), .Z(n19565) );
  ANDN U28725 ( .B(n20144), .A(n20145), .Z(n20142) );
  AND U28726 ( .A(a[40]), .B(b[57]), .Z(n20141) );
  XOR U28727 ( .A(n20147), .B(n20148), .Z(n19570) );
  ANDN U28728 ( .B(n20149), .A(n20150), .Z(n20147) );
  AND U28729 ( .A(a[41]), .B(b[56]), .Z(n20146) );
  XOR U28730 ( .A(n20152), .B(n20153), .Z(n19575) );
  ANDN U28731 ( .B(n20154), .A(n20155), .Z(n20152) );
  AND U28732 ( .A(a[42]), .B(b[55]), .Z(n20151) );
  XOR U28733 ( .A(n20157), .B(n20158), .Z(n19580) );
  ANDN U28734 ( .B(n20159), .A(n20160), .Z(n20157) );
  AND U28735 ( .A(a[43]), .B(b[54]), .Z(n20156) );
  XOR U28736 ( .A(n20162), .B(n20163), .Z(n19585) );
  ANDN U28737 ( .B(n20164), .A(n20165), .Z(n20162) );
  AND U28738 ( .A(a[44]), .B(b[53]), .Z(n20161) );
  XOR U28739 ( .A(n20167), .B(n20168), .Z(n19590) );
  ANDN U28740 ( .B(n20169), .A(n20170), .Z(n20167) );
  AND U28741 ( .A(a[45]), .B(b[52]), .Z(n20166) );
  XOR U28742 ( .A(n20172), .B(n20173), .Z(n19595) );
  ANDN U28743 ( .B(n20174), .A(n20175), .Z(n20172) );
  AND U28744 ( .A(a[46]), .B(b[51]), .Z(n20171) );
  XOR U28745 ( .A(n20177), .B(n20178), .Z(n19600) );
  ANDN U28746 ( .B(n20179), .A(n20180), .Z(n20177) );
  AND U28747 ( .A(a[47]), .B(b[50]), .Z(n20176) );
  XOR U28748 ( .A(n20182), .B(n20183), .Z(n19605) );
  ANDN U28749 ( .B(n20184), .A(n20185), .Z(n20182) );
  AND U28750 ( .A(a[48]), .B(b[49]), .Z(n20181) );
  XOR U28751 ( .A(n20187), .B(n20188), .Z(n19610) );
  ANDN U28752 ( .B(n20189), .A(n20190), .Z(n20187) );
  AND U28753 ( .A(a[49]), .B(b[48]), .Z(n20186) );
  XOR U28754 ( .A(n20192), .B(n20193), .Z(n19615) );
  ANDN U28755 ( .B(n20194), .A(n20195), .Z(n20192) );
  AND U28756 ( .A(a[50]), .B(b[47]), .Z(n20191) );
  XOR U28757 ( .A(n20197), .B(n20198), .Z(n19620) );
  ANDN U28758 ( .B(n20199), .A(n20200), .Z(n20197) );
  AND U28759 ( .A(a[51]), .B(b[46]), .Z(n20196) );
  XOR U28760 ( .A(n20202), .B(n20203), .Z(n19625) );
  ANDN U28761 ( .B(n20204), .A(n20205), .Z(n20202) );
  AND U28762 ( .A(a[52]), .B(b[45]), .Z(n20201) );
  XOR U28763 ( .A(n20207), .B(n20208), .Z(n19630) );
  ANDN U28764 ( .B(n20209), .A(n20210), .Z(n20207) );
  AND U28765 ( .A(a[53]), .B(b[44]), .Z(n20206) );
  XOR U28766 ( .A(n20212), .B(n20213), .Z(n19635) );
  ANDN U28767 ( .B(n20214), .A(n20215), .Z(n20212) );
  AND U28768 ( .A(a[54]), .B(b[43]), .Z(n20211) );
  XOR U28769 ( .A(n20217), .B(n20218), .Z(n19640) );
  ANDN U28770 ( .B(n20219), .A(n20220), .Z(n20217) );
  AND U28771 ( .A(a[55]), .B(b[42]), .Z(n20216) );
  XOR U28772 ( .A(n20222), .B(n20223), .Z(n19645) );
  ANDN U28773 ( .B(n20224), .A(n20225), .Z(n20222) );
  AND U28774 ( .A(a[56]), .B(b[41]), .Z(n20221) );
  XOR U28775 ( .A(n20227), .B(n20228), .Z(n19650) );
  ANDN U28776 ( .B(n20229), .A(n20230), .Z(n20227) );
  AND U28777 ( .A(a[57]), .B(b[40]), .Z(n20226) );
  XOR U28778 ( .A(n20232), .B(n20233), .Z(n19655) );
  ANDN U28779 ( .B(n20234), .A(n20235), .Z(n20232) );
  AND U28780 ( .A(a[58]), .B(b[39]), .Z(n20231) );
  XOR U28781 ( .A(n20237), .B(n20238), .Z(n19660) );
  ANDN U28782 ( .B(n20239), .A(n20240), .Z(n20237) );
  AND U28783 ( .A(a[59]), .B(b[38]), .Z(n20236) );
  XOR U28784 ( .A(n20242), .B(n20243), .Z(n19665) );
  ANDN U28785 ( .B(n20244), .A(n20245), .Z(n20242) );
  AND U28786 ( .A(a[60]), .B(b[37]), .Z(n20241) );
  XOR U28787 ( .A(n20247), .B(n20248), .Z(n19670) );
  ANDN U28788 ( .B(n20249), .A(n20250), .Z(n20247) );
  AND U28789 ( .A(a[61]), .B(b[36]), .Z(n20246) );
  XOR U28790 ( .A(n20252), .B(n20253), .Z(n19675) );
  ANDN U28791 ( .B(n20254), .A(n20255), .Z(n20252) );
  AND U28792 ( .A(a[62]), .B(b[35]), .Z(n20251) );
  XOR U28793 ( .A(n20257), .B(n20258), .Z(n19680) );
  ANDN U28794 ( .B(n20259), .A(n20260), .Z(n20257) );
  AND U28795 ( .A(a[63]), .B(b[34]), .Z(n20256) );
  XOR U28796 ( .A(n20262), .B(n20263), .Z(n19685) );
  ANDN U28797 ( .B(n20264), .A(n20265), .Z(n20262) );
  AND U28798 ( .A(a[64]), .B(b[33]), .Z(n20261) );
  XOR U28799 ( .A(n20267), .B(n20268), .Z(n19690) );
  ANDN U28800 ( .B(n20269), .A(n20270), .Z(n20267) );
  AND U28801 ( .A(a[65]), .B(b[32]), .Z(n20266) );
  XOR U28802 ( .A(n20272), .B(n20273), .Z(n19695) );
  ANDN U28803 ( .B(n20274), .A(n20275), .Z(n20272) );
  AND U28804 ( .A(a[66]), .B(b[31]), .Z(n20271) );
  XOR U28805 ( .A(n20277), .B(n20278), .Z(n19700) );
  ANDN U28806 ( .B(n20279), .A(n20280), .Z(n20277) );
  AND U28807 ( .A(a[67]), .B(b[30]), .Z(n20276) );
  XOR U28808 ( .A(n20282), .B(n20283), .Z(n19705) );
  ANDN U28809 ( .B(n20284), .A(n20285), .Z(n20282) );
  AND U28810 ( .A(a[68]), .B(b[29]), .Z(n20281) );
  XOR U28811 ( .A(n20287), .B(n20288), .Z(n19710) );
  ANDN U28812 ( .B(n20289), .A(n20290), .Z(n20287) );
  AND U28813 ( .A(a[69]), .B(b[28]), .Z(n20286) );
  XOR U28814 ( .A(n20292), .B(n20293), .Z(n19715) );
  ANDN U28815 ( .B(n20294), .A(n20295), .Z(n20292) );
  AND U28816 ( .A(a[70]), .B(b[27]), .Z(n20291) );
  XOR U28817 ( .A(n20297), .B(n20298), .Z(n19720) );
  ANDN U28818 ( .B(n20299), .A(n20300), .Z(n20297) );
  AND U28819 ( .A(a[71]), .B(b[26]), .Z(n20296) );
  XOR U28820 ( .A(n20302), .B(n20303), .Z(n19725) );
  ANDN U28821 ( .B(n20304), .A(n20305), .Z(n20302) );
  AND U28822 ( .A(a[72]), .B(b[25]), .Z(n20301) );
  XOR U28823 ( .A(n20307), .B(n20308), .Z(n19730) );
  ANDN U28824 ( .B(n20309), .A(n20310), .Z(n20307) );
  AND U28825 ( .A(a[73]), .B(b[24]), .Z(n20306) );
  XOR U28826 ( .A(n20312), .B(n20313), .Z(n19735) );
  ANDN U28827 ( .B(n20314), .A(n20315), .Z(n20312) );
  AND U28828 ( .A(a[74]), .B(b[23]), .Z(n20311) );
  XOR U28829 ( .A(n20317), .B(n20318), .Z(n19740) );
  ANDN U28830 ( .B(n20319), .A(n20320), .Z(n20317) );
  AND U28831 ( .A(a[75]), .B(b[22]), .Z(n20316) );
  XOR U28832 ( .A(n20322), .B(n20323), .Z(n19745) );
  ANDN U28833 ( .B(n20324), .A(n20325), .Z(n20322) );
  AND U28834 ( .A(a[76]), .B(b[21]), .Z(n20321) );
  XOR U28835 ( .A(n20327), .B(n20328), .Z(n19750) );
  ANDN U28836 ( .B(n20329), .A(n20330), .Z(n20327) );
  AND U28837 ( .A(a[77]), .B(b[20]), .Z(n20326) );
  XOR U28838 ( .A(n20332), .B(n20333), .Z(n19755) );
  ANDN U28839 ( .B(n20334), .A(n20335), .Z(n20332) );
  AND U28840 ( .A(a[78]), .B(b[19]), .Z(n20331) );
  XOR U28841 ( .A(n20337), .B(n20338), .Z(n19760) );
  ANDN U28842 ( .B(n20339), .A(n20340), .Z(n20337) );
  AND U28843 ( .A(a[79]), .B(b[18]), .Z(n20336) );
  XOR U28844 ( .A(n20342), .B(n20343), .Z(n19765) );
  ANDN U28845 ( .B(n20344), .A(n20345), .Z(n20342) );
  AND U28846 ( .A(a[80]), .B(b[17]), .Z(n20341) );
  XOR U28847 ( .A(n20347), .B(n20348), .Z(n19770) );
  ANDN U28848 ( .B(n20349), .A(n20350), .Z(n20347) );
  AND U28849 ( .A(a[81]), .B(b[16]), .Z(n20346) );
  XOR U28850 ( .A(n20352), .B(n20353), .Z(n19775) );
  ANDN U28851 ( .B(n20354), .A(n20355), .Z(n20352) );
  AND U28852 ( .A(a[82]), .B(b[15]), .Z(n20351) );
  XOR U28853 ( .A(n20357), .B(n20358), .Z(n19780) );
  ANDN U28854 ( .B(n20359), .A(n20360), .Z(n20357) );
  AND U28855 ( .A(a[83]), .B(b[14]), .Z(n20356) );
  XOR U28856 ( .A(n20362), .B(n20363), .Z(n19785) );
  ANDN U28857 ( .B(n20364), .A(n20365), .Z(n20362) );
  AND U28858 ( .A(a[84]), .B(b[13]), .Z(n20361) );
  XOR U28859 ( .A(n20367), .B(n20368), .Z(n19790) );
  ANDN U28860 ( .B(n20369), .A(n20370), .Z(n20367) );
  AND U28861 ( .A(a[85]), .B(b[12]), .Z(n20366) );
  XOR U28862 ( .A(n20372), .B(n20373), .Z(n19795) );
  ANDN U28863 ( .B(n20374), .A(n20375), .Z(n20372) );
  AND U28864 ( .A(a[86]), .B(b[11]), .Z(n20371) );
  XOR U28865 ( .A(n20377), .B(n20378), .Z(n19800) );
  ANDN U28866 ( .B(n20379), .A(n20380), .Z(n20377) );
  AND U28867 ( .A(a[87]), .B(b[10]), .Z(n20376) );
  XOR U28868 ( .A(n20382), .B(n20383), .Z(n19805) );
  ANDN U28869 ( .B(n20384), .A(n20385), .Z(n20382) );
  AND U28870 ( .A(b[9]), .B(a[88]), .Z(n20381) );
  XOR U28871 ( .A(n20387), .B(n20388), .Z(n19810) );
  ANDN U28872 ( .B(n20389), .A(n20390), .Z(n20387) );
  AND U28873 ( .A(b[8]), .B(a[89]), .Z(n20386) );
  XOR U28874 ( .A(n20392), .B(n20393), .Z(n19815) );
  ANDN U28875 ( .B(n20394), .A(n20395), .Z(n20392) );
  AND U28876 ( .A(b[7]), .B(a[90]), .Z(n20391) );
  XOR U28877 ( .A(n20397), .B(n20398), .Z(n19820) );
  ANDN U28878 ( .B(n20399), .A(n20400), .Z(n20397) );
  AND U28879 ( .A(b[6]), .B(a[91]), .Z(n20396) );
  XOR U28880 ( .A(n20402), .B(n20403), .Z(n19825) );
  ANDN U28881 ( .B(n20404), .A(n20405), .Z(n20402) );
  AND U28882 ( .A(b[5]), .B(a[92]), .Z(n20401) );
  XOR U28883 ( .A(n20407), .B(n20408), .Z(n19830) );
  ANDN U28884 ( .B(n20409), .A(n20410), .Z(n20407) );
  AND U28885 ( .A(b[4]), .B(a[93]), .Z(n20406) );
  XOR U28886 ( .A(n20412), .B(n20413), .Z(n19835) );
  ANDN U28887 ( .B(n19847), .A(n19848), .Z(n20412) );
  AND U28888 ( .A(b[2]), .B(a[94]), .Z(n20414) );
  XNOR U28889 ( .A(n20409), .B(n20413), .Z(n20415) );
  XOR U28890 ( .A(n20416), .B(n20417), .Z(n20413) );
  OR U28891 ( .A(n19850), .B(n19851), .Z(n20417) );
  XNOR U28892 ( .A(n20419), .B(n20420), .Z(n20418) );
  XOR U28893 ( .A(n20419), .B(n20422), .Z(n19850) );
  NAND U28894 ( .A(b[1]), .B(a[94]), .Z(n20422) );
  IV U28895 ( .A(n20416), .Z(n20419) );
  NANDN U28896 ( .A(n13), .B(n14), .Z(n20416) );
  XOR U28897 ( .A(n20423), .B(n20424), .Z(n14) );
  NAND U28898 ( .A(a[94]), .B(b[0]), .Z(n13) );
  XNOR U28899 ( .A(n20404), .B(n20408), .Z(n20425) );
  XNOR U28900 ( .A(n20399), .B(n20403), .Z(n20426) );
  XNOR U28901 ( .A(n20394), .B(n20398), .Z(n20427) );
  XNOR U28902 ( .A(n20389), .B(n20393), .Z(n20428) );
  XNOR U28903 ( .A(n20384), .B(n20388), .Z(n20429) );
  XNOR U28904 ( .A(n20379), .B(n20383), .Z(n20430) );
  XNOR U28905 ( .A(n20374), .B(n20378), .Z(n20431) );
  XNOR U28906 ( .A(n20369), .B(n20373), .Z(n20432) );
  XNOR U28907 ( .A(n20364), .B(n20368), .Z(n20433) );
  XNOR U28908 ( .A(n20359), .B(n20363), .Z(n20434) );
  XNOR U28909 ( .A(n20354), .B(n20358), .Z(n20435) );
  XNOR U28910 ( .A(n20349), .B(n20353), .Z(n20436) );
  XNOR U28911 ( .A(n20344), .B(n20348), .Z(n20437) );
  XNOR U28912 ( .A(n20339), .B(n20343), .Z(n20438) );
  XNOR U28913 ( .A(n20334), .B(n20338), .Z(n20439) );
  XNOR U28914 ( .A(n20329), .B(n20333), .Z(n20440) );
  XNOR U28915 ( .A(n20324), .B(n20328), .Z(n20441) );
  XNOR U28916 ( .A(n20319), .B(n20323), .Z(n20442) );
  XNOR U28917 ( .A(n20314), .B(n20318), .Z(n20443) );
  XNOR U28918 ( .A(n20309), .B(n20313), .Z(n20444) );
  XNOR U28919 ( .A(n20304), .B(n20308), .Z(n20445) );
  XNOR U28920 ( .A(n20299), .B(n20303), .Z(n20446) );
  XNOR U28921 ( .A(n20294), .B(n20298), .Z(n20447) );
  XNOR U28922 ( .A(n20289), .B(n20293), .Z(n20448) );
  XNOR U28923 ( .A(n20284), .B(n20288), .Z(n20449) );
  XNOR U28924 ( .A(n20279), .B(n20283), .Z(n20450) );
  XNOR U28925 ( .A(n20274), .B(n20278), .Z(n20451) );
  XNOR U28926 ( .A(n20269), .B(n20273), .Z(n20452) );
  XNOR U28927 ( .A(n20264), .B(n20268), .Z(n20453) );
  XNOR U28928 ( .A(n20259), .B(n20263), .Z(n20454) );
  XNOR U28929 ( .A(n20254), .B(n20258), .Z(n20455) );
  XNOR U28930 ( .A(n20249), .B(n20253), .Z(n20456) );
  XNOR U28931 ( .A(n20244), .B(n20248), .Z(n20457) );
  XNOR U28932 ( .A(n20239), .B(n20243), .Z(n20458) );
  XNOR U28933 ( .A(n20234), .B(n20238), .Z(n20459) );
  XNOR U28934 ( .A(n20229), .B(n20233), .Z(n20460) );
  XNOR U28935 ( .A(n20224), .B(n20228), .Z(n20461) );
  XNOR U28936 ( .A(n20219), .B(n20223), .Z(n20462) );
  XNOR U28937 ( .A(n20214), .B(n20218), .Z(n20463) );
  XNOR U28938 ( .A(n20209), .B(n20213), .Z(n20464) );
  XNOR U28939 ( .A(n20204), .B(n20208), .Z(n20465) );
  XNOR U28940 ( .A(n20199), .B(n20203), .Z(n20466) );
  XNOR U28941 ( .A(n20194), .B(n20198), .Z(n20467) );
  XNOR U28942 ( .A(n20189), .B(n20193), .Z(n20468) );
  XNOR U28943 ( .A(n20184), .B(n20188), .Z(n20469) );
  XNOR U28944 ( .A(n20179), .B(n20183), .Z(n20470) );
  XNOR U28945 ( .A(n20174), .B(n20178), .Z(n20471) );
  XNOR U28946 ( .A(n20169), .B(n20173), .Z(n20472) );
  XNOR U28947 ( .A(n20164), .B(n20168), .Z(n20473) );
  XNOR U28948 ( .A(n20159), .B(n20163), .Z(n20474) );
  XNOR U28949 ( .A(n20154), .B(n20158), .Z(n20475) );
  XNOR U28950 ( .A(n20149), .B(n20153), .Z(n20476) );
  XNOR U28951 ( .A(n20144), .B(n20148), .Z(n20477) );
  XNOR U28952 ( .A(n20139), .B(n20143), .Z(n20478) );
  XNOR U28953 ( .A(n20134), .B(n20138), .Z(n20479) );
  XNOR U28954 ( .A(n20129), .B(n20133), .Z(n20480) );
  XNOR U28955 ( .A(n20124), .B(n20128), .Z(n20481) );
  XNOR U28956 ( .A(n20119), .B(n20123), .Z(n20482) );
  XNOR U28957 ( .A(n20114), .B(n20118), .Z(n20483) );
  XNOR U28958 ( .A(n20109), .B(n20113), .Z(n20484) );
  XNOR U28959 ( .A(n20104), .B(n20108), .Z(n20485) );
  XNOR U28960 ( .A(n20099), .B(n20103), .Z(n20486) );
  XNOR U28961 ( .A(n20094), .B(n20098), .Z(n20487) );
  XNOR U28962 ( .A(n20089), .B(n20093), .Z(n20488) );
  XNOR U28963 ( .A(n20084), .B(n20088), .Z(n20489) );
  XNOR U28964 ( .A(n20079), .B(n20083), .Z(n20490) );
  XNOR U28965 ( .A(n20074), .B(n20078), .Z(n20491) );
  XNOR U28966 ( .A(n20069), .B(n20073), .Z(n20492) );
  XNOR U28967 ( .A(n20064), .B(n20068), .Z(n20493) );
  XNOR U28968 ( .A(n20059), .B(n20063), .Z(n20494) );
  XNOR U28969 ( .A(n20054), .B(n20058), .Z(n20495) );
  XNOR U28970 ( .A(n20049), .B(n20053), .Z(n20496) );
  XNOR U28971 ( .A(n20044), .B(n20048), .Z(n20497) );
  XNOR U28972 ( .A(n20039), .B(n20043), .Z(n20498) );
  XNOR U28973 ( .A(n20034), .B(n20038), .Z(n20499) );
  XNOR U28974 ( .A(n20029), .B(n20033), .Z(n20500) );
  XNOR U28975 ( .A(n20024), .B(n20028), .Z(n20501) );
  XNOR U28976 ( .A(n20019), .B(n20023), .Z(n20502) );
  XNOR U28977 ( .A(n20014), .B(n20018), .Z(n20503) );
  XNOR U28978 ( .A(n20009), .B(n20013), .Z(n20504) );
  XNOR U28979 ( .A(n20004), .B(n20008), .Z(n20505) );
  XNOR U28980 ( .A(n19999), .B(n20003), .Z(n20506) );
  XNOR U28981 ( .A(n19994), .B(n19998), .Z(n20507) );
  XNOR U28982 ( .A(n19989), .B(n19993), .Z(n20508) );
  XNOR U28983 ( .A(n19984), .B(n19988), .Z(n20509) );
  XNOR U28984 ( .A(n19979), .B(n19983), .Z(n20510) );
  XNOR U28985 ( .A(n19974), .B(n19978), .Z(n20511) );
  XNOR U28986 ( .A(n19969), .B(n19973), .Z(n20512) );
  XNOR U28987 ( .A(n19964), .B(n19968), .Z(n20513) );
  XNOR U28988 ( .A(n19959), .B(n19963), .Z(n20514) );
  XNOR U28989 ( .A(n19954), .B(n19958), .Z(n20515) );
  XNOR U28990 ( .A(n19949), .B(n19953), .Z(n20516) );
  XOR U28991 ( .A(n20517), .B(n19948), .Z(n19949) );
  AND U28992 ( .A(a[0]), .B(b[96]), .Z(n20517) );
  XNOR U28993 ( .A(n20518), .B(n19948), .Z(n19950) );
  XNOR U28994 ( .A(n20519), .B(n20520), .Z(n19948) );
  ANDN U28995 ( .B(n20521), .A(n20522), .Z(n20519) );
  AND U28996 ( .A(a[1]), .B(b[95]), .Z(n20518) );
  XOR U28997 ( .A(n20524), .B(n20525), .Z(n19953) );
  ANDN U28998 ( .B(n20526), .A(n20527), .Z(n20524) );
  AND U28999 ( .A(a[2]), .B(b[94]), .Z(n20523) );
  XOR U29000 ( .A(n20529), .B(n20530), .Z(n19958) );
  ANDN U29001 ( .B(n20531), .A(n20532), .Z(n20529) );
  AND U29002 ( .A(a[3]), .B(b[93]), .Z(n20528) );
  XOR U29003 ( .A(n20534), .B(n20535), .Z(n19963) );
  ANDN U29004 ( .B(n20536), .A(n20537), .Z(n20534) );
  AND U29005 ( .A(a[4]), .B(b[92]), .Z(n20533) );
  XOR U29006 ( .A(n20539), .B(n20540), .Z(n19968) );
  ANDN U29007 ( .B(n20541), .A(n20542), .Z(n20539) );
  AND U29008 ( .A(a[5]), .B(b[91]), .Z(n20538) );
  XOR U29009 ( .A(n20544), .B(n20545), .Z(n19973) );
  ANDN U29010 ( .B(n20546), .A(n20547), .Z(n20544) );
  AND U29011 ( .A(a[6]), .B(b[90]), .Z(n20543) );
  XOR U29012 ( .A(n20549), .B(n20550), .Z(n19978) );
  ANDN U29013 ( .B(n20551), .A(n20552), .Z(n20549) );
  AND U29014 ( .A(a[7]), .B(b[89]), .Z(n20548) );
  XOR U29015 ( .A(n20554), .B(n20555), .Z(n19983) );
  ANDN U29016 ( .B(n20556), .A(n20557), .Z(n20554) );
  AND U29017 ( .A(a[8]), .B(b[88]), .Z(n20553) );
  XOR U29018 ( .A(n20559), .B(n20560), .Z(n19988) );
  ANDN U29019 ( .B(n20561), .A(n20562), .Z(n20559) );
  AND U29020 ( .A(a[9]), .B(b[87]), .Z(n20558) );
  XOR U29021 ( .A(n20564), .B(n20565), .Z(n19993) );
  ANDN U29022 ( .B(n20566), .A(n20567), .Z(n20564) );
  AND U29023 ( .A(a[10]), .B(b[86]), .Z(n20563) );
  XOR U29024 ( .A(n20569), .B(n20570), .Z(n19998) );
  ANDN U29025 ( .B(n20571), .A(n20572), .Z(n20569) );
  AND U29026 ( .A(a[11]), .B(b[85]), .Z(n20568) );
  XOR U29027 ( .A(n20574), .B(n20575), .Z(n20003) );
  ANDN U29028 ( .B(n20576), .A(n20577), .Z(n20574) );
  AND U29029 ( .A(a[12]), .B(b[84]), .Z(n20573) );
  XOR U29030 ( .A(n20579), .B(n20580), .Z(n20008) );
  ANDN U29031 ( .B(n20581), .A(n20582), .Z(n20579) );
  AND U29032 ( .A(a[13]), .B(b[83]), .Z(n20578) );
  XOR U29033 ( .A(n20584), .B(n20585), .Z(n20013) );
  ANDN U29034 ( .B(n20586), .A(n20587), .Z(n20584) );
  AND U29035 ( .A(a[14]), .B(b[82]), .Z(n20583) );
  XOR U29036 ( .A(n20589), .B(n20590), .Z(n20018) );
  ANDN U29037 ( .B(n20591), .A(n20592), .Z(n20589) );
  AND U29038 ( .A(a[15]), .B(b[81]), .Z(n20588) );
  XOR U29039 ( .A(n20594), .B(n20595), .Z(n20023) );
  ANDN U29040 ( .B(n20596), .A(n20597), .Z(n20594) );
  AND U29041 ( .A(a[16]), .B(b[80]), .Z(n20593) );
  XOR U29042 ( .A(n20599), .B(n20600), .Z(n20028) );
  ANDN U29043 ( .B(n20601), .A(n20602), .Z(n20599) );
  AND U29044 ( .A(a[17]), .B(b[79]), .Z(n20598) );
  XOR U29045 ( .A(n20604), .B(n20605), .Z(n20033) );
  ANDN U29046 ( .B(n20606), .A(n20607), .Z(n20604) );
  AND U29047 ( .A(a[18]), .B(b[78]), .Z(n20603) );
  XOR U29048 ( .A(n20609), .B(n20610), .Z(n20038) );
  ANDN U29049 ( .B(n20611), .A(n20612), .Z(n20609) );
  AND U29050 ( .A(a[19]), .B(b[77]), .Z(n20608) );
  XOR U29051 ( .A(n20614), .B(n20615), .Z(n20043) );
  ANDN U29052 ( .B(n20616), .A(n20617), .Z(n20614) );
  AND U29053 ( .A(a[20]), .B(b[76]), .Z(n20613) );
  XOR U29054 ( .A(n20619), .B(n20620), .Z(n20048) );
  ANDN U29055 ( .B(n20621), .A(n20622), .Z(n20619) );
  AND U29056 ( .A(a[21]), .B(b[75]), .Z(n20618) );
  XOR U29057 ( .A(n20624), .B(n20625), .Z(n20053) );
  ANDN U29058 ( .B(n20626), .A(n20627), .Z(n20624) );
  AND U29059 ( .A(a[22]), .B(b[74]), .Z(n20623) );
  XOR U29060 ( .A(n20629), .B(n20630), .Z(n20058) );
  ANDN U29061 ( .B(n20631), .A(n20632), .Z(n20629) );
  AND U29062 ( .A(a[23]), .B(b[73]), .Z(n20628) );
  XOR U29063 ( .A(n20634), .B(n20635), .Z(n20063) );
  ANDN U29064 ( .B(n20636), .A(n20637), .Z(n20634) );
  AND U29065 ( .A(a[24]), .B(b[72]), .Z(n20633) );
  XOR U29066 ( .A(n20639), .B(n20640), .Z(n20068) );
  ANDN U29067 ( .B(n20641), .A(n20642), .Z(n20639) );
  AND U29068 ( .A(a[25]), .B(b[71]), .Z(n20638) );
  XOR U29069 ( .A(n20644), .B(n20645), .Z(n20073) );
  ANDN U29070 ( .B(n20646), .A(n20647), .Z(n20644) );
  AND U29071 ( .A(a[26]), .B(b[70]), .Z(n20643) );
  XOR U29072 ( .A(n20649), .B(n20650), .Z(n20078) );
  ANDN U29073 ( .B(n20651), .A(n20652), .Z(n20649) );
  AND U29074 ( .A(a[27]), .B(b[69]), .Z(n20648) );
  XOR U29075 ( .A(n20654), .B(n20655), .Z(n20083) );
  ANDN U29076 ( .B(n20656), .A(n20657), .Z(n20654) );
  AND U29077 ( .A(a[28]), .B(b[68]), .Z(n20653) );
  XOR U29078 ( .A(n20659), .B(n20660), .Z(n20088) );
  ANDN U29079 ( .B(n20661), .A(n20662), .Z(n20659) );
  AND U29080 ( .A(a[29]), .B(b[67]), .Z(n20658) );
  XOR U29081 ( .A(n20664), .B(n20665), .Z(n20093) );
  ANDN U29082 ( .B(n20666), .A(n20667), .Z(n20664) );
  AND U29083 ( .A(a[30]), .B(b[66]), .Z(n20663) );
  XOR U29084 ( .A(n20669), .B(n20670), .Z(n20098) );
  ANDN U29085 ( .B(n20671), .A(n20672), .Z(n20669) );
  AND U29086 ( .A(a[31]), .B(b[65]), .Z(n20668) );
  XOR U29087 ( .A(n20674), .B(n20675), .Z(n20103) );
  ANDN U29088 ( .B(n20676), .A(n20677), .Z(n20674) );
  AND U29089 ( .A(a[32]), .B(b[64]), .Z(n20673) );
  XOR U29090 ( .A(n20679), .B(n20680), .Z(n20108) );
  ANDN U29091 ( .B(n20681), .A(n20682), .Z(n20679) );
  AND U29092 ( .A(a[33]), .B(b[63]), .Z(n20678) );
  XOR U29093 ( .A(n20684), .B(n20685), .Z(n20113) );
  ANDN U29094 ( .B(n20686), .A(n20687), .Z(n20684) );
  AND U29095 ( .A(a[34]), .B(b[62]), .Z(n20683) );
  XOR U29096 ( .A(n20689), .B(n20690), .Z(n20118) );
  ANDN U29097 ( .B(n20691), .A(n20692), .Z(n20689) );
  AND U29098 ( .A(a[35]), .B(b[61]), .Z(n20688) );
  XOR U29099 ( .A(n20694), .B(n20695), .Z(n20123) );
  ANDN U29100 ( .B(n20696), .A(n20697), .Z(n20694) );
  AND U29101 ( .A(a[36]), .B(b[60]), .Z(n20693) );
  XOR U29102 ( .A(n20699), .B(n20700), .Z(n20128) );
  ANDN U29103 ( .B(n20701), .A(n20702), .Z(n20699) );
  AND U29104 ( .A(a[37]), .B(b[59]), .Z(n20698) );
  XOR U29105 ( .A(n20704), .B(n20705), .Z(n20133) );
  ANDN U29106 ( .B(n20706), .A(n20707), .Z(n20704) );
  AND U29107 ( .A(a[38]), .B(b[58]), .Z(n20703) );
  XOR U29108 ( .A(n20709), .B(n20710), .Z(n20138) );
  ANDN U29109 ( .B(n20711), .A(n20712), .Z(n20709) );
  AND U29110 ( .A(a[39]), .B(b[57]), .Z(n20708) );
  XOR U29111 ( .A(n20714), .B(n20715), .Z(n20143) );
  ANDN U29112 ( .B(n20716), .A(n20717), .Z(n20714) );
  AND U29113 ( .A(a[40]), .B(b[56]), .Z(n20713) );
  XOR U29114 ( .A(n20719), .B(n20720), .Z(n20148) );
  ANDN U29115 ( .B(n20721), .A(n20722), .Z(n20719) );
  AND U29116 ( .A(a[41]), .B(b[55]), .Z(n20718) );
  XOR U29117 ( .A(n20724), .B(n20725), .Z(n20153) );
  ANDN U29118 ( .B(n20726), .A(n20727), .Z(n20724) );
  AND U29119 ( .A(a[42]), .B(b[54]), .Z(n20723) );
  XOR U29120 ( .A(n20729), .B(n20730), .Z(n20158) );
  ANDN U29121 ( .B(n20731), .A(n20732), .Z(n20729) );
  AND U29122 ( .A(a[43]), .B(b[53]), .Z(n20728) );
  XOR U29123 ( .A(n20734), .B(n20735), .Z(n20163) );
  ANDN U29124 ( .B(n20736), .A(n20737), .Z(n20734) );
  AND U29125 ( .A(a[44]), .B(b[52]), .Z(n20733) );
  XOR U29126 ( .A(n20739), .B(n20740), .Z(n20168) );
  ANDN U29127 ( .B(n20741), .A(n20742), .Z(n20739) );
  AND U29128 ( .A(a[45]), .B(b[51]), .Z(n20738) );
  XOR U29129 ( .A(n20744), .B(n20745), .Z(n20173) );
  ANDN U29130 ( .B(n20746), .A(n20747), .Z(n20744) );
  AND U29131 ( .A(a[46]), .B(b[50]), .Z(n20743) );
  XOR U29132 ( .A(n20749), .B(n20750), .Z(n20178) );
  ANDN U29133 ( .B(n20751), .A(n20752), .Z(n20749) );
  AND U29134 ( .A(a[47]), .B(b[49]), .Z(n20748) );
  XOR U29135 ( .A(n20754), .B(n20755), .Z(n20183) );
  ANDN U29136 ( .B(n20756), .A(n20757), .Z(n20754) );
  AND U29137 ( .A(a[48]), .B(b[48]), .Z(n20753) );
  XOR U29138 ( .A(n20759), .B(n20760), .Z(n20188) );
  ANDN U29139 ( .B(n20761), .A(n20762), .Z(n20759) );
  AND U29140 ( .A(a[49]), .B(b[47]), .Z(n20758) );
  XOR U29141 ( .A(n20764), .B(n20765), .Z(n20193) );
  ANDN U29142 ( .B(n20766), .A(n20767), .Z(n20764) );
  AND U29143 ( .A(a[50]), .B(b[46]), .Z(n20763) );
  XOR U29144 ( .A(n20769), .B(n20770), .Z(n20198) );
  ANDN U29145 ( .B(n20771), .A(n20772), .Z(n20769) );
  AND U29146 ( .A(a[51]), .B(b[45]), .Z(n20768) );
  XOR U29147 ( .A(n20774), .B(n20775), .Z(n20203) );
  ANDN U29148 ( .B(n20776), .A(n20777), .Z(n20774) );
  AND U29149 ( .A(a[52]), .B(b[44]), .Z(n20773) );
  XOR U29150 ( .A(n20779), .B(n20780), .Z(n20208) );
  ANDN U29151 ( .B(n20781), .A(n20782), .Z(n20779) );
  AND U29152 ( .A(a[53]), .B(b[43]), .Z(n20778) );
  XOR U29153 ( .A(n20784), .B(n20785), .Z(n20213) );
  ANDN U29154 ( .B(n20786), .A(n20787), .Z(n20784) );
  AND U29155 ( .A(a[54]), .B(b[42]), .Z(n20783) );
  XOR U29156 ( .A(n20789), .B(n20790), .Z(n20218) );
  ANDN U29157 ( .B(n20791), .A(n20792), .Z(n20789) );
  AND U29158 ( .A(a[55]), .B(b[41]), .Z(n20788) );
  XOR U29159 ( .A(n20794), .B(n20795), .Z(n20223) );
  ANDN U29160 ( .B(n20796), .A(n20797), .Z(n20794) );
  AND U29161 ( .A(a[56]), .B(b[40]), .Z(n20793) );
  XOR U29162 ( .A(n20799), .B(n20800), .Z(n20228) );
  ANDN U29163 ( .B(n20801), .A(n20802), .Z(n20799) );
  AND U29164 ( .A(a[57]), .B(b[39]), .Z(n20798) );
  XOR U29165 ( .A(n20804), .B(n20805), .Z(n20233) );
  ANDN U29166 ( .B(n20806), .A(n20807), .Z(n20804) );
  AND U29167 ( .A(a[58]), .B(b[38]), .Z(n20803) );
  XOR U29168 ( .A(n20809), .B(n20810), .Z(n20238) );
  ANDN U29169 ( .B(n20811), .A(n20812), .Z(n20809) );
  AND U29170 ( .A(a[59]), .B(b[37]), .Z(n20808) );
  XOR U29171 ( .A(n20814), .B(n20815), .Z(n20243) );
  ANDN U29172 ( .B(n20816), .A(n20817), .Z(n20814) );
  AND U29173 ( .A(a[60]), .B(b[36]), .Z(n20813) );
  XOR U29174 ( .A(n20819), .B(n20820), .Z(n20248) );
  ANDN U29175 ( .B(n20821), .A(n20822), .Z(n20819) );
  AND U29176 ( .A(a[61]), .B(b[35]), .Z(n20818) );
  XOR U29177 ( .A(n20824), .B(n20825), .Z(n20253) );
  ANDN U29178 ( .B(n20826), .A(n20827), .Z(n20824) );
  AND U29179 ( .A(a[62]), .B(b[34]), .Z(n20823) );
  XOR U29180 ( .A(n20829), .B(n20830), .Z(n20258) );
  ANDN U29181 ( .B(n20831), .A(n20832), .Z(n20829) );
  AND U29182 ( .A(a[63]), .B(b[33]), .Z(n20828) );
  XOR U29183 ( .A(n20834), .B(n20835), .Z(n20263) );
  ANDN U29184 ( .B(n20836), .A(n20837), .Z(n20834) );
  AND U29185 ( .A(a[64]), .B(b[32]), .Z(n20833) );
  XOR U29186 ( .A(n20839), .B(n20840), .Z(n20268) );
  ANDN U29187 ( .B(n20841), .A(n20842), .Z(n20839) );
  AND U29188 ( .A(a[65]), .B(b[31]), .Z(n20838) );
  XOR U29189 ( .A(n20844), .B(n20845), .Z(n20273) );
  ANDN U29190 ( .B(n20846), .A(n20847), .Z(n20844) );
  AND U29191 ( .A(a[66]), .B(b[30]), .Z(n20843) );
  XOR U29192 ( .A(n20849), .B(n20850), .Z(n20278) );
  ANDN U29193 ( .B(n20851), .A(n20852), .Z(n20849) );
  AND U29194 ( .A(a[67]), .B(b[29]), .Z(n20848) );
  XOR U29195 ( .A(n20854), .B(n20855), .Z(n20283) );
  ANDN U29196 ( .B(n20856), .A(n20857), .Z(n20854) );
  AND U29197 ( .A(a[68]), .B(b[28]), .Z(n20853) );
  XOR U29198 ( .A(n20859), .B(n20860), .Z(n20288) );
  ANDN U29199 ( .B(n20861), .A(n20862), .Z(n20859) );
  AND U29200 ( .A(a[69]), .B(b[27]), .Z(n20858) );
  XOR U29201 ( .A(n20864), .B(n20865), .Z(n20293) );
  ANDN U29202 ( .B(n20866), .A(n20867), .Z(n20864) );
  AND U29203 ( .A(a[70]), .B(b[26]), .Z(n20863) );
  XOR U29204 ( .A(n20869), .B(n20870), .Z(n20298) );
  ANDN U29205 ( .B(n20871), .A(n20872), .Z(n20869) );
  AND U29206 ( .A(a[71]), .B(b[25]), .Z(n20868) );
  XOR U29207 ( .A(n20874), .B(n20875), .Z(n20303) );
  ANDN U29208 ( .B(n20876), .A(n20877), .Z(n20874) );
  AND U29209 ( .A(a[72]), .B(b[24]), .Z(n20873) );
  XOR U29210 ( .A(n20879), .B(n20880), .Z(n20308) );
  ANDN U29211 ( .B(n20881), .A(n20882), .Z(n20879) );
  AND U29212 ( .A(a[73]), .B(b[23]), .Z(n20878) );
  XOR U29213 ( .A(n20884), .B(n20885), .Z(n20313) );
  ANDN U29214 ( .B(n20886), .A(n20887), .Z(n20884) );
  AND U29215 ( .A(a[74]), .B(b[22]), .Z(n20883) );
  XOR U29216 ( .A(n20889), .B(n20890), .Z(n20318) );
  ANDN U29217 ( .B(n20891), .A(n20892), .Z(n20889) );
  AND U29218 ( .A(a[75]), .B(b[21]), .Z(n20888) );
  XOR U29219 ( .A(n20894), .B(n20895), .Z(n20323) );
  ANDN U29220 ( .B(n20896), .A(n20897), .Z(n20894) );
  AND U29221 ( .A(a[76]), .B(b[20]), .Z(n20893) );
  XOR U29222 ( .A(n20899), .B(n20900), .Z(n20328) );
  ANDN U29223 ( .B(n20901), .A(n20902), .Z(n20899) );
  AND U29224 ( .A(a[77]), .B(b[19]), .Z(n20898) );
  XOR U29225 ( .A(n20904), .B(n20905), .Z(n20333) );
  ANDN U29226 ( .B(n20906), .A(n20907), .Z(n20904) );
  AND U29227 ( .A(a[78]), .B(b[18]), .Z(n20903) );
  XOR U29228 ( .A(n20909), .B(n20910), .Z(n20338) );
  ANDN U29229 ( .B(n20911), .A(n20912), .Z(n20909) );
  AND U29230 ( .A(a[79]), .B(b[17]), .Z(n20908) );
  XOR U29231 ( .A(n20914), .B(n20915), .Z(n20343) );
  ANDN U29232 ( .B(n20916), .A(n20917), .Z(n20914) );
  AND U29233 ( .A(a[80]), .B(b[16]), .Z(n20913) );
  XOR U29234 ( .A(n20919), .B(n20920), .Z(n20348) );
  ANDN U29235 ( .B(n20921), .A(n20922), .Z(n20919) );
  AND U29236 ( .A(a[81]), .B(b[15]), .Z(n20918) );
  XOR U29237 ( .A(n20924), .B(n20925), .Z(n20353) );
  ANDN U29238 ( .B(n20926), .A(n20927), .Z(n20924) );
  AND U29239 ( .A(a[82]), .B(b[14]), .Z(n20923) );
  XOR U29240 ( .A(n20929), .B(n20930), .Z(n20358) );
  ANDN U29241 ( .B(n20931), .A(n20932), .Z(n20929) );
  AND U29242 ( .A(a[83]), .B(b[13]), .Z(n20928) );
  XOR U29243 ( .A(n20934), .B(n20935), .Z(n20363) );
  ANDN U29244 ( .B(n20936), .A(n20937), .Z(n20934) );
  AND U29245 ( .A(a[84]), .B(b[12]), .Z(n20933) );
  XOR U29246 ( .A(n20939), .B(n20940), .Z(n20368) );
  ANDN U29247 ( .B(n20941), .A(n20942), .Z(n20939) );
  AND U29248 ( .A(a[85]), .B(b[11]), .Z(n20938) );
  XOR U29249 ( .A(n20944), .B(n20945), .Z(n20373) );
  ANDN U29250 ( .B(n20946), .A(n20947), .Z(n20944) );
  AND U29251 ( .A(a[86]), .B(b[10]), .Z(n20943) );
  XOR U29252 ( .A(n20949), .B(n20950), .Z(n20378) );
  ANDN U29253 ( .B(n20951), .A(n20952), .Z(n20949) );
  AND U29254 ( .A(b[9]), .B(a[87]), .Z(n20948) );
  XOR U29255 ( .A(n20954), .B(n20955), .Z(n20383) );
  ANDN U29256 ( .B(n20956), .A(n20957), .Z(n20954) );
  AND U29257 ( .A(b[8]), .B(a[88]), .Z(n20953) );
  XOR U29258 ( .A(n20959), .B(n20960), .Z(n20388) );
  ANDN U29259 ( .B(n20961), .A(n20962), .Z(n20959) );
  AND U29260 ( .A(b[7]), .B(a[89]), .Z(n20958) );
  XOR U29261 ( .A(n20964), .B(n20965), .Z(n20393) );
  ANDN U29262 ( .B(n20966), .A(n20967), .Z(n20964) );
  AND U29263 ( .A(b[6]), .B(a[90]), .Z(n20963) );
  XOR U29264 ( .A(n20969), .B(n20970), .Z(n20398) );
  ANDN U29265 ( .B(n20971), .A(n20972), .Z(n20969) );
  AND U29266 ( .A(b[5]), .B(a[91]), .Z(n20968) );
  XOR U29267 ( .A(n20974), .B(n20975), .Z(n20403) );
  ANDN U29268 ( .B(n20976), .A(n20977), .Z(n20974) );
  AND U29269 ( .A(b[4]), .B(a[92]), .Z(n20973) );
  XOR U29270 ( .A(n20979), .B(n20980), .Z(n20408) );
  ANDN U29271 ( .B(n20420), .A(n20421), .Z(n20979) );
  AND U29272 ( .A(b[2]), .B(a[93]), .Z(n20981) );
  XNOR U29273 ( .A(n20976), .B(n20980), .Z(n20982) );
  XOR U29274 ( .A(n20983), .B(n20984), .Z(n20980) );
  OR U29275 ( .A(n20423), .B(n20424), .Z(n20984) );
  XNOR U29276 ( .A(n20986), .B(n20987), .Z(n20985) );
  XOR U29277 ( .A(n20986), .B(n20989), .Z(n20423) );
  NAND U29278 ( .A(b[1]), .B(a[93]), .Z(n20989) );
  IV U29279 ( .A(n20983), .Z(n20986) );
  NANDN U29280 ( .A(n15), .B(n16), .Z(n20983) );
  XOR U29281 ( .A(n20990), .B(n20991), .Z(n16) );
  NAND U29282 ( .A(a[93]), .B(b[0]), .Z(n15) );
  XNOR U29283 ( .A(n20971), .B(n20975), .Z(n20992) );
  XNOR U29284 ( .A(n20966), .B(n20970), .Z(n20993) );
  XNOR U29285 ( .A(n20961), .B(n20965), .Z(n20994) );
  XNOR U29286 ( .A(n20956), .B(n20960), .Z(n20995) );
  XNOR U29287 ( .A(n20951), .B(n20955), .Z(n20996) );
  XNOR U29288 ( .A(n20946), .B(n20950), .Z(n20997) );
  XNOR U29289 ( .A(n20941), .B(n20945), .Z(n20998) );
  XNOR U29290 ( .A(n20936), .B(n20940), .Z(n20999) );
  XNOR U29291 ( .A(n20931), .B(n20935), .Z(n21000) );
  XNOR U29292 ( .A(n20926), .B(n20930), .Z(n21001) );
  XNOR U29293 ( .A(n20921), .B(n20925), .Z(n21002) );
  XNOR U29294 ( .A(n20916), .B(n20920), .Z(n21003) );
  XNOR U29295 ( .A(n20911), .B(n20915), .Z(n21004) );
  XNOR U29296 ( .A(n20906), .B(n20910), .Z(n21005) );
  XNOR U29297 ( .A(n20901), .B(n20905), .Z(n21006) );
  XNOR U29298 ( .A(n20896), .B(n20900), .Z(n21007) );
  XNOR U29299 ( .A(n20891), .B(n20895), .Z(n21008) );
  XNOR U29300 ( .A(n20886), .B(n20890), .Z(n21009) );
  XNOR U29301 ( .A(n20881), .B(n20885), .Z(n21010) );
  XNOR U29302 ( .A(n20876), .B(n20880), .Z(n21011) );
  XNOR U29303 ( .A(n20871), .B(n20875), .Z(n21012) );
  XNOR U29304 ( .A(n20866), .B(n20870), .Z(n21013) );
  XNOR U29305 ( .A(n20861), .B(n20865), .Z(n21014) );
  XNOR U29306 ( .A(n20856), .B(n20860), .Z(n21015) );
  XNOR U29307 ( .A(n20851), .B(n20855), .Z(n21016) );
  XNOR U29308 ( .A(n20846), .B(n20850), .Z(n21017) );
  XNOR U29309 ( .A(n20841), .B(n20845), .Z(n21018) );
  XNOR U29310 ( .A(n20836), .B(n20840), .Z(n21019) );
  XNOR U29311 ( .A(n20831), .B(n20835), .Z(n21020) );
  XNOR U29312 ( .A(n20826), .B(n20830), .Z(n21021) );
  XNOR U29313 ( .A(n20821), .B(n20825), .Z(n21022) );
  XNOR U29314 ( .A(n20816), .B(n20820), .Z(n21023) );
  XNOR U29315 ( .A(n20811), .B(n20815), .Z(n21024) );
  XNOR U29316 ( .A(n20806), .B(n20810), .Z(n21025) );
  XNOR U29317 ( .A(n20801), .B(n20805), .Z(n21026) );
  XNOR U29318 ( .A(n20796), .B(n20800), .Z(n21027) );
  XNOR U29319 ( .A(n20791), .B(n20795), .Z(n21028) );
  XNOR U29320 ( .A(n20786), .B(n20790), .Z(n21029) );
  XNOR U29321 ( .A(n20781), .B(n20785), .Z(n21030) );
  XNOR U29322 ( .A(n20776), .B(n20780), .Z(n21031) );
  XNOR U29323 ( .A(n20771), .B(n20775), .Z(n21032) );
  XNOR U29324 ( .A(n20766), .B(n20770), .Z(n21033) );
  XNOR U29325 ( .A(n20761), .B(n20765), .Z(n21034) );
  XNOR U29326 ( .A(n20756), .B(n20760), .Z(n21035) );
  XNOR U29327 ( .A(n20751), .B(n20755), .Z(n21036) );
  XNOR U29328 ( .A(n20746), .B(n20750), .Z(n21037) );
  XNOR U29329 ( .A(n20741), .B(n20745), .Z(n21038) );
  XNOR U29330 ( .A(n20736), .B(n20740), .Z(n21039) );
  XNOR U29331 ( .A(n20731), .B(n20735), .Z(n21040) );
  XNOR U29332 ( .A(n20726), .B(n20730), .Z(n21041) );
  XNOR U29333 ( .A(n20721), .B(n20725), .Z(n21042) );
  XNOR U29334 ( .A(n20716), .B(n20720), .Z(n21043) );
  XNOR U29335 ( .A(n20711), .B(n20715), .Z(n21044) );
  XNOR U29336 ( .A(n20706), .B(n20710), .Z(n21045) );
  XNOR U29337 ( .A(n20701), .B(n20705), .Z(n21046) );
  XNOR U29338 ( .A(n21047), .B(n21048), .Z(n20701) );
  XNOR U29339 ( .A(n20696), .B(n20700), .Z(n21048) );
  XNOR U29340 ( .A(n20691), .B(n20695), .Z(n21049) );
  XNOR U29341 ( .A(n20686), .B(n20690), .Z(n21050) );
  XNOR U29342 ( .A(n20681), .B(n20685), .Z(n21051) );
  XNOR U29343 ( .A(n20676), .B(n20680), .Z(n21052) );
  XNOR U29344 ( .A(n20671), .B(n20675), .Z(n21053) );
  XNOR U29345 ( .A(n20666), .B(n20670), .Z(n21054) );
  XNOR U29346 ( .A(n20661), .B(n20665), .Z(n21055) );
  XNOR U29347 ( .A(n20656), .B(n20660), .Z(n21056) );
  XNOR U29348 ( .A(n20651), .B(n20655), .Z(n21057) );
  XNOR U29349 ( .A(n20646), .B(n20650), .Z(n21058) );
  XNOR U29350 ( .A(n20641), .B(n20645), .Z(n21059) );
  XNOR U29351 ( .A(n20636), .B(n20640), .Z(n21060) );
  XNOR U29352 ( .A(n20631), .B(n20635), .Z(n21061) );
  XNOR U29353 ( .A(n20626), .B(n20630), .Z(n21062) );
  XNOR U29354 ( .A(n20621), .B(n20625), .Z(n21063) );
  XNOR U29355 ( .A(n20616), .B(n20620), .Z(n21064) );
  XNOR U29356 ( .A(n20611), .B(n20615), .Z(n21065) );
  XNOR U29357 ( .A(n20606), .B(n20610), .Z(n21066) );
  XNOR U29358 ( .A(n20601), .B(n20605), .Z(n21067) );
  XNOR U29359 ( .A(n20596), .B(n20600), .Z(n21068) );
  XNOR U29360 ( .A(n20591), .B(n20595), .Z(n21069) );
  XNOR U29361 ( .A(n20586), .B(n20590), .Z(n21070) );
  XNOR U29362 ( .A(n20581), .B(n20585), .Z(n21071) );
  XNOR U29363 ( .A(n20576), .B(n20580), .Z(n21072) );
  XNOR U29364 ( .A(n20571), .B(n20575), .Z(n21073) );
  XNOR U29365 ( .A(n20566), .B(n20570), .Z(n21074) );
  XNOR U29366 ( .A(n20561), .B(n20565), .Z(n21075) );
  XNOR U29367 ( .A(n20556), .B(n20560), .Z(n21076) );
  XNOR U29368 ( .A(n20551), .B(n20555), .Z(n21077) );
  XNOR U29369 ( .A(n20546), .B(n20550), .Z(n21078) );
  XNOR U29370 ( .A(n20541), .B(n20545), .Z(n21079) );
  XNOR U29371 ( .A(n20536), .B(n20540), .Z(n21080) );
  XNOR U29372 ( .A(n20531), .B(n20535), .Z(n21081) );
  XNOR U29373 ( .A(n20526), .B(n20530), .Z(n21082) );
  XNOR U29374 ( .A(n20521), .B(n20525), .Z(n21083) );
  XNOR U29375 ( .A(n21084), .B(n20520), .Z(n20521) );
  AND U29376 ( .A(a[0]), .B(b[95]), .Z(n21084) );
  XOR U29377 ( .A(n21085), .B(n20520), .Z(n20522) );
  XNOR U29378 ( .A(n21086), .B(n21087), .Z(n20520) );
  ANDN U29379 ( .B(n21088), .A(n21089), .Z(n21086) );
  AND U29380 ( .A(a[1]), .B(b[94]), .Z(n21085) );
  XOR U29381 ( .A(n21091), .B(n21092), .Z(n20525) );
  ANDN U29382 ( .B(n21093), .A(n21094), .Z(n21091) );
  AND U29383 ( .A(a[2]), .B(b[93]), .Z(n21090) );
  XOR U29384 ( .A(n21096), .B(n21097), .Z(n20530) );
  ANDN U29385 ( .B(n21098), .A(n21099), .Z(n21096) );
  AND U29386 ( .A(a[3]), .B(b[92]), .Z(n21095) );
  XOR U29387 ( .A(n21101), .B(n21102), .Z(n20535) );
  ANDN U29388 ( .B(n21103), .A(n21104), .Z(n21101) );
  AND U29389 ( .A(a[4]), .B(b[91]), .Z(n21100) );
  XOR U29390 ( .A(n21106), .B(n21107), .Z(n20540) );
  ANDN U29391 ( .B(n21108), .A(n21109), .Z(n21106) );
  AND U29392 ( .A(a[5]), .B(b[90]), .Z(n21105) );
  XOR U29393 ( .A(n21111), .B(n21112), .Z(n20545) );
  ANDN U29394 ( .B(n21113), .A(n21114), .Z(n21111) );
  AND U29395 ( .A(a[6]), .B(b[89]), .Z(n21110) );
  XOR U29396 ( .A(n21116), .B(n21117), .Z(n20550) );
  ANDN U29397 ( .B(n21118), .A(n21119), .Z(n21116) );
  AND U29398 ( .A(a[7]), .B(b[88]), .Z(n21115) );
  XOR U29399 ( .A(n21121), .B(n21122), .Z(n20555) );
  ANDN U29400 ( .B(n21123), .A(n21124), .Z(n21121) );
  AND U29401 ( .A(a[8]), .B(b[87]), .Z(n21120) );
  XOR U29402 ( .A(n21126), .B(n21127), .Z(n20560) );
  ANDN U29403 ( .B(n21128), .A(n21129), .Z(n21126) );
  AND U29404 ( .A(a[9]), .B(b[86]), .Z(n21125) );
  XOR U29405 ( .A(n21131), .B(n21132), .Z(n20565) );
  ANDN U29406 ( .B(n21133), .A(n21134), .Z(n21131) );
  AND U29407 ( .A(a[10]), .B(b[85]), .Z(n21130) );
  XOR U29408 ( .A(n21136), .B(n21137), .Z(n20570) );
  ANDN U29409 ( .B(n21138), .A(n21139), .Z(n21136) );
  AND U29410 ( .A(a[11]), .B(b[84]), .Z(n21135) );
  XOR U29411 ( .A(n21141), .B(n21142), .Z(n20575) );
  ANDN U29412 ( .B(n21143), .A(n21144), .Z(n21141) );
  AND U29413 ( .A(a[12]), .B(b[83]), .Z(n21140) );
  XOR U29414 ( .A(n21146), .B(n21147), .Z(n20580) );
  ANDN U29415 ( .B(n21148), .A(n21149), .Z(n21146) );
  AND U29416 ( .A(a[13]), .B(b[82]), .Z(n21145) );
  XOR U29417 ( .A(n21151), .B(n21152), .Z(n20585) );
  ANDN U29418 ( .B(n21153), .A(n21154), .Z(n21151) );
  AND U29419 ( .A(a[14]), .B(b[81]), .Z(n21150) );
  XOR U29420 ( .A(n21156), .B(n21157), .Z(n20590) );
  ANDN U29421 ( .B(n21158), .A(n21159), .Z(n21156) );
  AND U29422 ( .A(a[15]), .B(b[80]), .Z(n21155) );
  XOR U29423 ( .A(n21161), .B(n21162), .Z(n20595) );
  ANDN U29424 ( .B(n21163), .A(n21164), .Z(n21161) );
  AND U29425 ( .A(a[16]), .B(b[79]), .Z(n21160) );
  XOR U29426 ( .A(n21166), .B(n21167), .Z(n20600) );
  ANDN U29427 ( .B(n21168), .A(n21169), .Z(n21166) );
  AND U29428 ( .A(a[17]), .B(b[78]), .Z(n21165) );
  XOR U29429 ( .A(n21171), .B(n21172), .Z(n20605) );
  ANDN U29430 ( .B(n21173), .A(n21174), .Z(n21171) );
  AND U29431 ( .A(a[18]), .B(b[77]), .Z(n21170) );
  XOR U29432 ( .A(n21176), .B(n21177), .Z(n20610) );
  ANDN U29433 ( .B(n21178), .A(n21179), .Z(n21176) );
  AND U29434 ( .A(a[19]), .B(b[76]), .Z(n21175) );
  XOR U29435 ( .A(n21181), .B(n21182), .Z(n20615) );
  ANDN U29436 ( .B(n21183), .A(n21184), .Z(n21181) );
  AND U29437 ( .A(a[20]), .B(b[75]), .Z(n21180) );
  XOR U29438 ( .A(n21186), .B(n21187), .Z(n20620) );
  ANDN U29439 ( .B(n21188), .A(n21189), .Z(n21186) );
  AND U29440 ( .A(a[21]), .B(b[74]), .Z(n21185) );
  XOR U29441 ( .A(n21191), .B(n21192), .Z(n20625) );
  ANDN U29442 ( .B(n21193), .A(n21194), .Z(n21191) );
  AND U29443 ( .A(a[22]), .B(b[73]), .Z(n21190) );
  XOR U29444 ( .A(n21196), .B(n21197), .Z(n20630) );
  ANDN U29445 ( .B(n21198), .A(n21199), .Z(n21196) );
  AND U29446 ( .A(a[23]), .B(b[72]), .Z(n21195) );
  XOR U29447 ( .A(n21201), .B(n21202), .Z(n20635) );
  ANDN U29448 ( .B(n21203), .A(n21204), .Z(n21201) );
  AND U29449 ( .A(a[24]), .B(b[71]), .Z(n21200) );
  XOR U29450 ( .A(n21206), .B(n21207), .Z(n20640) );
  ANDN U29451 ( .B(n21208), .A(n21209), .Z(n21206) );
  AND U29452 ( .A(a[25]), .B(b[70]), .Z(n21205) );
  XOR U29453 ( .A(n21211), .B(n21212), .Z(n20645) );
  ANDN U29454 ( .B(n21213), .A(n21214), .Z(n21211) );
  AND U29455 ( .A(a[26]), .B(b[69]), .Z(n21210) );
  XOR U29456 ( .A(n21216), .B(n21217), .Z(n20650) );
  ANDN U29457 ( .B(n21218), .A(n21219), .Z(n21216) );
  AND U29458 ( .A(a[27]), .B(b[68]), .Z(n21215) );
  XOR U29459 ( .A(n21221), .B(n21222), .Z(n20655) );
  ANDN U29460 ( .B(n21223), .A(n21224), .Z(n21221) );
  AND U29461 ( .A(a[28]), .B(b[67]), .Z(n21220) );
  XOR U29462 ( .A(n21226), .B(n21227), .Z(n20660) );
  ANDN U29463 ( .B(n21228), .A(n21229), .Z(n21226) );
  AND U29464 ( .A(a[29]), .B(b[66]), .Z(n21225) );
  XOR U29465 ( .A(n21231), .B(n21232), .Z(n20665) );
  ANDN U29466 ( .B(n21233), .A(n21234), .Z(n21231) );
  AND U29467 ( .A(a[30]), .B(b[65]), .Z(n21230) );
  XOR U29468 ( .A(n21236), .B(n21237), .Z(n20670) );
  ANDN U29469 ( .B(n21238), .A(n21239), .Z(n21236) );
  AND U29470 ( .A(a[31]), .B(b[64]), .Z(n21235) );
  XOR U29471 ( .A(n21241), .B(n21242), .Z(n20675) );
  ANDN U29472 ( .B(n21243), .A(n21244), .Z(n21241) );
  AND U29473 ( .A(a[32]), .B(b[63]), .Z(n21240) );
  XOR U29474 ( .A(n21246), .B(n21247), .Z(n20680) );
  ANDN U29475 ( .B(n21248), .A(n21249), .Z(n21246) );
  AND U29476 ( .A(a[33]), .B(b[62]), .Z(n21245) );
  XOR U29477 ( .A(n21251), .B(n21252), .Z(n20685) );
  ANDN U29478 ( .B(n21253), .A(n21254), .Z(n21251) );
  AND U29479 ( .A(a[34]), .B(b[61]), .Z(n21250) );
  XOR U29480 ( .A(n21256), .B(n21257), .Z(n20690) );
  ANDN U29481 ( .B(n21258), .A(n21259), .Z(n21256) );
  AND U29482 ( .A(a[35]), .B(b[60]), .Z(n21255) );
  IV U29483 ( .A(n20697), .Z(n21047) );
  XOR U29484 ( .A(n21261), .B(n21262), .Z(n20695) );
  ANDN U29485 ( .B(n21263), .A(n21264), .Z(n21261) );
  AND U29486 ( .A(a[36]), .B(b[59]), .Z(n21260) );
  XOR U29487 ( .A(n21266), .B(n21267), .Z(n20700) );
  ANDN U29488 ( .B(n21268), .A(n21269), .Z(n21266) );
  AND U29489 ( .A(a[37]), .B(b[58]), .Z(n21265) );
  XOR U29490 ( .A(n21271), .B(n21272), .Z(n20705) );
  ANDN U29491 ( .B(n21273), .A(n21274), .Z(n21271) );
  AND U29492 ( .A(a[38]), .B(b[57]), .Z(n21270) );
  XOR U29493 ( .A(n21276), .B(n21277), .Z(n20710) );
  ANDN U29494 ( .B(n21278), .A(n21279), .Z(n21276) );
  AND U29495 ( .A(a[39]), .B(b[56]), .Z(n21275) );
  XOR U29496 ( .A(n21281), .B(n21282), .Z(n20715) );
  ANDN U29497 ( .B(n21283), .A(n21284), .Z(n21281) );
  AND U29498 ( .A(a[40]), .B(b[55]), .Z(n21280) );
  XOR U29499 ( .A(n21286), .B(n21287), .Z(n20720) );
  ANDN U29500 ( .B(n21288), .A(n21289), .Z(n21286) );
  AND U29501 ( .A(a[41]), .B(b[54]), .Z(n21285) );
  XOR U29502 ( .A(n21291), .B(n21292), .Z(n20725) );
  ANDN U29503 ( .B(n21293), .A(n21294), .Z(n21291) );
  AND U29504 ( .A(a[42]), .B(b[53]), .Z(n21290) );
  XOR U29505 ( .A(n21296), .B(n21297), .Z(n20730) );
  ANDN U29506 ( .B(n21298), .A(n21299), .Z(n21296) );
  AND U29507 ( .A(a[43]), .B(b[52]), .Z(n21295) );
  XOR U29508 ( .A(n21301), .B(n21302), .Z(n20735) );
  ANDN U29509 ( .B(n21303), .A(n21304), .Z(n21301) );
  AND U29510 ( .A(a[44]), .B(b[51]), .Z(n21300) );
  XOR U29511 ( .A(n21306), .B(n21307), .Z(n20740) );
  ANDN U29512 ( .B(n21308), .A(n21309), .Z(n21306) );
  AND U29513 ( .A(a[45]), .B(b[50]), .Z(n21305) );
  XOR U29514 ( .A(n21311), .B(n21312), .Z(n20745) );
  ANDN U29515 ( .B(n21313), .A(n21314), .Z(n21311) );
  AND U29516 ( .A(a[46]), .B(b[49]), .Z(n21310) );
  XOR U29517 ( .A(n21316), .B(n21317), .Z(n20750) );
  ANDN U29518 ( .B(n21318), .A(n21319), .Z(n21316) );
  AND U29519 ( .A(a[47]), .B(b[48]), .Z(n21315) );
  XOR U29520 ( .A(n21321), .B(n21322), .Z(n20755) );
  ANDN U29521 ( .B(n21323), .A(n21324), .Z(n21321) );
  AND U29522 ( .A(a[48]), .B(b[47]), .Z(n21320) );
  XOR U29523 ( .A(n21326), .B(n21327), .Z(n20760) );
  ANDN U29524 ( .B(n21328), .A(n21329), .Z(n21326) );
  AND U29525 ( .A(a[49]), .B(b[46]), .Z(n21325) );
  XOR U29526 ( .A(n21331), .B(n21332), .Z(n20765) );
  ANDN U29527 ( .B(n21333), .A(n21334), .Z(n21331) );
  AND U29528 ( .A(a[50]), .B(b[45]), .Z(n21330) );
  XOR U29529 ( .A(n21336), .B(n21337), .Z(n20770) );
  ANDN U29530 ( .B(n21338), .A(n21339), .Z(n21336) );
  AND U29531 ( .A(a[51]), .B(b[44]), .Z(n21335) );
  XOR U29532 ( .A(n21341), .B(n21342), .Z(n20775) );
  ANDN U29533 ( .B(n21343), .A(n21344), .Z(n21341) );
  AND U29534 ( .A(a[52]), .B(b[43]), .Z(n21340) );
  XOR U29535 ( .A(n21346), .B(n21347), .Z(n20780) );
  ANDN U29536 ( .B(n21348), .A(n21349), .Z(n21346) );
  AND U29537 ( .A(a[53]), .B(b[42]), .Z(n21345) );
  XOR U29538 ( .A(n21351), .B(n21352), .Z(n20785) );
  ANDN U29539 ( .B(n21353), .A(n21354), .Z(n21351) );
  AND U29540 ( .A(a[54]), .B(b[41]), .Z(n21350) );
  XOR U29541 ( .A(n21356), .B(n21357), .Z(n20790) );
  ANDN U29542 ( .B(n21358), .A(n21359), .Z(n21356) );
  AND U29543 ( .A(a[55]), .B(b[40]), .Z(n21355) );
  XOR U29544 ( .A(n21361), .B(n21362), .Z(n20795) );
  ANDN U29545 ( .B(n21363), .A(n21364), .Z(n21361) );
  AND U29546 ( .A(a[56]), .B(b[39]), .Z(n21360) );
  XOR U29547 ( .A(n21366), .B(n21367), .Z(n20800) );
  ANDN U29548 ( .B(n21368), .A(n21369), .Z(n21366) );
  AND U29549 ( .A(a[57]), .B(b[38]), .Z(n21365) );
  XOR U29550 ( .A(n21371), .B(n21372), .Z(n20805) );
  ANDN U29551 ( .B(n21373), .A(n21374), .Z(n21371) );
  AND U29552 ( .A(a[58]), .B(b[37]), .Z(n21370) );
  XOR U29553 ( .A(n21376), .B(n21377), .Z(n20810) );
  ANDN U29554 ( .B(n21378), .A(n21379), .Z(n21376) );
  AND U29555 ( .A(a[59]), .B(b[36]), .Z(n21375) );
  XOR U29556 ( .A(n21381), .B(n21382), .Z(n20815) );
  ANDN U29557 ( .B(n21383), .A(n21384), .Z(n21381) );
  AND U29558 ( .A(a[60]), .B(b[35]), .Z(n21380) );
  XOR U29559 ( .A(n21386), .B(n21387), .Z(n20820) );
  ANDN U29560 ( .B(n21388), .A(n21389), .Z(n21386) );
  AND U29561 ( .A(a[61]), .B(b[34]), .Z(n21385) );
  XOR U29562 ( .A(n21391), .B(n21392), .Z(n20825) );
  ANDN U29563 ( .B(n21393), .A(n21394), .Z(n21391) );
  AND U29564 ( .A(a[62]), .B(b[33]), .Z(n21390) );
  XOR U29565 ( .A(n21396), .B(n21397), .Z(n20830) );
  ANDN U29566 ( .B(n21398), .A(n21399), .Z(n21396) );
  AND U29567 ( .A(a[63]), .B(b[32]), .Z(n21395) );
  XOR U29568 ( .A(n21401), .B(n21402), .Z(n20835) );
  ANDN U29569 ( .B(n21403), .A(n21404), .Z(n21401) );
  AND U29570 ( .A(a[64]), .B(b[31]), .Z(n21400) );
  XOR U29571 ( .A(n21406), .B(n21407), .Z(n20840) );
  ANDN U29572 ( .B(n21408), .A(n21409), .Z(n21406) );
  AND U29573 ( .A(a[65]), .B(b[30]), .Z(n21405) );
  XOR U29574 ( .A(n21411), .B(n21412), .Z(n20845) );
  ANDN U29575 ( .B(n21413), .A(n21414), .Z(n21411) );
  AND U29576 ( .A(a[66]), .B(b[29]), .Z(n21410) );
  XOR U29577 ( .A(n21416), .B(n21417), .Z(n20850) );
  ANDN U29578 ( .B(n21418), .A(n21419), .Z(n21416) );
  AND U29579 ( .A(a[67]), .B(b[28]), .Z(n21415) );
  XOR U29580 ( .A(n21421), .B(n21422), .Z(n20855) );
  ANDN U29581 ( .B(n21423), .A(n21424), .Z(n21421) );
  AND U29582 ( .A(a[68]), .B(b[27]), .Z(n21420) );
  XOR U29583 ( .A(n21426), .B(n21427), .Z(n20860) );
  ANDN U29584 ( .B(n21428), .A(n21429), .Z(n21426) );
  AND U29585 ( .A(a[69]), .B(b[26]), .Z(n21425) );
  XOR U29586 ( .A(n21431), .B(n21432), .Z(n20865) );
  ANDN U29587 ( .B(n21433), .A(n21434), .Z(n21431) );
  AND U29588 ( .A(a[70]), .B(b[25]), .Z(n21430) );
  XOR U29589 ( .A(n21436), .B(n21437), .Z(n20870) );
  ANDN U29590 ( .B(n21438), .A(n21439), .Z(n21436) );
  AND U29591 ( .A(a[71]), .B(b[24]), .Z(n21435) );
  XOR U29592 ( .A(n21441), .B(n21442), .Z(n20875) );
  ANDN U29593 ( .B(n21443), .A(n21444), .Z(n21441) );
  AND U29594 ( .A(a[72]), .B(b[23]), .Z(n21440) );
  XOR U29595 ( .A(n21446), .B(n21447), .Z(n20880) );
  ANDN U29596 ( .B(n21448), .A(n21449), .Z(n21446) );
  AND U29597 ( .A(a[73]), .B(b[22]), .Z(n21445) );
  XOR U29598 ( .A(n21451), .B(n21452), .Z(n20885) );
  ANDN U29599 ( .B(n21453), .A(n21454), .Z(n21451) );
  AND U29600 ( .A(a[74]), .B(b[21]), .Z(n21450) );
  XOR U29601 ( .A(n21456), .B(n21457), .Z(n20890) );
  ANDN U29602 ( .B(n21458), .A(n21459), .Z(n21456) );
  AND U29603 ( .A(a[75]), .B(b[20]), .Z(n21455) );
  XOR U29604 ( .A(n21461), .B(n21462), .Z(n20895) );
  ANDN U29605 ( .B(n21463), .A(n21464), .Z(n21461) );
  AND U29606 ( .A(a[76]), .B(b[19]), .Z(n21460) );
  XOR U29607 ( .A(n21466), .B(n21467), .Z(n20900) );
  ANDN U29608 ( .B(n21468), .A(n21469), .Z(n21466) );
  AND U29609 ( .A(a[77]), .B(b[18]), .Z(n21465) );
  XOR U29610 ( .A(n21471), .B(n21472), .Z(n20905) );
  ANDN U29611 ( .B(n21473), .A(n21474), .Z(n21471) );
  AND U29612 ( .A(a[78]), .B(b[17]), .Z(n21470) );
  XOR U29613 ( .A(n21476), .B(n21477), .Z(n20910) );
  ANDN U29614 ( .B(n21478), .A(n21479), .Z(n21476) );
  AND U29615 ( .A(a[79]), .B(b[16]), .Z(n21475) );
  XOR U29616 ( .A(n21481), .B(n21482), .Z(n20915) );
  ANDN U29617 ( .B(n21483), .A(n21484), .Z(n21481) );
  AND U29618 ( .A(a[80]), .B(b[15]), .Z(n21480) );
  XOR U29619 ( .A(n21486), .B(n21487), .Z(n20920) );
  ANDN U29620 ( .B(n21488), .A(n21489), .Z(n21486) );
  AND U29621 ( .A(a[81]), .B(b[14]), .Z(n21485) );
  XOR U29622 ( .A(n21491), .B(n21492), .Z(n20925) );
  ANDN U29623 ( .B(n21493), .A(n21494), .Z(n21491) );
  AND U29624 ( .A(a[82]), .B(b[13]), .Z(n21490) );
  XOR U29625 ( .A(n21496), .B(n21497), .Z(n20930) );
  ANDN U29626 ( .B(n21498), .A(n21499), .Z(n21496) );
  AND U29627 ( .A(a[83]), .B(b[12]), .Z(n21495) );
  XOR U29628 ( .A(n21501), .B(n21502), .Z(n20935) );
  ANDN U29629 ( .B(n21503), .A(n21504), .Z(n21501) );
  AND U29630 ( .A(a[84]), .B(b[11]), .Z(n21500) );
  XOR U29631 ( .A(n21506), .B(n21507), .Z(n20940) );
  ANDN U29632 ( .B(n21508), .A(n21509), .Z(n21506) );
  AND U29633 ( .A(a[85]), .B(b[10]), .Z(n21505) );
  XOR U29634 ( .A(n21511), .B(n21512), .Z(n20945) );
  ANDN U29635 ( .B(n21513), .A(n21514), .Z(n21511) );
  AND U29636 ( .A(b[9]), .B(a[86]), .Z(n21510) );
  XOR U29637 ( .A(n21516), .B(n21517), .Z(n20950) );
  ANDN U29638 ( .B(n21518), .A(n21519), .Z(n21516) );
  AND U29639 ( .A(b[8]), .B(a[87]), .Z(n21515) );
  XOR U29640 ( .A(n21521), .B(n21522), .Z(n20955) );
  ANDN U29641 ( .B(n21523), .A(n21524), .Z(n21521) );
  AND U29642 ( .A(b[7]), .B(a[88]), .Z(n21520) );
  XOR U29643 ( .A(n21526), .B(n21527), .Z(n20960) );
  ANDN U29644 ( .B(n21528), .A(n21529), .Z(n21526) );
  AND U29645 ( .A(b[6]), .B(a[89]), .Z(n21525) );
  XOR U29646 ( .A(n21531), .B(n21532), .Z(n20965) );
  ANDN U29647 ( .B(n21533), .A(n21534), .Z(n21531) );
  AND U29648 ( .A(b[5]), .B(a[90]), .Z(n21530) );
  XOR U29649 ( .A(n21536), .B(n21537), .Z(n20970) );
  ANDN U29650 ( .B(n21538), .A(n21539), .Z(n21536) );
  AND U29651 ( .A(b[4]), .B(a[91]), .Z(n21535) );
  XOR U29652 ( .A(n21541), .B(n21542), .Z(n20975) );
  ANDN U29653 ( .B(n20987), .A(n20988), .Z(n21541) );
  AND U29654 ( .A(b[2]), .B(a[92]), .Z(n21543) );
  XNOR U29655 ( .A(n21538), .B(n21542), .Z(n21544) );
  XOR U29656 ( .A(n21545), .B(n21546), .Z(n21542) );
  OR U29657 ( .A(n20990), .B(n20991), .Z(n21546) );
  XNOR U29658 ( .A(n21548), .B(n21549), .Z(n21547) );
  XOR U29659 ( .A(n21548), .B(n21551), .Z(n20990) );
  NAND U29660 ( .A(b[1]), .B(a[92]), .Z(n21551) );
  IV U29661 ( .A(n21545), .Z(n21548) );
  NANDN U29662 ( .A(n17), .B(n18), .Z(n21545) );
  XOR U29663 ( .A(n21552), .B(n21553), .Z(n18) );
  NAND U29664 ( .A(a[92]), .B(b[0]), .Z(n17) );
  XNOR U29665 ( .A(n21533), .B(n21537), .Z(n21554) );
  XNOR U29666 ( .A(n21528), .B(n21532), .Z(n21555) );
  XNOR U29667 ( .A(n21523), .B(n21527), .Z(n21556) );
  XNOR U29668 ( .A(n21518), .B(n21522), .Z(n21557) );
  XNOR U29669 ( .A(n21513), .B(n21517), .Z(n21558) );
  XNOR U29670 ( .A(n21508), .B(n21512), .Z(n21559) );
  XNOR U29671 ( .A(n21503), .B(n21507), .Z(n21560) );
  XNOR U29672 ( .A(n21498), .B(n21502), .Z(n21561) );
  XNOR U29673 ( .A(n21493), .B(n21497), .Z(n21562) );
  XNOR U29674 ( .A(n21488), .B(n21492), .Z(n21563) );
  XNOR U29675 ( .A(n21483), .B(n21487), .Z(n21564) );
  XNOR U29676 ( .A(n21478), .B(n21482), .Z(n21565) );
  XNOR U29677 ( .A(n21473), .B(n21477), .Z(n21566) );
  XNOR U29678 ( .A(n21468), .B(n21472), .Z(n21567) );
  XNOR U29679 ( .A(n21463), .B(n21467), .Z(n21568) );
  XNOR U29680 ( .A(n21458), .B(n21462), .Z(n21569) );
  XNOR U29681 ( .A(n21453), .B(n21457), .Z(n21570) );
  XNOR U29682 ( .A(n21448), .B(n21452), .Z(n21571) );
  XNOR U29683 ( .A(n21443), .B(n21447), .Z(n21572) );
  XNOR U29684 ( .A(n21438), .B(n21442), .Z(n21573) );
  XNOR U29685 ( .A(n21433), .B(n21437), .Z(n21574) );
  XNOR U29686 ( .A(n21428), .B(n21432), .Z(n21575) );
  XNOR U29687 ( .A(n21423), .B(n21427), .Z(n21576) );
  XNOR U29688 ( .A(n21418), .B(n21422), .Z(n21577) );
  XNOR U29689 ( .A(n21413), .B(n21417), .Z(n21578) );
  XNOR U29690 ( .A(n21408), .B(n21412), .Z(n21579) );
  XNOR U29691 ( .A(n21403), .B(n21407), .Z(n21580) );
  XNOR U29692 ( .A(n21398), .B(n21402), .Z(n21581) );
  XNOR U29693 ( .A(n21393), .B(n21397), .Z(n21582) );
  XNOR U29694 ( .A(n21388), .B(n21392), .Z(n21583) );
  XNOR U29695 ( .A(n21383), .B(n21387), .Z(n21584) );
  XNOR U29696 ( .A(n21378), .B(n21382), .Z(n21585) );
  XNOR U29697 ( .A(n21373), .B(n21377), .Z(n21586) );
  XNOR U29698 ( .A(n21368), .B(n21372), .Z(n21587) );
  XNOR U29699 ( .A(n21363), .B(n21367), .Z(n21588) );
  XNOR U29700 ( .A(n21358), .B(n21362), .Z(n21589) );
  XNOR U29701 ( .A(n21353), .B(n21357), .Z(n21590) );
  XNOR U29702 ( .A(n21348), .B(n21352), .Z(n21591) );
  XNOR U29703 ( .A(n21343), .B(n21347), .Z(n21592) );
  XNOR U29704 ( .A(n21338), .B(n21342), .Z(n21593) );
  XNOR U29705 ( .A(n21333), .B(n21337), .Z(n21594) );
  XNOR U29706 ( .A(n21328), .B(n21332), .Z(n21595) );
  XNOR U29707 ( .A(n21323), .B(n21327), .Z(n21596) );
  XNOR U29708 ( .A(n21318), .B(n21322), .Z(n21597) );
  XNOR U29709 ( .A(n21313), .B(n21317), .Z(n21598) );
  XNOR U29710 ( .A(n21308), .B(n21312), .Z(n21599) );
  XNOR U29711 ( .A(n21303), .B(n21307), .Z(n21600) );
  XNOR U29712 ( .A(n21298), .B(n21302), .Z(n21601) );
  XNOR U29713 ( .A(n21293), .B(n21297), .Z(n21602) );
  XNOR U29714 ( .A(n21288), .B(n21292), .Z(n21603) );
  XNOR U29715 ( .A(n21283), .B(n21287), .Z(n21604) );
  XNOR U29716 ( .A(n21278), .B(n21282), .Z(n21605) );
  XNOR U29717 ( .A(n21273), .B(n21277), .Z(n21606) );
  XNOR U29718 ( .A(n21268), .B(n21272), .Z(n21607) );
  XNOR U29719 ( .A(n21263), .B(n21267), .Z(n21608) );
  XNOR U29720 ( .A(n21258), .B(n21262), .Z(n21609) );
  XNOR U29721 ( .A(n21253), .B(n21257), .Z(n21610) );
  XNOR U29722 ( .A(n21248), .B(n21252), .Z(n21611) );
  XNOR U29723 ( .A(n21243), .B(n21247), .Z(n21612) );
  XNOR U29724 ( .A(n21238), .B(n21242), .Z(n21613) );
  XNOR U29725 ( .A(n21233), .B(n21237), .Z(n21614) );
  XNOR U29726 ( .A(n21228), .B(n21232), .Z(n21615) );
  XNOR U29727 ( .A(n21223), .B(n21227), .Z(n21616) );
  XNOR U29728 ( .A(n21218), .B(n21222), .Z(n21617) );
  XNOR U29729 ( .A(n21213), .B(n21217), .Z(n21618) );
  XNOR U29730 ( .A(n21208), .B(n21212), .Z(n21619) );
  XNOR U29731 ( .A(n21203), .B(n21207), .Z(n21620) );
  XNOR U29732 ( .A(n21198), .B(n21202), .Z(n21621) );
  XNOR U29733 ( .A(n21193), .B(n21197), .Z(n21622) );
  XNOR U29734 ( .A(n21188), .B(n21192), .Z(n21623) );
  XNOR U29735 ( .A(n21183), .B(n21187), .Z(n21624) );
  XNOR U29736 ( .A(n21178), .B(n21182), .Z(n21625) );
  XNOR U29737 ( .A(n21173), .B(n21177), .Z(n21626) );
  XNOR U29738 ( .A(n21168), .B(n21172), .Z(n21627) );
  XNOR U29739 ( .A(n21163), .B(n21167), .Z(n21628) );
  XNOR U29740 ( .A(n21158), .B(n21162), .Z(n21629) );
  XNOR U29741 ( .A(n21153), .B(n21157), .Z(n21630) );
  XNOR U29742 ( .A(n21148), .B(n21152), .Z(n21631) );
  XNOR U29743 ( .A(n21143), .B(n21147), .Z(n21632) );
  XNOR U29744 ( .A(n21138), .B(n21142), .Z(n21633) );
  XNOR U29745 ( .A(n21133), .B(n21137), .Z(n21634) );
  XNOR U29746 ( .A(n21128), .B(n21132), .Z(n21635) );
  XNOR U29747 ( .A(n21123), .B(n21127), .Z(n21636) );
  XNOR U29748 ( .A(n21118), .B(n21122), .Z(n21637) );
  XNOR U29749 ( .A(n21113), .B(n21117), .Z(n21638) );
  XNOR U29750 ( .A(n21108), .B(n21112), .Z(n21639) );
  XNOR U29751 ( .A(n21103), .B(n21107), .Z(n21640) );
  XNOR U29752 ( .A(n21098), .B(n21102), .Z(n21641) );
  XNOR U29753 ( .A(n21093), .B(n21097), .Z(n21642) );
  XNOR U29754 ( .A(n21088), .B(n21092), .Z(n21643) );
  XOR U29755 ( .A(n21644), .B(n21087), .Z(n21088) );
  AND U29756 ( .A(a[0]), .B(b[94]), .Z(n21644) );
  XNOR U29757 ( .A(n21645), .B(n21087), .Z(n21089) );
  XNOR U29758 ( .A(n21646), .B(n21647), .Z(n21087) );
  ANDN U29759 ( .B(n21648), .A(n21649), .Z(n21646) );
  AND U29760 ( .A(a[1]), .B(b[93]), .Z(n21645) );
  XOR U29761 ( .A(n21651), .B(n21652), .Z(n21092) );
  ANDN U29762 ( .B(n21653), .A(n21654), .Z(n21651) );
  AND U29763 ( .A(a[2]), .B(b[92]), .Z(n21650) );
  XOR U29764 ( .A(n21656), .B(n21657), .Z(n21097) );
  ANDN U29765 ( .B(n21658), .A(n21659), .Z(n21656) );
  AND U29766 ( .A(a[3]), .B(b[91]), .Z(n21655) );
  XOR U29767 ( .A(n21661), .B(n21662), .Z(n21102) );
  ANDN U29768 ( .B(n21663), .A(n21664), .Z(n21661) );
  AND U29769 ( .A(a[4]), .B(b[90]), .Z(n21660) );
  XOR U29770 ( .A(n21666), .B(n21667), .Z(n21107) );
  ANDN U29771 ( .B(n21668), .A(n21669), .Z(n21666) );
  AND U29772 ( .A(a[5]), .B(b[89]), .Z(n21665) );
  XOR U29773 ( .A(n21671), .B(n21672), .Z(n21112) );
  ANDN U29774 ( .B(n21673), .A(n21674), .Z(n21671) );
  AND U29775 ( .A(a[6]), .B(b[88]), .Z(n21670) );
  XOR U29776 ( .A(n21676), .B(n21677), .Z(n21117) );
  ANDN U29777 ( .B(n21678), .A(n21679), .Z(n21676) );
  AND U29778 ( .A(a[7]), .B(b[87]), .Z(n21675) );
  XOR U29779 ( .A(n21681), .B(n21682), .Z(n21122) );
  ANDN U29780 ( .B(n21683), .A(n21684), .Z(n21681) );
  AND U29781 ( .A(a[8]), .B(b[86]), .Z(n21680) );
  XOR U29782 ( .A(n21686), .B(n21687), .Z(n21127) );
  ANDN U29783 ( .B(n21688), .A(n21689), .Z(n21686) );
  AND U29784 ( .A(a[9]), .B(b[85]), .Z(n21685) );
  XOR U29785 ( .A(n21691), .B(n21692), .Z(n21132) );
  ANDN U29786 ( .B(n21693), .A(n21694), .Z(n21691) );
  AND U29787 ( .A(a[10]), .B(b[84]), .Z(n21690) );
  XOR U29788 ( .A(n21696), .B(n21697), .Z(n21137) );
  ANDN U29789 ( .B(n21698), .A(n21699), .Z(n21696) );
  AND U29790 ( .A(a[11]), .B(b[83]), .Z(n21695) );
  XOR U29791 ( .A(n21701), .B(n21702), .Z(n21142) );
  ANDN U29792 ( .B(n21703), .A(n21704), .Z(n21701) );
  AND U29793 ( .A(a[12]), .B(b[82]), .Z(n21700) );
  XOR U29794 ( .A(n21706), .B(n21707), .Z(n21147) );
  ANDN U29795 ( .B(n21708), .A(n21709), .Z(n21706) );
  AND U29796 ( .A(a[13]), .B(b[81]), .Z(n21705) );
  XOR U29797 ( .A(n21711), .B(n21712), .Z(n21152) );
  ANDN U29798 ( .B(n21713), .A(n21714), .Z(n21711) );
  AND U29799 ( .A(a[14]), .B(b[80]), .Z(n21710) );
  XOR U29800 ( .A(n21716), .B(n21717), .Z(n21157) );
  ANDN U29801 ( .B(n21718), .A(n21719), .Z(n21716) );
  AND U29802 ( .A(a[15]), .B(b[79]), .Z(n21715) );
  XOR U29803 ( .A(n21721), .B(n21722), .Z(n21162) );
  ANDN U29804 ( .B(n21723), .A(n21724), .Z(n21721) );
  AND U29805 ( .A(a[16]), .B(b[78]), .Z(n21720) );
  XOR U29806 ( .A(n21726), .B(n21727), .Z(n21167) );
  ANDN U29807 ( .B(n21728), .A(n21729), .Z(n21726) );
  AND U29808 ( .A(a[17]), .B(b[77]), .Z(n21725) );
  XOR U29809 ( .A(n21731), .B(n21732), .Z(n21172) );
  ANDN U29810 ( .B(n21733), .A(n21734), .Z(n21731) );
  AND U29811 ( .A(a[18]), .B(b[76]), .Z(n21730) );
  XOR U29812 ( .A(n21736), .B(n21737), .Z(n21177) );
  ANDN U29813 ( .B(n21738), .A(n21739), .Z(n21736) );
  AND U29814 ( .A(a[19]), .B(b[75]), .Z(n21735) );
  XOR U29815 ( .A(n21741), .B(n21742), .Z(n21182) );
  ANDN U29816 ( .B(n21743), .A(n21744), .Z(n21741) );
  AND U29817 ( .A(a[20]), .B(b[74]), .Z(n21740) );
  XOR U29818 ( .A(n21746), .B(n21747), .Z(n21187) );
  ANDN U29819 ( .B(n21748), .A(n21749), .Z(n21746) );
  AND U29820 ( .A(a[21]), .B(b[73]), .Z(n21745) );
  XOR U29821 ( .A(n21751), .B(n21752), .Z(n21192) );
  ANDN U29822 ( .B(n21753), .A(n21754), .Z(n21751) );
  AND U29823 ( .A(a[22]), .B(b[72]), .Z(n21750) );
  XOR U29824 ( .A(n21756), .B(n21757), .Z(n21197) );
  ANDN U29825 ( .B(n21758), .A(n21759), .Z(n21756) );
  AND U29826 ( .A(a[23]), .B(b[71]), .Z(n21755) );
  XOR U29827 ( .A(n21761), .B(n21762), .Z(n21202) );
  ANDN U29828 ( .B(n21763), .A(n21764), .Z(n21761) );
  AND U29829 ( .A(a[24]), .B(b[70]), .Z(n21760) );
  XOR U29830 ( .A(n21766), .B(n21767), .Z(n21207) );
  ANDN U29831 ( .B(n21768), .A(n21769), .Z(n21766) );
  AND U29832 ( .A(a[25]), .B(b[69]), .Z(n21765) );
  XOR U29833 ( .A(n21771), .B(n21772), .Z(n21212) );
  ANDN U29834 ( .B(n21773), .A(n21774), .Z(n21771) );
  AND U29835 ( .A(a[26]), .B(b[68]), .Z(n21770) );
  XOR U29836 ( .A(n21776), .B(n21777), .Z(n21217) );
  ANDN U29837 ( .B(n21778), .A(n21779), .Z(n21776) );
  AND U29838 ( .A(a[27]), .B(b[67]), .Z(n21775) );
  XOR U29839 ( .A(n21781), .B(n21782), .Z(n21222) );
  ANDN U29840 ( .B(n21783), .A(n21784), .Z(n21781) );
  AND U29841 ( .A(a[28]), .B(b[66]), .Z(n21780) );
  XOR U29842 ( .A(n21786), .B(n21787), .Z(n21227) );
  ANDN U29843 ( .B(n21788), .A(n21789), .Z(n21786) );
  AND U29844 ( .A(a[29]), .B(b[65]), .Z(n21785) );
  XOR U29845 ( .A(n21791), .B(n21792), .Z(n21232) );
  ANDN U29846 ( .B(n21793), .A(n21794), .Z(n21791) );
  AND U29847 ( .A(a[30]), .B(b[64]), .Z(n21790) );
  XOR U29848 ( .A(n21796), .B(n21797), .Z(n21237) );
  ANDN U29849 ( .B(n21798), .A(n21799), .Z(n21796) );
  AND U29850 ( .A(a[31]), .B(b[63]), .Z(n21795) );
  XOR U29851 ( .A(n21801), .B(n21802), .Z(n21242) );
  ANDN U29852 ( .B(n21803), .A(n21804), .Z(n21801) );
  AND U29853 ( .A(a[32]), .B(b[62]), .Z(n21800) );
  XOR U29854 ( .A(n21806), .B(n21807), .Z(n21247) );
  ANDN U29855 ( .B(n21808), .A(n21809), .Z(n21806) );
  AND U29856 ( .A(a[33]), .B(b[61]), .Z(n21805) );
  XOR U29857 ( .A(n21811), .B(n21812), .Z(n21252) );
  ANDN U29858 ( .B(n21813), .A(n21814), .Z(n21811) );
  AND U29859 ( .A(a[34]), .B(b[60]), .Z(n21810) );
  XOR U29860 ( .A(n21816), .B(n21817), .Z(n21257) );
  ANDN U29861 ( .B(n21818), .A(n21819), .Z(n21816) );
  AND U29862 ( .A(a[35]), .B(b[59]), .Z(n21815) );
  XOR U29863 ( .A(n21821), .B(n21822), .Z(n21262) );
  ANDN U29864 ( .B(n21823), .A(n21824), .Z(n21821) );
  AND U29865 ( .A(a[36]), .B(b[58]), .Z(n21820) );
  XOR U29866 ( .A(n21826), .B(n21827), .Z(n21267) );
  ANDN U29867 ( .B(n21828), .A(n21829), .Z(n21826) );
  AND U29868 ( .A(a[37]), .B(b[57]), .Z(n21825) );
  XOR U29869 ( .A(n21831), .B(n21832), .Z(n21272) );
  ANDN U29870 ( .B(n21833), .A(n21834), .Z(n21831) );
  AND U29871 ( .A(a[38]), .B(b[56]), .Z(n21830) );
  XOR U29872 ( .A(n21836), .B(n21837), .Z(n21277) );
  ANDN U29873 ( .B(n21838), .A(n21839), .Z(n21836) );
  AND U29874 ( .A(a[39]), .B(b[55]), .Z(n21835) );
  XOR U29875 ( .A(n21841), .B(n21842), .Z(n21282) );
  ANDN U29876 ( .B(n21843), .A(n21844), .Z(n21841) );
  AND U29877 ( .A(a[40]), .B(b[54]), .Z(n21840) );
  XOR U29878 ( .A(n21846), .B(n21847), .Z(n21287) );
  ANDN U29879 ( .B(n21848), .A(n21849), .Z(n21846) );
  AND U29880 ( .A(a[41]), .B(b[53]), .Z(n21845) );
  XOR U29881 ( .A(n21851), .B(n21852), .Z(n21292) );
  ANDN U29882 ( .B(n21853), .A(n21854), .Z(n21851) );
  AND U29883 ( .A(a[42]), .B(b[52]), .Z(n21850) );
  XOR U29884 ( .A(n21856), .B(n21857), .Z(n21297) );
  ANDN U29885 ( .B(n21858), .A(n21859), .Z(n21856) );
  AND U29886 ( .A(a[43]), .B(b[51]), .Z(n21855) );
  XOR U29887 ( .A(n21861), .B(n21862), .Z(n21302) );
  ANDN U29888 ( .B(n21863), .A(n21864), .Z(n21861) );
  AND U29889 ( .A(a[44]), .B(b[50]), .Z(n21860) );
  XOR U29890 ( .A(n21866), .B(n21867), .Z(n21307) );
  ANDN U29891 ( .B(n21868), .A(n21869), .Z(n21866) );
  AND U29892 ( .A(a[45]), .B(b[49]), .Z(n21865) );
  XOR U29893 ( .A(n21871), .B(n21872), .Z(n21312) );
  ANDN U29894 ( .B(n21873), .A(n21874), .Z(n21871) );
  AND U29895 ( .A(a[46]), .B(b[48]), .Z(n21870) );
  XOR U29896 ( .A(n21876), .B(n21877), .Z(n21317) );
  ANDN U29897 ( .B(n21878), .A(n21879), .Z(n21876) );
  AND U29898 ( .A(a[47]), .B(b[47]), .Z(n21875) );
  XOR U29899 ( .A(n21881), .B(n21882), .Z(n21322) );
  ANDN U29900 ( .B(n21883), .A(n21884), .Z(n21881) );
  AND U29901 ( .A(a[48]), .B(b[46]), .Z(n21880) );
  XOR U29902 ( .A(n21886), .B(n21887), .Z(n21327) );
  ANDN U29903 ( .B(n21888), .A(n21889), .Z(n21886) );
  AND U29904 ( .A(a[49]), .B(b[45]), .Z(n21885) );
  XOR U29905 ( .A(n21891), .B(n21892), .Z(n21332) );
  ANDN U29906 ( .B(n21893), .A(n21894), .Z(n21891) );
  AND U29907 ( .A(a[50]), .B(b[44]), .Z(n21890) );
  XOR U29908 ( .A(n21896), .B(n21897), .Z(n21337) );
  ANDN U29909 ( .B(n21898), .A(n21899), .Z(n21896) );
  AND U29910 ( .A(a[51]), .B(b[43]), .Z(n21895) );
  XOR U29911 ( .A(n21901), .B(n21902), .Z(n21342) );
  ANDN U29912 ( .B(n21903), .A(n21904), .Z(n21901) );
  AND U29913 ( .A(a[52]), .B(b[42]), .Z(n21900) );
  XOR U29914 ( .A(n21906), .B(n21907), .Z(n21347) );
  ANDN U29915 ( .B(n21908), .A(n21909), .Z(n21906) );
  AND U29916 ( .A(a[53]), .B(b[41]), .Z(n21905) );
  XOR U29917 ( .A(n21911), .B(n21912), .Z(n21352) );
  ANDN U29918 ( .B(n21913), .A(n21914), .Z(n21911) );
  AND U29919 ( .A(a[54]), .B(b[40]), .Z(n21910) );
  XOR U29920 ( .A(n21916), .B(n21917), .Z(n21357) );
  ANDN U29921 ( .B(n21918), .A(n21919), .Z(n21916) );
  AND U29922 ( .A(a[55]), .B(b[39]), .Z(n21915) );
  XOR U29923 ( .A(n21921), .B(n21922), .Z(n21362) );
  ANDN U29924 ( .B(n21923), .A(n21924), .Z(n21921) );
  AND U29925 ( .A(a[56]), .B(b[38]), .Z(n21920) );
  XOR U29926 ( .A(n21926), .B(n21927), .Z(n21367) );
  ANDN U29927 ( .B(n21928), .A(n21929), .Z(n21926) );
  AND U29928 ( .A(a[57]), .B(b[37]), .Z(n21925) );
  XOR U29929 ( .A(n21931), .B(n21932), .Z(n21372) );
  ANDN U29930 ( .B(n21933), .A(n21934), .Z(n21931) );
  AND U29931 ( .A(a[58]), .B(b[36]), .Z(n21930) );
  XOR U29932 ( .A(n21936), .B(n21937), .Z(n21377) );
  ANDN U29933 ( .B(n21938), .A(n21939), .Z(n21936) );
  AND U29934 ( .A(a[59]), .B(b[35]), .Z(n21935) );
  XOR U29935 ( .A(n21941), .B(n21942), .Z(n21382) );
  ANDN U29936 ( .B(n21943), .A(n21944), .Z(n21941) );
  AND U29937 ( .A(a[60]), .B(b[34]), .Z(n21940) );
  XOR U29938 ( .A(n21946), .B(n21947), .Z(n21387) );
  ANDN U29939 ( .B(n21948), .A(n21949), .Z(n21946) );
  AND U29940 ( .A(a[61]), .B(b[33]), .Z(n21945) );
  XOR U29941 ( .A(n21951), .B(n21952), .Z(n21392) );
  ANDN U29942 ( .B(n21953), .A(n21954), .Z(n21951) );
  AND U29943 ( .A(a[62]), .B(b[32]), .Z(n21950) );
  XOR U29944 ( .A(n21956), .B(n21957), .Z(n21397) );
  ANDN U29945 ( .B(n21958), .A(n21959), .Z(n21956) );
  AND U29946 ( .A(a[63]), .B(b[31]), .Z(n21955) );
  XOR U29947 ( .A(n21961), .B(n21962), .Z(n21402) );
  ANDN U29948 ( .B(n21963), .A(n21964), .Z(n21961) );
  AND U29949 ( .A(a[64]), .B(b[30]), .Z(n21960) );
  XOR U29950 ( .A(n21966), .B(n21967), .Z(n21407) );
  ANDN U29951 ( .B(n21968), .A(n21969), .Z(n21966) );
  AND U29952 ( .A(a[65]), .B(b[29]), .Z(n21965) );
  XOR U29953 ( .A(n21971), .B(n21972), .Z(n21412) );
  ANDN U29954 ( .B(n21973), .A(n21974), .Z(n21971) );
  AND U29955 ( .A(a[66]), .B(b[28]), .Z(n21970) );
  XOR U29956 ( .A(n21976), .B(n21977), .Z(n21417) );
  ANDN U29957 ( .B(n21978), .A(n21979), .Z(n21976) );
  AND U29958 ( .A(a[67]), .B(b[27]), .Z(n21975) );
  XOR U29959 ( .A(n21981), .B(n21982), .Z(n21422) );
  ANDN U29960 ( .B(n21983), .A(n21984), .Z(n21981) );
  AND U29961 ( .A(a[68]), .B(b[26]), .Z(n21980) );
  XOR U29962 ( .A(n21986), .B(n21987), .Z(n21427) );
  ANDN U29963 ( .B(n21988), .A(n21989), .Z(n21986) );
  AND U29964 ( .A(a[69]), .B(b[25]), .Z(n21985) );
  XOR U29965 ( .A(n21991), .B(n21992), .Z(n21432) );
  ANDN U29966 ( .B(n21993), .A(n21994), .Z(n21991) );
  AND U29967 ( .A(a[70]), .B(b[24]), .Z(n21990) );
  XOR U29968 ( .A(n21996), .B(n21997), .Z(n21437) );
  ANDN U29969 ( .B(n21998), .A(n21999), .Z(n21996) );
  AND U29970 ( .A(a[71]), .B(b[23]), .Z(n21995) );
  XOR U29971 ( .A(n22001), .B(n22002), .Z(n21442) );
  ANDN U29972 ( .B(n22003), .A(n22004), .Z(n22001) );
  AND U29973 ( .A(a[72]), .B(b[22]), .Z(n22000) );
  XOR U29974 ( .A(n22006), .B(n22007), .Z(n21447) );
  ANDN U29975 ( .B(n22008), .A(n22009), .Z(n22006) );
  AND U29976 ( .A(a[73]), .B(b[21]), .Z(n22005) );
  XOR U29977 ( .A(n22011), .B(n22012), .Z(n21452) );
  ANDN U29978 ( .B(n22013), .A(n22014), .Z(n22011) );
  AND U29979 ( .A(a[74]), .B(b[20]), .Z(n22010) );
  XOR U29980 ( .A(n22016), .B(n22017), .Z(n21457) );
  ANDN U29981 ( .B(n22018), .A(n22019), .Z(n22016) );
  AND U29982 ( .A(a[75]), .B(b[19]), .Z(n22015) );
  XOR U29983 ( .A(n22021), .B(n22022), .Z(n21462) );
  ANDN U29984 ( .B(n22023), .A(n22024), .Z(n22021) );
  AND U29985 ( .A(a[76]), .B(b[18]), .Z(n22020) );
  XOR U29986 ( .A(n22026), .B(n22027), .Z(n21467) );
  ANDN U29987 ( .B(n22028), .A(n22029), .Z(n22026) );
  AND U29988 ( .A(a[77]), .B(b[17]), .Z(n22025) );
  XOR U29989 ( .A(n22031), .B(n22032), .Z(n21472) );
  ANDN U29990 ( .B(n22033), .A(n22034), .Z(n22031) );
  AND U29991 ( .A(a[78]), .B(b[16]), .Z(n22030) );
  XOR U29992 ( .A(n22036), .B(n22037), .Z(n21477) );
  ANDN U29993 ( .B(n22038), .A(n22039), .Z(n22036) );
  AND U29994 ( .A(a[79]), .B(b[15]), .Z(n22035) );
  XOR U29995 ( .A(n22041), .B(n22042), .Z(n21482) );
  ANDN U29996 ( .B(n22043), .A(n22044), .Z(n22041) );
  AND U29997 ( .A(a[80]), .B(b[14]), .Z(n22040) );
  XOR U29998 ( .A(n22046), .B(n22047), .Z(n21487) );
  ANDN U29999 ( .B(n22048), .A(n22049), .Z(n22046) );
  AND U30000 ( .A(a[81]), .B(b[13]), .Z(n22045) );
  XOR U30001 ( .A(n22051), .B(n22052), .Z(n21492) );
  ANDN U30002 ( .B(n22053), .A(n22054), .Z(n22051) );
  AND U30003 ( .A(a[82]), .B(b[12]), .Z(n22050) );
  XOR U30004 ( .A(n22056), .B(n22057), .Z(n21497) );
  ANDN U30005 ( .B(n22058), .A(n22059), .Z(n22056) );
  AND U30006 ( .A(a[83]), .B(b[11]), .Z(n22055) );
  XOR U30007 ( .A(n22061), .B(n22062), .Z(n21502) );
  ANDN U30008 ( .B(n22063), .A(n22064), .Z(n22061) );
  AND U30009 ( .A(a[84]), .B(b[10]), .Z(n22060) );
  XOR U30010 ( .A(n22066), .B(n22067), .Z(n21507) );
  ANDN U30011 ( .B(n22068), .A(n22069), .Z(n22066) );
  AND U30012 ( .A(b[9]), .B(a[85]), .Z(n22065) );
  XOR U30013 ( .A(n22071), .B(n22072), .Z(n21512) );
  ANDN U30014 ( .B(n22073), .A(n22074), .Z(n22071) );
  AND U30015 ( .A(b[8]), .B(a[86]), .Z(n22070) );
  XOR U30016 ( .A(n22076), .B(n22077), .Z(n21517) );
  ANDN U30017 ( .B(n22078), .A(n22079), .Z(n22076) );
  AND U30018 ( .A(b[7]), .B(a[87]), .Z(n22075) );
  XOR U30019 ( .A(n22081), .B(n22082), .Z(n21522) );
  ANDN U30020 ( .B(n22083), .A(n22084), .Z(n22081) );
  AND U30021 ( .A(b[6]), .B(a[88]), .Z(n22080) );
  XOR U30022 ( .A(n22086), .B(n22087), .Z(n21527) );
  ANDN U30023 ( .B(n22088), .A(n22089), .Z(n22086) );
  AND U30024 ( .A(b[5]), .B(a[89]), .Z(n22085) );
  XOR U30025 ( .A(n22091), .B(n22092), .Z(n21532) );
  ANDN U30026 ( .B(n22093), .A(n22094), .Z(n22091) );
  AND U30027 ( .A(b[4]), .B(a[90]), .Z(n22090) );
  XOR U30028 ( .A(n22096), .B(n22097), .Z(n21537) );
  ANDN U30029 ( .B(n21549), .A(n21550), .Z(n22096) );
  AND U30030 ( .A(b[2]), .B(a[91]), .Z(n22098) );
  XNOR U30031 ( .A(n22093), .B(n22097), .Z(n22099) );
  XOR U30032 ( .A(n22100), .B(n22101), .Z(n22097) );
  OR U30033 ( .A(n21552), .B(n21553), .Z(n22101) );
  XNOR U30034 ( .A(n22103), .B(n22104), .Z(n22102) );
  XOR U30035 ( .A(n22103), .B(n22106), .Z(n21552) );
  NAND U30036 ( .A(b[1]), .B(a[91]), .Z(n22106) );
  IV U30037 ( .A(n22100), .Z(n22103) );
  NANDN U30038 ( .A(n19), .B(n20), .Z(n22100) );
  XOR U30039 ( .A(n22107), .B(n22108), .Z(n20) );
  NAND U30040 ( .A(a[91]), .B(b[0]), .Z(n19) );
  XNOR U30041 ( .A(n22088), .B(n22092), .Z(n22109) );
  XNOR U30042 ( .A(n22083), .B(n22087), .Z(n22110) );
  XNOR U30043 ( .A(n22078), .B(n22082), .Z(n22111) );
  XNOR U30044 ( .A(n22073), .B(n22077), .Z(n22112) );
  XNOR U30045 ( .A(n22068), .B(n22072), .Z(n22113) );
  XNOR U30046 ( .A(n22063), .B(n22067), .Z(n22114) );
  XNOR U30047 ( .A(n22058), .B(n22062), .Z(n22115) );
  XNOR U30048 ( .A(n22053), .B(n22057), .Z(n22116) );
  XNOR U30049 ( .A(n22048), .B(n22052), .Z(n22117) );
  XNOR U30050 ( .A(n22043), .B(n22047), .Z(n22118) );
  XNOR U30051 ( .A(n22038), .B(n22042), .Z(n22119) );
  XNOR U30052 ( .A(n22033), .B(n22037), .Z(n22120) );
  XNOR U30053 ( .A(n22028), .B(n22032), .Z(n22121) );
  XNOR U30054 ( .A(n22023), .B(n22027), .Z(n22122) );
  XNOR U30055 ( .A(n22018), .B(n22022), .Z(n22123) );
  XNOR U30056 ( .A(n22013), .B(n22017), .Z(n22124) );
  XNOR U30057 ( .A(n22008), .B(n22012), .Z(n22125) );
  XNOR U30058 ( .A(n22003), .B(n22007), .Z(n22126) );
  XNOR U30059 ( .A(n21998), .B(n22002), .Z(n22127) );
  XNOR U30060 ( .A(n21993), .B(n21997), .Z(n22128) );
  XNOR U30061 ( .A(n21988), .B(n21992), .Z(n22129) );
  XNOR U30062 ( .A(n21983), .B(n21987), .Z(n22130) );
  XNOR U30063 ( .A(n21978), .B(n21982), .Z(n22131) );
  XNOR U30064 ( .A(n21973), .B(n21977), .Z(n22132) );
  XNOR U30065 ( .A(n21968), .B(n21972), .Z(n22133) );
  XNOR U30066 ( .A(n21963), .B(n21967), .Z(n22134) );
  XNOR U30067 ( .A(n21958), .B(n21962), .Z(n22135) );
  XNOR U30068 ( .A(n21953), .B(n21957), .Z(n22136) );
  XNOR U30069 ( .A(n21948), .B(n21952), .Z(n22137) );
  XNOR U30070 ( .A(n21943), .B(n21947), .Z(n22138) );
  XNOR U30071 ( .A(n21938), .B(n21942), .Z(n22139) );
  XNOR U30072 ( .A(n21933), .B(n21937), .Z(n22140) );
  XNOR U30073 ( .A(n21928), .B(n21932), .Z(n22141) );
  XNOR U30074 ( .A(n21923), .B(n21927), .Z(n22142) );
  XNOR U30075 ( .A(n21918), .B(n21922), .Z(n22143) );
  XNOR U30076 ( .A(n21913), .B(n21917), .Z(n22144) );
  XNOR U30077 ( .A(n21908), .B(n21912), .Z(n22145) );
  XNOR U30078 ( .A(n21903), .B(n21907), .Z(n22146) );
  XNOR U30079 ( .A(n21898), .B(n21902), .Z(n22147) );
  XNOR U30080 ( .A(n21893), .B(n21897), .Z(n22148) );
  XNOR U30081 ( .A(n21888), .B(n21892), .Z(n22149) );
  XNOR U30082 ( .A(n21883), .B(n21887), .Z(n22150) );
  XNOR U30083 ( .A(n21878), .B(n21882), .Z(n22151) );
  XNOR U30084 ( .A(n21873), .B(n21877), .Z(n22152) );
  XNOR U30085 ( .A(n21868), .B(n21872), .Z(n22153) );
  XNOR U30086 ( .A(n21863), .B(n21867), .Z(n22154) );
  XNOR U30087 ( .A(n21858), .B(n21862), .Z(n22155) );
  XNOR U30088 ( .A(n21853), .B(n21857), .Z(n22156) );
  XNOR U30089 ( .A(n21848), .B(n21852), .Z(n22157) );
  XNOR U30090 ( .A(n21843), .B(n21847), .Z(n22158) );
  XNOR U30091 ( .A(n21838), .B(n21842), .Z(n22159) );
  XNOR U30092 ( .A(n21833), .B(n21837), .Z(n22160) );
  XNOR U30093 ( .A(n21828), .B(n21832), .Z(n22161) );
  XNOR U30094 ( .A(n21823), .B(n21827), .Z(n22162) );
  XNOR U30095 ( .A(n21818), .B(n21822), .Z(n22163) );
  XNOR U30096 ( .A(n21813), .B(n21817), .Z(n22164) );
  XNOR U30097 ( .A(n21808), .B(n21812), .Z(n22165) );
  XNOR U30098 ( .A(n21803), .B(n21807), .Z(n22166) );
  XNOR U30099 ( .A(n21798), .B(n21802), .Z(n22167) );
  XNOR U30100 ( .A(n21793), .B(n21797), .Z(n22168) );
  XNOR U30101 ( .A(n21788), .B(n21792), .Z(n22169) );
  XNOR U30102 ( .A(n21783), .B(n21787), .Z(n22170) );
  XNOR U30103 ( .A(n21778), .B(n21782), .Z(n22171) );
  XNOR U30104 ( .A(n21773), .B(n21777), .Z(n22172) );
  XNOR U30105 ( .A(n21768), .B(n21772), .Z(n22173) );
  XNOR U30106 ( .A(n21763), .B(n21767), .Z(n22174) );
  XNOR U30107 ( .A(n21758), .B(n21762), .Z(n22175) );
  XNOR U30108 ( .A(n21753), .B(n21757), .Z(n22176) );
  XNOR U30109 ( .A(n21748), .B(n21752), .Z(n22177) );
  XNOR U30110 ( .A(n21743), .B(n21747), .Z(n22178) );
  XNOR U30111 ( .A(n21738), .B(n21742), .Z(n22179) );
  XNOR U30112 ( .A(n21733), .B(n21737), .Z(n22180) );
  XNOR U30113 ( .A(n21728), .B(n21732), .Z(n22181) );
  XNOR U30114 ( .A(n21723), .B(n21727), .Z(n22182) );
  XNOR U30115 ( .A(n21718), .B(n21722), .Z(n22183) );
  XNOR U30116 ( .A(n21713), .B(n21717), .Z(n22184) );
  XNOR U30117 ( .A(n21708), .B(n21712), .Z(n22185) );
  XNOR U30118 ( .A(n21703), .B(n21707), .Z(n22186) );
  XNOR U30119 ( .A(n21698), .B(n21702), .Z(n22187) );
  XNOR U30120 ( .A(n21693), .B(n21697), .Z(n22188) );
  XNOR U30121 ( .A(n21688), .B(n21692), .Z(n22189) );
  XNOR U30122 ( .A(n21683), .B(n21687), .Z(n22190) );
  XNOR U30123 ( .A(n21678), .B(n21682), .Z(n22191) );
  XNOR U30124 ( .A(n21673), .B(n21677), .Z(n22192) );
  XNOR U30125 ( .A(n21668), .B(n21672), .Z(n22193) );
  XNOR U30126 ( .A(n21663), .B(n21667), .Z(n22194) );
  XNOR U30127 ( .A(n21658), .B(n21662), .Z(n22195) );
  XNOR U30128 ( .A(n21653), .B(n21657), .Z(n22196) );
  XNOR U30129 ( .A(n21648), .B(n21652), .Z(n22197) );
  XNOR U30130 ( .A(n22198), .B(n21647), .Z(n21648) );
  AND U30131 ( .A(a[0]), .B(b[93]), .Z(n22198) );
  XOR U30132 ( .A(n22199), .B(n21647), .Z(n21649) );
  XNOR U30133 ( .A(n22200), .B(n22201), .Z(n21647) );
  ANDN U30134 ( .B(n22202), .A(n22203), .Z(n22200) );
  AND U30135 ( .A(a[1]), .B(b[92]), .Z(n22199) );
  XOR U30136 ( .A(n22205), .B(n22206), .Z(n21652) );
  ANDN U30137 ( .B(n22207), .A(n22208), .Z(n22205) );
  AND U30138 ( .A(a[2]), .B(b[91]), .Z(n22204) );
  XOR U30139 ( .A(n22210), .B(n22211), .Z(n21657) );
  ANDN U30140 ( .B(n22212), .A(n22213), .Z(n22210) );
  AND U30141 ( .A(a[3]), .B(b[90]), .Z(n22209) );
  XOR U30142 ( .A(n22215), .B(n22216), .Z(n21662) );
  ANDN U30143 ( .B(n22217), .A(n22218), .Z(n22215) );
  AND U30144 ( .A(a[4]), .B(b[89]), .Z(n22214) );
  XOR U30145 ( .A(n22220), .B(n22221), .Z(n21667) );
  ANDN U30146 ( .B(n22222), .A(n22223), .Z(n22220) );
  AND U30147 ( .A(a[5]), .B(b[88]), .Z(n22219) );
  XOR U30148 ( .A(n22225), .B(n22226), .Z(n21672) );
  ANDN U30149 ( .B(n22227), .A(n22228), .Z(n22225) );
  AND U30150 ( .A(a[6]), .B(b[87]), .Z(n22224) );
  XOR U30151 ( .A(n22230), .B(n22231), .Z(n21677) );
  ANDN U30152 ( .B(n22232), .A(n22233), .Z(n22230) );
  AND U30153 ( .A(a[7]), .B(b[86]), .Z(n22229) );
  XOR U30154 ( .A(n22235), .B(n22236), .Z(n21682) );
  ANDN U30155 ( .B(n22237), .A(n22238), .Z(n22235) );
  AND U30156 ( .A(a[8]), .B(b[85]), .Z(n22234) );
  XOR U30157 ( .A(n22240), .B(n22241), .Z(n21687) );
  ANDN U30158 ( .B(n22242), .A(n22243), .Z(n22240) );
  AND U30159 ( .A(a[9]), .B(b[84]), .Z(n22239) );
  XOR U30160 ( .A(n22245), .B(n22246), .Z(n21692) );
  ANDN U30161 ( .B(n22247), .A(n22248), .Z(n22245) );
  AND U30162 ( .A(a[10]), .B(b[83]), .Z(n22244) );
  XOR U30163 ( .A(n22250), .B(n22251), .Z(n21697) );
  ANDN U30164 ( .B(n22252), .A(n22253), .Z(n22250) );
  AND U30165 ( .A(a[11]), .B(b[82]), .Z(n22249) );
  XOR U30166 ( .A(n22255), .B(n22256), .Z(n21702) );
  ANDN U30167 ( .B(n22257), .A(n22258), .Z(n22255) );
  AND U30168 ( .A(a[12]), .B(b[81]), .Z(n22254) );
  XOR U30169 ( .A(n22260), .B(n22261), .Z(n21707) );
  ANDN U30170 ( .B(n22262), .A(n22263), .Z(n22260) );
  AND U30171 ( .A(a[13]), .B(b[80]), .Z(n22259) );
  XOR U30172 ( .A(n22265), .B(n22266), .Z(n21712) );
  ANDN U30173 ( .B(n22267), .A(n22268), .Z(n22265) );
  AND U30174 ( .A(a[14]), .B(b[79]), .Z(n22264) );
  XOR U30175 ( .A(n22270), .B(n22271), .Z(n21717) );
  ANDN U30176 ( .B(n22272), .A(n22273), .Z(n22270) );
  AND U30177 ( .A(a[15]), .B(b[78]), .Z(n22269) );
  XOR U30178 ( .A(n22275), .B(n22276), .Z(n21722) );
  ANDN U30179 ( .B(n22277), .A(n22278), .Z(n22275) );
  AND U30180 ( .A(a[16]), .B(b[77]), .Z(n22274) );
  XOR U30181 ( .A(n22280), .B(n22281), .Z(n21727) );
  ANDN U30182 ( .B(n22282), .A(n22283), .Z(n22280) );
  AND U30183 ( .A(a[17]), .B(b[76]), .Z(n22279) );
  XOR U30184 ( .A(n22285), .B(n22286), .Z(n21732) );
  ANDN U30185 ( .B(n22287), .A(n22288), .Z(n22285) );
  AND U30186 ( .A(a[18]), .B(b[75]), .Z(n22284) );
  XOR U30187 ( .A(n22290), .B(n22291), .Z(n21737) );
  ANDN U30188 ( .B(n22292), .A(n22293), .Z(n22290) );
  AND U30189 ( .A(a[19]), .B(b[74]), .Z(n22289) );
  XOR U30190 ( .A(n22295), .B(n22296), .Z(n21742) );
  ANDN U30191 ( .B(n22297), .A(n22298), .Z(n22295) );
  AND U30192 ( .A(a[20]), .B(b[73]), .Z(n22294) );
  XOR U30193 ( .A(n22300), .B(n22301), .Z(n21747) );
  ANDN U30194 ( .B(n22302), .A(n22303), .Z(n22300) );
  AND U30195 ( .A(a[21]), .B(b[72]), .Z(n22299) );
  XOR U30196 ( .A(n22305), .B(n22306), .Z(n21752) );
  ANDN U30197 ( .B(n22307), .A(n22308), .Z(n22305) );
  AND U30198 ( .A(a[22]), .B(b[71]), .Z(n22304) );
  XOR U30199 ( .A(n22310), .B(n22311), .Z(n21757) );
  ANDN U30200 ( .B(n22312), .A(n22313), .Z(n22310) );
  AND U30201 ( .A(a[23]), .B(b[70]), .Z(n22309) );
  XOR U30202 ( .A(n22315), .B(n22316), .Z(n21762) );
  ANDN U30203 ( .B(n22317), .A(n22318), .Z(n22315) );
  AND U30204 ( .A(a[24]), .B(b[69]), .Z(n22314) );
  XOR U30205 ( .A(n22320), .B(n22321), .Z(n21767) );
  ANDN U30206 ( .B(n22322), .A(n22323), .Z(n22320) );
  AND U30207 ( .A(a[25]), .B(b[68]), .Z(n22319) );
  XOR U30208 ( .A(n22325), .B(n22326), .Z(n21772) );
  ANDN U30209 ( .B(n22327), .A(n22328), .Z(n22325) );
  AND U30210 ( .A(a[26]), .B(b[67]), .Z(n22324) );
  XOR U30211 ( .A(n22330), .B(n22331), .Z(n21777) );
  ANDN U30212 ( .B(n22332), .A(n22333), .Z(n22330) );
  AND U30213 ( .A(a[27]), .B(b[66]), .Z(n22329) );
  XOR U30214 ( .A(n22335), .B(n22336), .Z(n21782) );
  ANDN U30215 ( .B(n22337), .A(n22338), .Z(n22335) );
  AND U30216 ( .A(a[28]), .B(b[65]), .Z(n22334) );
  XOR U30217 ( .A(n22340), .B(n22341), .Z(n21787) );
  ANDN U30218 ( .B(n22342), .A(n22343), .Z(n22340) );
  AND U30219 ( .A(a[29]), .B(b[64]), .Z(n22339) );
  XOR U30220 ( .A(n22345), .B(n22346), .Z(n21792) );
  ANDN U30221 ( .B(n22347), .A(n22348), .Z(n22345) );
  AND U30222 ( .A(a[30]), .B(b[63]), .Z(n22344) );
  XOR U30223 ( .A(n22350), .B(n22351), .Z(n21797) );
  ANDN U30224 ( .B(n22352), .A(n22353), .Z(n22350) );
  AND U30225 ( .A(a[31]), .B(b[62]), .Z(n22349) );
  XOR U30226 ( .A(n22355), .B(n22356), .Z(n21802) );
  ANDN U30227 ( .B(n22357), .A(n22358), .Z(n22355) );
  AND U30228 ( .A(a[32]), .B(b[61]), .Z(n22354) );
  XOR U30229 ( .A(n22360), .B(n22361), .Z(n21807) );
  ANDN U30230 ( .B(n22362), .A(n22363), .Z(n22360) );
  AND U30231 ( .A(a[33]), .B(b[60]), .Z(n22359) );
  XOR U30232 ( .A(n22365), .B(n22366), .Z(n21812) );
  ANDN U30233 ( .B(n22367), .A(n22368), .Z(n22365) );
  AND U30234 ( .A(a[34]), .B(b[59]), .Z(n22364) );
  XOR U30235 ( .A(n22370), .B(n22371), .Z(n21817) );
  ANDN U30236 ( .B(n22372), .A(n22373), .Z(n22370) );
  AND U30237 ( .A(a[35]), .B(b[58]), .Z(n22369) );
  XOR U30238 ( .A(n22375), .B(n22376), .Z(n21822) );
  ANDN U30239 ( .B(n22377), .A(n22378), .Z(n22375) );
  AND U30240 ( .A(a[36]), .B(b[57]), .Z(n22374) );
  XOR U30241 ( .A(n22380), .B(n22381), .Z(n21827) );
  ANDN U30242 ( .B(n22382), .A(n22383), .Z(n22380) );
  AND U30243 ( .A(a[37]), .B(b[56]), .Z(n22379) );
  XOR U30244 ( .A(n22385), .B(n22386), .Z(n21832) );
  ANDN U30245 ( .B(n22387), .A(n22388), .Z(n22385) );
  AND U30246 ( .A(a[38]), .B(b[55]), .Z(n22384) );
  XOR U30247 ( .A(n22390), .B(n22391), .Z(n21837) );
  ANDN U30248 ( .B(n22392), .A(n22393), .Z(n22390) );
  AND U30249 ( .A(a[39]), .B(b[54]), .Z(n22389) );
  XOR U30250 ( .A(n22395), .B(n22396), .Z(n21842) );
  ANDN U30251 ( .B(n22397), .A(n22398), .Z(n22395) );
  AND U30252 ( .A(a[40]), .B(b[53]), .Z(n22394) );
  XOR U30253 ( .A(n22400), .B(n22401), .Z(n21847) );
  ANDN U30254 ( .B(n22402), .A(n22403), .Z(n22400) );
  AND U30255 ( .A(a[41]), .B(b[52]), .Z(n22399) );
  XOR U30256 ( .A(n22405), .B(n22406), .Z(n21852) );
  ANDN U30257 ( .B(n22407), .A(n22408), .Z(n22405) );
  AND U30258 ( .A(a[42]), .B(b[51]), .Z(n22404) );
  XOR U30259 ( .A(n22410), .B(n22411), .Z(n21857) );
  ANDN U30260 ( .B(n22412), .A(n22413), .Z(n22410) );
  AND U30261 ( .A(a[43]), .B(b[50]), .Z(n22409) );
  XOR U30262 ( .A(n22415), .B(n22416), .Z(n21862) );
  ANDN U30263 ( .B(n22417), .A(n22418), .Z(n22415) );
  AND U30264 ( .A(a[44]), .B(b[49]), .Z(n22414) );
  XOR U30265 ( .A(n22420), .B(n22421), .Z(n21867) );
  ANDN U30266 ( .B(n22422), .A(n22423), .Z(n22420) );
  AND U30267 ( .A(a[45]), .B(b[48]), .Z(n22419) );
  XOR U30268 ( .A(n22425), .B(n22426), .Z(n21872) );
  ANDN U30269 ( .B(n22427), .A(n22428), .Z(n22425) );
  AND U30270 ( .A(a[46]), .B(b[47]), .Z(n22424) );
  XOR U30271 ( .A(n22430), .B(n22431), .Z(n21877) );
  ANDN U30272 ( .B(n22432), .A(n22433), .Z(n22430) );
  AND U30273 ( .A(a[47]), .B(b[46]), .Z(n22429) );
  XOR U30274 ( .A(n22435), .B(n22436), .Z(n21882) );
  ANDN U30275 ( .B(n22437), .A(n22438), .Z(n22435) );
  AND U30276 ( .A(a[48]), .B(b[45]), .Z(n22434) );
  XOR U30277 ( .A(n22440), .B(n22441), .Z(n21887) );
  ANDN U30278 ( .B(n22442), .A(n22443), .Z(n22440) );
  AND U30279 ( .A(a[49]), .B(b[44]), .Z(n22439) );
  XOR U30280 ( .A(n22445), .B(n22446), .Z(n21892) );
  ANDN U30281 ( .B(n22447), .A(n22448), .Z(n22445) );
  AND U30282 ( .A(a[50]), .B(b[43]), .Z(n22444) );
  XOR U30283 ( .A(n22450), .B(n22451), .Z(n21897) );
  ANDN U30284 ( .B(n22452), .A(n22453), .Z(n22450) );
  AND U30285 ( .A(a[51]), .B(b[42]), .Z(n22449) );
  XOR U30286 ( .A(n22455), .B(n22456), .Z(n21902) );
  ANDN U30287 ( .B(n22457), .A(n22458), .Z(n22455) );
  AND U30288 ( .A(a[52]), .B(b[41]), .Z(n22454) );
  XOR U30289 ( .A(n22460), .B(n22461), .Z(n21907) );
  ANDN U30290 ( .B(n22462), .A(n22463), .Z(n22460) );
  AND U30291 ( .A(a[53]), .B(b[40]), .Z(n22459) );
  XOR U30292 ( .A(n22465), .B(n22466), .Z(n21912) );
  ANDN U30293 ( .B(n22467), .A(n22468), .Z(n22465) );
  AND U30294 ( .A(a[54]), .B(b[39]), .Z(n22464) );
  XOR U30295 ( .A(n22470), .B(n22471), .Z(n21917) );
  ANDN U30296 ( .B(n22472), .A(n22473), .Z(n22470) );
  AND U30297 ( .A(a[55]), .B(b[38]), .Z(n22469) );
  XOR U30298 ( .A(n22475), .B(n22476), .Z(n21922) );
  ANDN U30299 ( .B(n22477), .A(n22478), .Z(n22475) );
  AND U30300 ( .A(a[56]), .B(b[37]), .Z(n22474) );
  XOR U30301 ( .A(n22480), .B(n22481), .Z(n21927) );
  ANDN U30302 ( .B(n22482), .A(n22483), .Z(n22480) );
  AND U30303 ( .A(a[57]), .B(b[36]), .Z(n22479) );
  XOR U30304 ( .A(n22485), .B(n22486), .Z(n21932) );
  ANDN U30305 ( .B(n22487), .A(n22488), .Z(n22485) );
  AND U30306 ( .A(a[58]), .B(b[35]), .Z(n22484) );
  XOR U30307 ( .A(n22490), .B(n22491), .Z(n21937) );
  ANDN U30308 ( .B(n22492), .A(n22493), .Z(n22490) );
  AND U30309 ( .A(a[59]), .B(b[34]), .Z(n22489) );
  XOR U30310 ( .A(n22495), .B(n22496), .Z(n21942) );
  ANDN U30311 ( .B(n22497), .A(n22498), .Z(n22495) );
  AND U30312 ( .A(a[60]), .B(b[33]), .Z(n22494) );
  XOR U30313 ( .A(n22500), .B(n22501), .Z(n21947) );
  ANDN U30314 ( .B(n22502), .A(n22503), .Z(n22500) );
  AND U30315 ( .A(a[61]), .B(b[32]), .Z(n22499) );
  XOR U30316 ( .A(n22505), .B(n22506), .Z(n21952) );
  ANDN U30317 ( .B(n22507), .A(n22508), .Z(n22505) );
  AND U30318 ( .A(a[62]), .B(b[31]), .Z(n22504) );
  XOR U30319 ( .A(n22510), .B(n22511), .Z(n21957) );
  ANDN U30320 ( .B(n22512), .A(n22513), .Z(n22510) );
  AND U30321 ( .A(a[63]), .B(b[30]), .Z(n22509) );
  XOR U30322 ( .A(n22515), .B(n22516), .Z(n21962) );
  ANDN U30323 ( .B(n22517), .A(n22518), .Z(n22515) );
  AND U30324 ( .A(a[64]), .B(b[29]), .Z(n22514) );
  XOR U30325 ( .A(n22520), .B(n22521), .Z(n21967) );
  ANDN U30326 ( .B(n22522), .A(n22523), .Z(n22520) );
  AND U30327 ( .A(a[65]), .B(b[28]), .Z(n22519) );
  XOR U30328 ( .A(n22525), .B(n22526), .Z(n21972) );
  ANDN U30329 ( .B(n22527), .A(n22528), .Z(n22525) );
  AND U30330 ( .A(a[66]), .B(b[27]), .Z(n22524) );
  XOR U30331 ( .A(n22530), .B(n22531), .Z(n21977) );
  ANDN U30332 ( .B(n22532), .A(n22533), .Z(n22530) );
  AND U30333 ( .A(a[67]), .B(b[26]), .Z(n22529) );
  XOR U30334 ( .A(n22535), .B(n22536), .Z(n21982) );
  ANDN U30335 ( .B(n22537), .A(n22538), .Z(n22535) );
  AND U30336 ( .A(a[68]), .B(b[25]), .Z(n22534) );
  XOR U30337 ( .A(n22540), .B(n22541), .Z(n21987) );
  ANDN U30338 ( .B(n22542), .A(n22543), .Z(n22540) );
  AND U30339 ( .A(a[69]), .B(b[24]), .Z(n22539) );
  XOR U30340 ( .A(n22545), .B(n22546), .Z(n21992) );
  ANDN U30341 ( .B(n22547), .A(n22548), .Z(n22545) );
  AND U30342 ( .A(a[70]), .B(b[23]), .Z(n22544) );
  XOR U30343 ( .A(n22550), .B(n22551), .Z(n21997) );
  ANDN U30344 ( .B(n22552), .A(n22553), .Z(n22550) );
  AND U30345 ( .A(a[71]), .B(b[22]), .Z(n22549) );
  XOR U30346 ( .A(n22555), .B(n22556), .Z(n22002) );
  ANDN U30347 ( .B(n22557), .A(n22558), .Z(n22555) );
  AND U30348 ( .A(a[72]), .B(b[21]), .Z(n22554) );
  XOR U30349 ( .A(n22560), .B(n22561), .Z(n22007) );
  ANDN U30350 ( .B(n22562), .A(n22563), .Z(n22560) );
  AND U30351 ( .A(a[73]), .B(b[20]), .Z(n22559) );
  XOR U30352 ( .A(n22565), .B(n22566), .Z(n22012) );
  ANDN U30353 ( .B(n22567), .A(n22568), .Z(n22565) );
  AND U30354 ( .A(a[74]), .B(b[19]), .Z(n22564) );
  XOR U30355 ( .A(n22570), .B(n22571), .Z(n22017) );
  ANDN U30356 ( .B(n22572), .A(n22573), .Z(n22570) );
  AND U30357 ( .A(a[75]), .B(b[18]), .Z(n22569) );
  XOR U30358 ( .A(n22575), .B(n22576), .Z(n22022) );
  ANDN U30359 ( .B(n22577), .A(n22578), .Z(n22575) );
  AND U30360 ( .A(a[76]), .B(b[17]), .Z(n22574) );
  XOR U30361 ( .A(n22580), .B(n22581), .Z(n22027) );
  ANDN U30362 ( .B(n22582), .A(n22583), .Z(n22580) );
  AND U30363 ( .A(a[77]), .B(b[16]), .Z(n22579) );
  XOR U30364 ( .A(n22585), .B(n22586), .Z(n22032) );
  ANDN U30365 ( .B(n22587), .A(n22588), .Z(n22585) );
  AND U30366 ( .A(a[78]), .B(b[15]), .Z(n22584) );
  XOR U30367 ( .A(n22590), .B(n22591), .Z(n22037) );
  ANDN U30368 ( .B(n22592), .A(n22593), .Z(n22590) );
  AND U30369 ( .A(a[79]), .B(b[14]), .Z(n22589) );
  XOR U30370 ( .A(n22595), .B(n22596), .Z(n22042) );
  ANDN U30371 ( .B(n22597), .A(n22598), .Z(n22595) );
  AND U30372 ( .A(a[80]), .B(b[13]), .Z(n22594) );
  XOR U30373 ( .A(n22600), .B(n22601), .Z(n22047) );
  ANDN U30374 ( .B(n22602), .A(n22603), .Z(n22600) );
  AND U30375 ( .A(a[81]), .B(b[12]), .Z(n22599) );
  XOR U30376 ( .A(n22605), .B(n22606), .Z(n22052) );
  ANDN U30377 ( .B(n22607), .A(n22608), .Z(n22605) );
  AND U30378 ( .A(a[82]), .B(b[11]), .Z(n22604) );
  XOR U30379 ( .A(n22610), .B(n22611), .Z(n22057) );
  ANDN U30380 ( .B(n22612), .A(n22613), .Z(n22610) );
  AND U30381 ( .A(a[83]), .B(b[10]), .Z(n22609) );
  XOR U30382 ( .A(n22615), .B(n22616), .Z(n22062) );
  ANDN U30383 ( .B(n22617), .A(n22618), .Z(n22615) );
  AND U30384 ( .A(b[9]), .B(a[84]), .Z(n22614) );
  XOR U30385 ( .A(n22620), .B(n22621), .Z(n22067) );
  ANDN U30386 ( .B(n22622), .A(n22623), .Z(n22620) );
  AND U30387 ( .A(b[8]), .B(a[85]), .Z(n22619) );
  XOR U30388 ( .A(n22625), .B(n22626), .Z(n22072) );
  ANDN U30389 ( .B(n22627), .A(n22628), .Z(n22625) );
  AND U30390 ( .A(b[7]), .B(a[86]), .Z(n22624) );
  XOR U30391 ( .A(n22630), .B(n22631), .Z(n22077) );
  ANDN U30392 ( .B(n22632), .A(n22633), .Z(n22630) );
  AND U30393 ( .A(b[6]), .B(a[87]), .Z(n22629) );
  XOR U30394 ( .A(n22635), .B(n22636), .Z(n22082) );
  ANDN U30395 ( .B(n22637), .A(n22638), .Z(n22635) );
  AND U30396 ( .A(b[5]), .B(a[88]), .Z(n22634) );
  XOR U30397 ( .A(n22640), .B(n22641), .Z(n22087) );
  ANDN U30398 ( .B(n22642), .A(n22643), .Z(n22640) );
  AND U30399 ( .A(b[4]), .B(a[89]), .Z(n22639) );
  XOR U30400 ( .A(n22645), .B(n22646), .Z(n22092) );
  ANDN U30401 ( .B(n22104), .A(n22105), .Z(n22645) );
  AND U30402 ( .A(b[2]), .B(a[90]), .Z(n22647) );
  XNOR U30403 ( .A(n22642), .B(n22646), .Z(n22648) );
  XOR U30404 ( .A(n22649), .B(n22650), .Z(n22646) );
  OR U30405 ( .A(n22107), .B(n22108), .Z(n22650) );
  XNOR U30406 ( .A(n22652), .B(n22653), .Z(n22651) );
  XOR U30407 ( .A(n22652), .B(n22655), .Z(n22107) );
  NAND U30408 ( .A(b[1]), .B(a[90]), .Z(n22655) );
  IV U30409 ( .A(n22649), .Z(n22652) );
  NANDN U30410 ( .A(n21), .B(n22), .Z(n22649) );
  XOR U30411 ( .A(n22656), .B(n22657), .Z(n22) );
  NAND U30412 ( .A(a[90]), .B(b[0]), .Z(n21) );
  XNOR U30413 ( .A(n22637), .B(n22641), .Z(n22658) );
  XNOR U30414 ( .A(n22632), .B(n22636), .Z(n22659) );
  XNOR U30415 ( .A(n22627), .B(n22631), .Z(n22660) );
  XNOR U30416 ( .A(n22622), .B(n22626), .Z(n22661) );
  XNOR U30417 ( .A(n22617), .B(n22621), .Z(n22662) );
  XNOR U30418 ( .A(n22612), .B(n22616), .Z(n22663) );
  XNOR U30419 ( .A(n22607), .B(n22611), .Z(n22664) );
  XNOR U30420 ( .A(n22602), .B(n22606), .Z(n22665) );
  XNOR U30421 ( .A(n22597), .B(n22601), .Z(n22666) );
  XNOR U30422 ( .A(n22592), .B(n22596), .Z(n22667) );
  XNOR U30423 ( .A(n22587), .B(n22591), .Z(n22668) );
  XNOR U30424 ( .A(n22582), .B(n22586), .Z(n22669) );
  XNOR U30425 ( .A(n22577), .B(n22581), .Z(n22670) );
  XNOR U30426 ( .A(n22572), .B(n22576), .Z(n22671) );
  XNOR U30427 ( .A(n22567), .B(n22571), .Z(n22672) );
  XNOR U30428 ( .A(n22562), .B(n22566), .Z(n22673) );
  XNOR U30429 ( .A(n22557), .B(n22561), .Z(n22674) );
  XNOR U30430 ( .A(n22552), .B(n22556), .Z(n22675) );
  XNOR U30431 ( .A(n22547), .B(n22551), .Z(n22676) );
  XNOR U30432 ( .A(n22542), .B(n22546), .Z(n22677) );
  XNOR U30433 ( .A(n22537), .B(n22541), .Z(n22678) );
  XNOR U30434 ( .A(n22532), .B(n22536), .Z(n22679) );
  XNOR U30435 ( .A(n22527), .B(n22531), .Z(n22680) );
  XNOR U30436 ( .A(n22522), .B(n22526), .Z(n22681) );
  XNOR U30437 ( .A(n22517), .B(n22521), .Z(n22682) );
  XNOR U30438 ( .A(n22512), .B(n22516), .Z(n22683) );
  XNOR U30439 ( .A(n22507), .B(n22511), .Z(n22684) );
  XNOR U30440 ( .A(n22502), .B(n22506), .Z(n22685) );
  XNOR U30441 ( .A(n22497), .B(n22501), .Z(n22686) );
  XNOR U30442 ( .A(n22492), .B(n22496), .Z(n22687) );
  XNOR U30443 ( .A(n22487), .B(n22491), .Z(n22688) );
  XNOR U30444 ( .A(n22482), .B(n22486), .Z(n22689) );
  XNOR U30445 ( .A(n22477), .B(n22481), .Z(n22690) );
  XNOR U30446 ( .A(n22472), .B(n22476), .Z(n22691) );
  XNOR U30447 ( .A(n22467), .B(n22471), .Z(n22692) );
  XNOR U30448 ( .A(n22462), .B(n22466), .Z(n22693) );
  XNOR U30449 ( .A(n22457), .B(n22461), .Z(n22694) );
  XNOR U30450 ( .A(n22452), .B(n22456), .Z(n22695) );
  XNOR U30451 ( .A(n22447), .B(n22451), .Z(n22696) );
  XNOR U30452 ( .A(n22442), .B(n22446), .Z(n22697) );
  XNOR U30453 ( .A(n22437), .B(n22441), .Z(n22698) );
  XNOR U30454 ( .A(n22432), .B(n22436), .Z(n22699) );
  XNOR U30455 ( .A(n22427), .B(n22431), .Z(n22700) );
  XNOR U30456 ( .A(n22422), .B(n22426), .Z(n22701) );
  XNOR U30457 ( .A(n22417), .B(n22421), .Z(n22702) );
  XNOR U30458 ( .A(n22412), .B(n22416), .Z(n22703) );
  XNOR U30459 ( .A(n22407), .B(n22411), .Z(n22704) );
  XNOR U30460 ( .A(n22402), .B(n22406), .Z(n22705) );
  XNOR U30461 ( .A(n22397), .B(n22401), .Z(n22706) );
  XNOR U30462 ( .A(n22392), .B(n22396), .Z(n22707) );
  XNOR U30463 ( .A(n22387), .B(n22391), .Z(n22708) );
  XNOR U30464 ( .A(n22382), .B(n22386), .Z(n22709) );
  XNOR U30465 ( .A(n22377), .B(n22381), .Z(n22710) );
  XNOR U30466 ( .A(n22372), .B(n22376), .Z(n22711) );
  XNOR U30467 ( .A(n22367), .B(n22371), .Z(n22712) );
  XNOR U30468 ( .A(n22362), .B(n22366), .Z(n22713) );
  XNOR U30469 ( .A(n22357), .B(n22361), .Z(n22714) );
  XNOR U30470 ( .A(n22352), .B(n22356), .Z(n22715) );
  XNOR U30471 ( .A(n22716), .B(n22717), .Z(n22352) );
  XNOR U30472 ( .A(n22347), .B(n22351), .Z(n22717) );
  XNOR U30473 ( .A(n22342), .B(n22346), .Z(n22718) );
  XNOR U30474 ( .A(n22337), .B(n22341), .Z(n22719) );
  XNOR U30475 ( .A(n22332), .B(n22336), .Z(n22720) );
  XNOR U30476 ( .A(n22327), .B(n22331), .Z(n22721) );
  XNOR U30477 ( .A(n22322), .B(n22326), .Z(n22722) );
  XNOR U30478 ( .A(n22317), .B(n22321), .Z(n22723) );
  XNOR U30479 ( .A(n22312), .B(n22316), .Z(n22724) );
  XNOR U30480 ( .A(n22307), .B(n22311), .Z(n22725) );
  XNOR U30481 ( .A(n22302), .B(n22306), .Z(n22726) );
  XNOR U30482 ( .A(n22297), .B(n22301), .Z(n22727) );
  XNOR U30483 ( .A(n22292), .B(n22296), .Z(n22728) );
  XNOR U30484 ( .A(n22287), .B(n22291), .Z(n22729) );
  XNOR U30485 ( .A(n22282), .B(n22286), .Z(n22730) );
  XNOR U30486 ( .A(n22277), .B(n22281), .Z(n22731) );
  XNOR U30487 ( .A(n22272), .B(n22276), .Z(n22732) );
  XNOR U30488 ( .A(n22267), .B(n22271), .Z(n22733) );
  XNOR U30489 ( .A(n22262), .B(n22266), .Z(n22734) );
  XNOR U30490 ( .A(n22257), .B(n22261), .Z(n22735) );
  XNOR U30491 ( .A(n22252), .B(n22256), .Z(n22736) );
  XNOR U30492 ( .A(n22247), .B(n22251), .Z(n22737) );
  XNOR U30493 ( .A(n22242), .B(n22246), .Z(n22738) );
  XNOR U30494 ( .A(n22237), .B(n22241), .Z(n22739) );
  XNOR U30495 ( .A(n22232), .B(n22236), .Z(n22740) );
  XNOR U30496 ( .A(n22227), .B(n22231), .Z(n22741) );
  XNOR U30497 ( .A(n22222), .B(n22226), .Z(n22742) );
  XNOR U30498 ( .A(n22217), .B(n22221), .Z(n22743) );
  XNOR U30499 ( .A(n22212), .B(n22216), .Z(n22744) );
  XNOR U30500 ( .A(n22207), .B(n22211), .Z(n22745) );
  XNOR U30501 ( .A(n22202), .B(n22206), .Z(n22746) );
  XOR U30502 ( .A(n22747), .B(n22201), .Z(n22202) );
  AND U30503 ( .A(a[0]), .B(b[92]), .Z(n22747) );
  XNOR U30504 ( .A(n22748), .B(n22201), .Z(n22203) );
  XNOR U30505 ( .A(n22749), .B(n22750), .Z(n22201) );
  ANDN U30506 ( .B(n22751), .A(n22752), .Z(n22749) );
  AND U30507 ( .A(a[1]), .B(b[91]), .Z(n22748) );
  XOR U30508 ( .A(n22754), .B(n22755), .Z(n22206) );
  ANDN U30509 ( .B(n22756), .A(n22757), .Z(n22754) );
  AND U30510 ( .A(a[2]), .B(b[90]), .Z(n22753) );
  XOR U30511 ( .A(n22759), .B(n22760), .Z(n22211) );
  ANDN U30512 ( .B(n22761), .A(n22762), .Z(n22759) );
  AND U30513 ( .A(a[3]), .B(b[89]), .Z(n22758) );
  XOR U30514 ( .A(n22764), .B(n22765), .Z(n22216) );
  ANDN U30515 ( .B(n22766), .A(n22767), .Z(n22764) );
  AND U30516 ( .A(a[4]), .B(b[88]), .Z(n22763) );
  XOR U30517 ( .A(n22769), .B(n22770), .Z(n22221) );
  ANDN U30518 ( .B(n22771), .A(n22772), .Z(n22769) );
  AND U30519 ( .A(a[5]), .B(b[87]), .Z(n22768) );
  XOR U30520 ( .A(n22774), .B(n22775), .Z(n22226) );
  ANDN U30521 ( .B(n22776), .A(n22777), .Z(n22774) );
  AND U30522 ( .A(a[6]), .B(b[86]), .Z(n22773) );
  XOR U30523 ( .A(n22779), .B(n22780), .Z(n22231) );
  ANDN U30524 ( .B(n22781), .A(n22782), .Z(n22779) );
  AND U30525 ( .A(a[7]), .B(b[85]), .Z(n22778) );
  XOR U30526 ( .A(n22784), .B(n22785), .Z(n22236) );
  ANDN U30527 ( .B(n22786), .A(n22787), .Z(n22784) );
  AND U30528 ( .A(a[8]), .B(b[84]), .Z(n22783) );
  XOR U30529 ( .A(n22789), .B(n22790), .Z(n22241) );
  ANDN U30530 ( .B(n22791), .A(n22792), .Z(n22789) );
  AND U30531 ( .A(a[9]), .B(b[83]), .Z(n22788) );
  XOR U30532 ( .A(n22794), .B(n22795), .Z(n22246) );
  ANDN U30533 ( .B(n22796), .A(n22797), .Z(n22794) );
  AND U30534 ( .A(a[10]), .B(b[82]), .Z(n22793) );
  XOR U30535 ( .A(n22799), .B(n22800), .Z(n22251) );
  ANDN U30536 ( .B(n22801), .A(n22802), .Z(n22799) );
  AND U30537 ( .A(a[11]), .B(b[81]), .Z(n22798) );
  XOR U30538 ( .A(n22804), .B(n22805), .Z(n22256) );
  ANDN U30539 ( .B(n22806), .A(n22807), .Z(n22804) );
  AND U30540 ( .A(a[12]), .B(b[80]), .Z(n22803) );
  XOR U30541 ( .A(n22809), .B(n22810), .Z(n22261) );
  ANDN U30542 ( .B(n22811), .A(n22812), .Z(n22809) );
  AND U30543 ( .A(a[13]), .B(b[79]), .Z(n22808) );
  XOR U30544 ( .A(n22814), .B(n22815), .Z(n22266) );
  ANDN U30545 ( .B(n22816), .A(n22817), .Z(n22814) );
  AND U30546 ( .A(a[14]), .B(b[78]), .Z(n22813) );
  XOR U30547 ( .A(n22819), .B(n22820), .Z(n22271) );
  ANDN U30548 ( .B(n22821), .A(n22822), .Z(n22819) );
  AND U30549 ( .A(a[15]), .B(b[77]), .Z(n22818) );
  XOR U30550 ( .A(n22824), .B(n22825), .Z(n22276) );
  ANDN U30551 ( .B(n22826), .A(n22827), .Z(n22824) );
  AND U30552 ( .A(a[16]), .B(b[76]), .Z(n22823) );
  XOR U30553 ( .A(n22829), .B(n22830), .Z(n22281) );
  ANDN U30554 ( .B(n22831), .A(n22832), .Z(n22829) );
  AND U30555 ( .A(a[17]), .B(b[75]), .Z(n22828) );
  XOR U30556 ( .A(n22834), .B(n22835), .Z(n22286) );
  ANDN U30557 ( .B(n22836), .A(n22837), .Z(n22834) );
  AND U30558 ( .A(a[18]), .B(b[74]), .Z(n22833) );
  XOR U30559 ( .A(n22839), .B(n22840), .Z(n22291) );
  ANDN U30560 ( .B(n22841), .A(n22842), .Z(n22839) );
  AND U30561 ( .A(a[19]), .B(b[73]), .Z(n22838) );
  XOR U30562 ( .A(n22844), .B(n22845), .Z(n22296) );
  ANDN U30563 ( .B(n22846), .A(n22847), .Z(n22844) );
  AND U30564 ( .A(a[20]), .B(b[72]), .Z(n22843) );
  XOR U30565 ( .A(n22849), .B(n22850), .Z(n22301) );
  ANDN U30566 ( .B(n22851), .A(n22852), .Z(n22849) );
  AND U30567 ( .A(a[21]), .B(b[71]), .Z(n22848) );
  XOR U30568 ( .A(n22854), .B(n22855), .Z(n22306) );
  ANDN U30569 ( .B(n22856), .A(n22857), .Z(n22854) );
  AND U30570 ( .A(a[22]), .B(b[70]), .Z(n22853) );
  XOR U30571 ( .A(n22859), .B(n22860), .Z(n22311) );
  ANDN U30572 ( .B(n22861), .A(n22862), .Z(n22859) );
  AND U30573 ( .A(a[23]), .B(b[69]), .Z(n22858) );
  XOR U30574 ( .A(n22864), .B(n22865), .Z(n22316) );
  ANDN U30575 ( .B(n22866), .A(n22867), .Z(n22864) );
  AND U30576 ( .A(a[24]), .B(b[68]), .Z(n22863) );
  XOR U30577 ( .A(n22869), .B(n22870), .Z(n22321) );
  ANDN U30578 ( .B(n22871), .A(n22872), .Z(n22869) );
  AND U30579 ( .A(a[25]), .B(b[67]), .Z(n22868) );
  XOR U30580 ( .A(n22874), .B(n22875), .Z(n22326) );
  ANDN U30581 ( .B(n22876), .A(n22877), .Z(n22874) );
  AND U30582 ( .A(a[26]), .B(b[66]), .Z(n22873) );
  XOR U30583 ( .A(n22879), .B(n22880), .Z(n22331) );
  ANDN U30584 ( .B(n22881), .A(n22882), .Z(n22879) );
  AND U30585 ( .A(a[27]), .B(b[65]), .Z(n22878) );
  XOR U30586 ( .A(n22884), .B(n22885), .Z(n22336) );
  ANDN U30587 ( .B(n22886), .A(n22887), .Z(n22884) );
  AND U30588 ( .A(a[28]), .B(b[64]), .Z(n22883) );
  XOR U30589 ( .A(n22889), .B(n22890), .Z(n22341) );
  ANDN U30590 ( .B(n22891), .A(n22892), .Z(n22889) );
  AND U30591 ( .A(a[29]), .B(b[63]), .Z(n22888) );
  IV U30592 ( .A(n22348), .Z(n22716) );
  XOR U30593 ( .A(n22894), .B(n22895), .Z(n22346) );
  ANDN U30594 ( .B(n22896), .A(n22897), .Z(n22894) );
  AND U30595 ( .A(a[30]), .B(b[62]), .Z(n22893) );
  XOR U30596 ( .A(n22899), .B(n22900), .Z(n22351) );
  ANDN U30597 ( .B(n22901), .A(n22902), .Z(n22899) );
  AND U30598 ( .A(a[31]), .B(b[61]), .Z(n22898) );
  XOR U30599 ( .A(n22904), .B(n22905), .Z(n22356) );
  ANDN U30600 ( .B(n22906), .A(n22907), .Z(n22904) );
  AND U30601 ( .A(a[32]), .B(b[60]), .Z(n22903) );
  XOR U30602 ( .A(n22909), .B(n22910), .Z(n22361) );
  ANDN U30603 ( .B(n22911), .A(n22912), .Z(n22909) );
  AND U30604 ( .A(a[33]), .B(b[59]), .Z(n22908) );
  XOR U30605 ( .A(n22914), .B(n22915), .Z(n22366) );
  ANDN U30606 ( .B(n22916), .A(n22917), .Z(n22914) );
  AND U30607 ( .A(a[34]), .B(b[58]), .Z(n22913) );
  XOR U30608 ( .A(n22919), .B(n22920), .Z(n22371) );
  ANDN U30609 ( .B(n22921), .A(n22922), .Z(n22919) );
  AND U30610 ( .A(a[35]), .B(b[57]), .Z(n22918) );
  XOR U30611 ( .A(n22924), .B(n22925), .Z(n22376) );
  ANDN U30612 ( .B(n22926), .A(n22927), .Z(n22924) );
  AND U30613 ( .A(a[36]), .B(b[56]), .Z(n22923) );
  XOR U30614 ( .A(n22929), .B(n22930), .Z(n22381) );
  ANDN U30615 ( .B(n22931), .A(n22932), .Z(n22929) );
  AND U30616 ( .A(a[37]), .B(b[55]), .Z(n22928) );
  XOR U30617 ( .A(n22934), .B(n22935), .Z(n22386) );
  ANDN U30618 ( .B(n22936), .A(n22937), .Z(n22934) );
  AND U30619 ( .A(a[38]), .B(b[54]), .Z(n22933) );
  XOR U30620 ( .A(n22939), .B(n22940), .Z(n22391) );
  ANDN U30621 ( .B(n22941), .A(n22942), .Z(n22939) );
  AND U30622 ( .A(a[39]), .B(b[53]), .Z(n22938) );
  XOR U30623 ( .A(n22944), .B(n22945), .Z(n22396) );
  ANDN U30624 ( .B(n22946), .A(n22947), .Z(n22944) );
  AND U30625 ( .A(a[40]), .B(b[52]), .Z(n22943) );
  XOR U30626 ( .A(n22949), .B(n22950), .Z(n22401) );
  ANDN U30627 ( .B(n22951), .A(n22952), .Z(n22949) );
  AND U30628 ( .A(a[41]), .B(b[51]), .Z(n22948) );
  XOR U30629 ( .A(n22954), .B(n22955), .Z(n22406) );
  ANDN U30630 ( .B(n22956), .A(n22957), .Z(n22954) );
  AND U30631 ( .A(a[42]), .B(b[50]), .Z(n22953) );
  XOR U30632 ( .A(n22959), .B(n22960), .Z(n22411) );
  ANDN U30633 ( .B(n22961), .A(n22962), .Z(n22959) );
  AND U30634 ( .A(a[43]), .B(b[49]), .Z(n22958) );
  XOR U30635 ( .A(n22964), .B(n22965), .Z(n22416) );
  ANDN U30636 ( .B(n22966), .A(n22967), .Z(n22964) );
  AND U30637 ( .A(a[44]), .B(b[48]), .Z(n22963) );
  XOR U30638 ( .A(n22969), .B(n22970), .Z(n22421) );
  ANDN U30639 ( .B(n22971), .A(n22972), .Z(n22969) );
  AND U30640 ( .A(a[45]), .B(b[47]), .Z(n22968) );
  XOR U30641 ( .A(n22974), .B(n22975), .Z(n22426) );
  ANDN U30642 ( .B(n22976), .A(n22977), .Z(n22974) );
  AND U30643 ( .A(a[46]), .B(b[46]), .Z(n22973) );
  XOR U30644 ( .A(n22979), .B(n22980), .Z(n22431) );
  ANDN U30645 ( .B(n22981), .A(n22982), .Z(n22979) );
  AND U30646 ( .A(a[47]), .B(b[45]), .Z(n22978) );
  XOR U30647 ( .A(n22984), .B(n22985), .Z(n22436) );
  ANDN U30648 ( .B(n22986), .A(n22987), .Z(n22984) );
  AND U30649 ( .A(a[48]), .B(b[44]), .Z(n22983) );
  XOR U30650 ( .A(n22989), .B(n22990), .Z(n22441) );
  ANDN U30651 ( .B(n22991), .A(n22992), .Z(n22989) );
  AND U30652 ( .A(a[49]), .B(b[43]), .Z(n22988) );
  XOR U30653 ( .A(n22994), .B(n22995), .Z(n22446) );
  ANDN U30654 ( .B(n22996), .A(n22997), .Z(n22994) );
  AND U30655 ( .A(a[50]), .B(b[42]), .Z(n22993) );
  XOR U30656 ( .A(n22999), .B(n23000), .Z(n22451) );
  ANDN U30657 ( .B(n23001), .A(n23002), .Z(n22999) );
  AND U30658 ( .A(a[51]), .B(b[41]), .Z(n22998) );
  XOR U30659 ( .A(n23004), .B(n23005), .Z(n22456) );
  ANDN U30660 ( .B(n23006), .A(n23007), .Z(n23004) );
  AND U30661 ( .A(a[52]), .B(b[40]), .Z(n23003) );
  XOR U30662 ( .A(n23009), .B(n23010), .Z(n22461) );
  ANDN U30663 ( .B(n23011), .A(n23012), .Z(n23009) );
  AND U30664 ( .A(a[53]), .B(b[39]), .Z(n23008) );
  XOR U30665 ( .A(n23014), .B(n23015), .Z(n22466) );
  ANDN U30666 ( .B(n23016), .A(n23017), .Z(n23014) );
  AND U30667 ( .A(a[54]), .B(b[38]), .Z(n23013) );
  XOR U30668 ( .A(n23019), .B(n23020), .Z(n22471) );
  ANDN U30669 ( .B(n23021), .A(n23022), .Z(n23019) );
  AND U30670 ( .A(a[55]), .B(b[37]), .Z(n23018) );
  XOR U30671 ( .A(n23024), .B(n23025), .Z(n22476) );
  ANDN U30672 ( .B(n23026), .A(n23027), .Z(n23024) );
  AND U30673 ( .A(a[56]), .B(b[36]), .Z(n23023) );
  XOR U30674 ( .A(n23029), .B(n23030), .Z(n22481) );
  ANDN U30675 ( .B(n23031), .A(n23032), .Z(n23029) );
  AND U30676 ( .A(a[57]), .B(b[35]), .Z(n23028) );
  XOR U30677 ( .A(n23034), .B(n23035), .Z(n22486) );
  ANDN U30678 ( .B(n23036), .A(n23037), .Z(n23034) );
  AND U30679 ( .A(a[58]), .B(b[34]), .Z(n23033) );
  XOR U30680 ( .A(n23039), .B(n23040), .Z(n22491) );
  ANDN U30681 ( .B(n23041), .A(n23042), .Z(n23039) );
  AND U30682 ( .A(a[59]), .B(b[33]), .Z(n23038) );
  XOR U30683 ( .A(n23044), .B(n23045), .Z(n22496) );
  ANDN U30684 ( .B(n23046), .A(n23047), .Z(n23044) );
  AND U30685 ( .A(a[60]), .B(b[32]), .Z(n23043) );
  XOR U30686 ( .A(n23049), .B(n23050), .Z(n22501) );
  ANDN U30687 ( .B(n23051), .A(n23052), .Z(n23049) );
  AND U30688 ( .A(a[61]), .B(b[31]), .Z(n23048) );
  XOR U30689 ( .A(n23054), .B(n23055), .Z(n22506) );
  ANDN U30690 ( .B(n23056), .A(n23057), .Z(n23054) );
  AND U30691 ( .A(a[62]), .B(b[30]), .Z(n23053) );
  XOR U30692 ( .A(n23059), .B(n23060), .Z(n22511) );
  ANDN U30693 ( .B(n23061), .A(n23062), .Z(n23059) );
  AND U30694 ( .A(a[63]), .B(b[29]), .Z(n23058) );
  XOR U30695 ( .A(n23064), .B(n23065), .Z(n22516) );
  ANDN U30696 ( .B(n23066), .A(n23067), .Z(n23064) );
  AND U30697 ( .A(a[64]), .B(b[28]), .Z(n23063) );
  XOR U30698 ( .A(n23069), .B(n23070), .Z(n22521) );
  ANDN U30699 ( .B(n23071), .A(n23072), .Z(n23069) );
  AND U30700 ( .A(a[65]), .B(b[27]), .Z(n23068) );
  XOR U30701 ( .A(n23074), .B(n23075), .Z(n22526) );
  ANDN U30702 ( .B(n23076), .A(n23077), .Z(n23074) );
  AND U30703 ( .A(a[66]), .B(b[26]), .Z(n23073) );
  XOR U30704 ( .A(n23079), .B(n23080), .Z(n22531) );
  ANDN U30705 ( .B(n23081), .A(n23082), .Z(n23079) );
  AND U30706 ( .A(a[67]), .B(b[25]), .Z(n23078) );
  XOR U30707 ( .A(n23084), .B(n23085), .Z(n22536) );
  ANDN U30708 ( .B(n23086), .A(n23087), .Z(n23084) );
  AND U30709 ( .A(a[68]), .B(b[24]), .Z(n23083) );
  XOR U30710 ( .A(n23089), .B(n23090), .Z(n22541) );
  ANDN U30711 ( .B(n23091), .A(n23092), .Z(n23089) );
  AND U30712 ( .A(a[69]), .B(b[23]), .Z(n23088) );
  XOR U30713 ( .A(n23094), .B(n23095), .Z(n22546) );
  ANDN U30714 ( .B(n23096), .A(n23097), .Z(n23094) );
  AND U30715 ( .A(a[70]), .B(b[22]), .Z(n23093) );
  XOR U30716 ( .A(n23099), .B(n23100), .Z(n22551) );
  ANDN U30717 ( .B(n23101), .A(n23102), .Z(n23099) );
  AND U30718 ( .A(a[71]), .B(b[21]), .Z(n23098) );
  XOR U30719 ( .A(n23104), .B(n23105), .Z(n22556) );
  ANDN U30720 ( .B(n23106), .A(n23107), .Z(n23104) );
  AND U30721 ( .A(a[72]), .B(b[20]), .Z(n23103) );
  XOR U30722 ( .A(n23109), .B(n23110), .Z(n22561) );
  ANDN U30723 ( .B(n23111), .A(n23112), .Z(n23109) );
  AND U30724 ( .A(a[73]), .B(b[19]), .Z(n23108) );
  XOR U30725 ( .A(n23114), .B(n23115), .Z(n22566) );
  ANDN U30726 ( .B(n23116), .A(n23117), .Z(n23114) );
  AND U30727 ( .A(a[74]), .B(b[18]), .Z(n23113) );
  XOR U30728 ( .A(n23119), .B(n23120), .Z(n22571) );
  ANDN U30729 ( .B(n23121), .A(n23122), .Z(n23119) );
  AND U30730 ( .A(a[75]), .B(b[17]), .Z(n23118) );
  XOR U30731 ( .A(n23124), .B(n23125), .Z(n22576) );
  ANDN U30732 ( .B(n23126), .A(n23127), .Z(n23124) );
  AND U30733 ( .A(a[76]), .B(b[16]), .Z(n23123) );
  XOR U30734 ( .A(n23129), .B(n23130), .Z(n22581) );
  ANDN U30735 ( .B(n23131), .A(n23132), .Z(n23129) );
  AND U30736 ( .A(a[77]), .B(b[15]), .Z(n23128) );
  XOR U30737 ( .A(n23134), .B(n23135), .Z(n22586) );
  ANDN U30738 ( .B(n23136), .A(n23137), .Z(n23134) );
  AND U30739 ( .A(a[78]), .B(b[14]), .Z(n23133) );
  XOR U30740 ( .A(n23139), .B(n23140), .Z(n22591) );
  ANDN U30741 ( .B(n23141), .A(n23142), .Z(n23139) );
  AND U30742 ( .A(a[79]), .B(b[13]), .Z(n23138) );
  XOR U30743 ( .A(n23144), .B(n23145), .Z(n22596) );
  ANDN U30744 ( .B(n23146), .A(n23147), .Z(n23144) );
  AND U30745 ( .A(a[80]), .B(b[12]), .Z(n23143) );
  XOR U30746 ( .A(n23149), .B(n23150), .Z(n22601) );
  ANDN U30747 ( .B(n23151), .A(n23152), .Z(n23149) );
  AND U30748 ( .A(a[81]), .B(b[11]), .Z(n23148) );
  XOR U30749 ( .A(n23154), .B(n23155), .Z(n22606) );
  ANDN U30750 ( .B(n23156), .A(n23157), .Z(n23154) );
  AND U30751 ( .A(a[82]), .B(b[10]), .Z(n23153) );
  XOR U30752 ( .A(n23159), .B(n23160), .Z(n22611) );
  ANDN U30753 ( .B(n23161), .A(n23162), .Z(n23159) );
  AND U30754 ( .A(b[9]), .B(a[83]), .Z(n23158) );
  XOR U30755 ( .A(n23164), .B(n23165), .Z(n22616) );
  ANDN U30756 ( .B(n23166), .A(n23167), .Z(n23164) );
  AND U30757 ( .A(b[8]), .B(a[84]), .Z(n23163) );
  XOR U30758 ( .A(n23169), .B(n23170), .Z(n22621) );
  ANDN U30759 ( .B(n23171), .A(n23172), .Z(n23169) );
  AND U30760 ( .A(b[7]), .B(a[85]), .Z(n23168) );
  XOR U30761 ( .A(n23174), .B(n23175), .Z(n22626) );
  ANDN U30762 ( .B(n23176), .A(n23177), .Z(n23174) );
  AND U30763 ( .A(b[6]), .B(a[86]), .Z(n23173) );
  XOR U30764 ( .A(n23179), .B(n23180), .Z(n22631) );
  ANDN U30765 ( .B(n23181), .A(n23182), .Z(n23179) );
  AND U30766 ( .A(b[5]), .B(a[87]), .Z(n23178) );
  XOR U30767 ( .A(n23184), .B(n23185), .Z(n22636) );
  ANDN U30768 ( .B(n23186), .A(n23187), .Z(n23184) );
  AND U30769 ( .A(b[4]), .B(a[88]), .Z(n23183) );
  XOR U30770 ( .A(n23189), .B(n23190), .Z(n22641) );
  ANDN U30771 ( .B(n22653), .A(n22654), .Z(n23189) );
  AND U30772 ( .A(b[2]), .B(a[89]), .Z(n23191) );
  XNOR U30773 ( .A(n23186), .B(n23190), .Z(n23192) );
  XOR U30774 ( .A(n23193), .B(n23194), .Z(n23190) );
  OR U30775 ( .A(n22656), .B(n22657), .Z(n23194) );
  XNOR U30776 ( .A(n23196), .B(n23197), .Z(n23195) );
  XOR U30777 ( .A(n23196), .B(n23199), .Z(n22656) );
  NAND U30778 ( .A(b[1]), .B(a[89]), .Z(n23199) );
  IV U30779 ( .A(n23193), .Z(n23196) );
  NANDN U30780 ( .A(n25), .B(n26), .Z(n23193) );
  XOR U30781 ( .A(n23200), .B(n23201), .Z(n26) );
  NAND U30782 ( .A(a[89]), .B(b[0]), .Z(n25) );
  XNOR U30783 ( .A(n23181), .B(n23185), .Z(n23202) );
  XNOR U30784 ( .A(n23176), .B(n23180), .Z(n23203) );
  XNOR U30785 ( .A(n23171), .B(n23175), .Z(n23204) );
  XNOR U30786 ( .A(n23166), .B(n23170), .Z(n23205) );
  XNOR U30787 ( .A(n23161), .B(n23165), .Z(n23206) );
  XNOR U30788 ( .A(n23156), .B(n23160), .Z(n23207) );
  XNOR U30789 ( .A(n23151), .B(n23155), .Z(n23208) );
  XNOR U30790 ( .A(n23146), .B(n23150), .Z(n23209) );
  XNOR U30791 ( .A(n23141), .B(n23145), .Z(n23210) );
  XNOR U30792 ( .A(n23136), .B(n23140), .Z(n23211) );
  XNOR U30793 ( .A(n23131), .B(n23135), .Z(n23212) );
  XNOR U30794 ( .A(n23126), .B(n23130), .Z(n23213) );
  XNOR U30795 ( .A(n23121), .B(n23125), .Z(n23214) );
  XNOR U30796 ( .A(n23116), .B(n23120), .Z(n23215) );
  XNOR U30797 ( .A(n23111), .B(n23115), .Z(n23216) );
  XNOR U30798 ( .A(n23106), .B(n23110), .Z(n23217) );
  XNOR U30799 ( .A(n23101), .B(n23105), .Z(n23218) );
  XNOR U30800 ( .A(n23096), .B(n23100), .Z(n23219) );
  XNOR U30801 ( .A(n23091), .B(n23095), .Z(n23220) );
  XNOR U30802 ( .A(n23086), .B(n23090), .Z(n23221) );
  XNOR U30803 ( .A(n23081), .B(n23085), .Z(n23222) );
  XNOR U30804 ( .A(n23076), .B(n23080), .Z(n23223) );
  XNOR U30805 ( .A(n23071), .B(n23075), .Z(n23224) );
  XNOR U30806 ( .A(n23066), .B(n23070), .Z(n23225) );
  XNOR U30807 ( .A(n23061), .B(n23065), .Z(n23226) );
  XNOR U30808 ( .A(n23056), .B(n23060), .Z(n23227) );
  XNOR U30809 ( .A(n23051), .B(n23055), .Z(n23228) );
  XNOR U30810 ( .A(n23046), .B(n23050), .Z(n23229) );
  XNOR U30811 ( .A(n23041), .B(n23045), .Z(n23230) );
  XNOR U30812 ( .A(n23036), .B(n23040), .Z(n23231) );
  XNOR U30813 ( .A(n23031), .B(n23035), .Z(n23232) );
  XNOR U30814 ( .A(n23026), .B(n23030), .Z(n23233) );
  XNOR U30815 ( .A(n23021), .B(n23025), .Z(n23234) );
  XNOR U30816 ( .A(n23016), .B(n23020), .Z(n23235) );
  XNOR U30817 ( .A(n23011), .B(n23015), .Z(n23236) );
  XNOR U30818 ( .A(n23006), .B(n23010), .Z(n23237) );
  XNOR U30819 ( .A(n23001), .B(n23005), .Z(n23238) );
  XNOR U30820 ( .A(n22996), .B(n23000), .Z(n23239) );
  XNOR U30821 ( .A(n22991), .B(n22995), .Z(n23240) );
  XNOR U30822 ( .A(n22986), .B(n22990), .Z(n23241) );
  XNOR U30823 ( .A(n22981), .B(n22985), .Z(n23242) );
  XNOR U30824 ( .A(n22976), .B(n22980), .Z(n23243) );
  XNOR U30825 ( .A(n22971), .B(n22975), .Z(n23244) );
  XNOR U30826 ( .A(n22966), .B(n22970), .Z(n23245) );
  XNOR U30827 ( .A(n22961), .B(n22965), .Z(n23246) );
  XNOR U30828 ( .A(n22956), .B(n22960), .Z(n23247) );
  XNOR U30829 ( .A(n22951), .B(n22955), .Z(n23248) );
  XNOR U30830 ( .A(n22946), .B(n22950), .Z(n23249) );
  XNOR U30831 ( .A(n22941), .B(n22945), .Z(n23250) );
  XNOR U30832 ( .A(n22936), .B(n22940), .Z(n23251) );
  XNOR U30833 ( .A(n22931), .B(n22935), .Z(n23252) );
  XNOR U30834 ( .A(n22926), .B(n22930), .Z(n23253) );
  XNOR U30835 ( .A(n22921), .B(n22925), .Z(n23254) );
  XNOR U30836 ( .A(n22916), .B(n22920), .Z(n23255) );
  XNOR U30837 ( .A(n22911), .B(n22915), .Z(n23256) );
  XNOR U30838 ( .A(n22906), .B(n22910), .Z(n23257) );
  XNOR U30839 ( .A(n22901), .B(n22905), .Z(n23258) );
  XNOR U30840 ( .A(n22896), .B(n22900), .Z(n23259) );
  XNOR U30841 ( .A(n22891), .B(n22895), .Z(n23260) );
  XNOR U30842 ( .A(n22886), .B(n22890), .Z(n23261) );
  XNOR U30843 ( .A(n22881), .B(n22885), .Z(n23262) );
  XNOR U30844 ( .A(n22876), .B(n22880), .Z(n23263) );
  XNOR U30845 ( .A(n22871), .B(n22875), .Z(n23264) );
  XNOR U30846 ( .A(n23265), .B(n23266), .Z(n22871) );
  XNOR U30847 ( .A(n22866), .B(n22870), .Z(n23266) );
  XNOR U30848 ( .A(n22861), .B(n22865), .Z(n23267) );
  XNOR U30849 ( .A(n22856), .B(n22860), .Z(n23268) );
  XNOR U30850 ( .A(n22851), .B(n22855), .Z(n23269) );
  XNOR U30851 ( .A(n22846), .B(n22850), .Z(n23270) );
  XNOR U30852 ( .A(n22841), .B(n22845), .Z(n23271) );
  XNOR U30853 ( .A(n22836), .B(n22840), .Z(n23272) );
  XNOR U30854 ( .A(n22831), .B(n22835), .Z(n23273) );
  XNOR U30855 ( .A(n22826), .B(n22830), .Z(n23274) );
  XNOR U30856 ( .A(n22821), .B(n22825), .Z(n23275) );
  XNOR U30857 ( .A(n22816), .B(n22820), .Z(n23276) );
  XNOR U30858 ( .A(n22811), .B(n22815), .Z(n23277) );
  XNOR U30859 ( .A(n22806), .B(n22810), .Z(n23278) );
  XNOR U30860 ( .A(n22801), .B(n22805), .Z(n23279) );
  XNOR U30861 ( .A(n22796), .B(n22800), .Z(n23280) );
  XNOR U30862 ( .A(n22791), .B(n22795), .Z(n23281) );
  XNOR U30863 ( .A(n22786), .B(n22790), .Z(n23282) );
  XNOR U30864 ( .A(n22781), .B(n22785), .Z(n23283) );
  XNOR U30865 ( .A(n22776), .B(n22780), .Z(n23284) );
  XNOR U30866 ( .A(n22771), .B(n22775), .Z(n23285) );
  XNOR U30867 ( .A(n22766), .B(n22770), .Z(n23286) );
  XNOR U30868 ( .A(n22761), .B(n22765), .Z(n23287) );
  XNOR U30869 ( .A(n22756), .B(n22760), .Z(n23288) );
  XNOR U30870 ( .A(n22751), .B(n22755), .Z(n23289) );
  XNOR U30871 ( .A(n23290), .B(n22750), .Z(n22751) );
  AND U30872 ( .A(a[0]), .B(b[91]), .Z(n23290) );
  XOR U30873 ( .A(n23291), .B(n22750), .Z(n22752) );
  XNOR U30874 ( .A(n23292), .B(n23293), .Z(n22750) );
  ANDN U30875 ( .B(n23294), .A(n23295), .Z(n23292) );
  AND U30876 ( .A(a[1]), .B(b[90]), .Z(n23291) );
  XOR U30877 ( .A(n23297), .B(n23298), .Z(n22755) );
  ANDN U30878 ( .B(n23299), .A(n23300), .Z(n23297) );
  AND U30879 ( .A(a[2]), .B(b[89]), .Z(n23296) );
  XOR U30880 ( .A(n23302), .B(n23303), .Z(n22760) );
  ANDN U30881 ( .B(n23304), .A(n23305), .Z(n23302) );
  AND U30882 ( .A(a[3]), .B(b[88]), .Z(n23301) );
  XOR U30883 ( .A(n23307), .B(n23308), .Z(n22765) );
  ANDN U30884 ( .B(n23309), .A(n23310), .Z(n23307) );
  AND U30885 ( .A(a[4]), .B(b[87]), .Z(n23306) );
  XOR U30886 ( .A(n23312), .B(n23313), .Z(n22770) );
  ANDN U30887 ( .B(n23314), .A(n23315), .Z(n23312) );
  AND U30888 ( .A(a[5]), .B(b[86]), .Z(n23311) );
  XOR U30889 ( .A(n23317), .B(n23318), .Z(n22775) );
  ANDN U30890 ( .B(n23319), .A(n23320), .Z(n23317) );
  AND U30891 ( .A(a[6]), .B(b[85]), .Z(n23316) );
  XOR U30892 ( .A(n23322), .B(n23323), .Z(n22780) );
  ANDN U30893 ( .B(n23324), .A(n23325), .Z(n23322) );
  AND U30894 ( .A(a[7]), .B(b[84]), .Z(n23321) );
  XOR U30895 ( .A(n23327), .B(n23328), .Z(n22785) );
  ANDN U30896 ( .B(n23329), .A(n23330), .Z(n23327) );
  AND U30897 ( .A(a[8]), .B(b[83]), .Z(n23326) );
  XOR U30898 ( .A(n23332), .B(n23333), .Z(n22790) );
  ANDN U30899 ( .B(n23334), .A(n23335), .Z(n23332) );
  AND U30900 ( .A(a[9]), .B(b[82]), .Z(n23331) );
  XOR U30901 ( .A(n23337), .B(n23338), .Z(n22795) );
  ANDN U30902 ( .B(n23339), .A(n23340), .Z(n23337) );
  AND U30903 ( .A(a[10]), .B(b[81]), .Z(n23336) );
  XOR U30904 ( .A(n23342), .B(n23343), .Z(n22800) );
  ANDN U30905 ( .B(n23344), .A(n23345), .Z(n23342) );
  AND U30906 ( .A(a[11]), .B(b[80]), .Z(n23341) );
  XOR U30907 ( .A(n23347), .B(n23348), .Z(n22805) );
  ANDN U30908 ( .B(n23349), .A(n23350), .Z(n23347) );
  AND U30909 ( .A(a[12]), .B(b[79]), .Z(n23346) );
  XOR U30910 ( .A(n23352), .B(n23353), .Z(n22810) );
  ANDN U30911 ( .B(n23354), .A(n23355), .Z(n23352) );
  AND U30912 ( .A(a[13]), .B(b[78]), .Z(n23351) );
  XOR U30913 ( .A(n23357), .B(n23358), .Z(n22815) );
  ANDN U30914 ( .B(n23359), .A(n23360), .Z(n23357) );
  AND U30915 ( .A(a[14]), .B(b[77]), .Z(n23356) );
  XOR U30916 ( .A(n23362), .B(n23363), .Z(n22820) );
  ANDN U30917 ( .B(n23364), .A(n23365), .Z(n23362) );
  AND U30918 ( .A(a[15]), .B(b[76]), .Z(n23361) );
  XOR U30919 ( .A(n23367), .B(n23368), .Z(n22825) );
  ANDN U30920 ( .B(n23369), .A(n23370), .Z(n23367) );
  AND U30921 ( .A(a[16]), .B(b[75]), .Z(n23366) );
  XOR U30922 ( .A(n23372), .B(n23373), .Z(n22830) );
  ANDN U30923 ( .B(n23374), .A(n23375), .Z(n23372) );
  AND U30924 ( .A(a[17]), .B(b[74]), .Z(n23371) );
  XOR U30925 ( .A(n23377), .B(n23378), .Z(n22835) );
  ANDN U30926 ( .B(n23379), .A(n23380), .Z(n23377) );
  AND U30927 ( .A(a[18]), .B(b[73]), .Z(n23376) );
  XOR U30928 ( .A(n23382), .B(n23383), .Z(n22840) );
  ANDN U30929 ( .B(n23384), .A(n23385), .Z(n23382) );
  AND U30930 ( .A(a[19]), .B(b[72]), .Z(n23381) );
  XOR U30931 ( .A(n23387), .B(n23388), .Z(n22845) );
  ANDN U30932 ( .B(n23389), .A(n23390), .Z(n23387) );
  AND U30933 ( .A(a[20]), .B(b[71]), .Z(n23386) );
  XOR U30934 ( .A(n23392), .B(n23393), .Z(n22850) );
  ANDN U30935 ( .B(n23394), .A(n23395), .Z(n23392) );
  AND U30936 ( .A(a[21]), .B(b[70]), .Z(n23391) );
  XOR U30937 ( .A(n23397), .B(n23398), .Z(n22855) );
  ANDN U30938 ( .B(n23399), .A(n23400), .Z(n23397) );
  AND U30939 ( .A(a[22]), .B(b[69]), .Z(n23396) );
  XOR U30940 ( .A(n23402), .B(n23403), .Z(n22860) );
  ANDN U30941 ( .B(n23404), .A(n23405), .Z(n23402) );
  AND U30942 ( .A(a[23]), .B(b[68]), .Z(n23401) );
  IV U30943 ( .A(n22867), .Z(n23265) );
  XOR U30944 ( .A(n23407), .B(n23408), .Z(n22865) );
  ANDN U30945 ( .B(n23409), .A(n23410), .Z(n23407) );
  AND U30946 ( .A(a[24]), .B(b[67]), .Z(n23406) );
  XOR U30947 ( .A(n23412), .B(n23413), .Z(n22870) );
  ANDN U30948 ( .B(n23414), .A(n23415), .Z(n23412) );
  AND U30949 ( .A(a[25]), .B(b[66]), .Z(n23411) );
  XOR U30950 ( .A(n23417), .B(n23418), .Z(n22875) );
  ANDN U30951 ( .B(n23419), .A(n23420), .Z(n23417) );
  AND U30952 ( .A(a[26]), .B(b[65]), .Z(n23416) );
  XOR U30953 ( .A(n23422), .B(n23423), .Z(n22880) );
  ANDN U30954 ( .B(n23424), .A(n23425), .Z(n23422) );
  AND U30955 ( .A(a[27]), .B(b[64]), .Z(n23421) );
  XOR U30956 ( .A(n23427), .B(n23428), .Z(n22885) );
  ANDN U30957 ( .B(n23429), .A(n23430), .Z(n23427) );
  AND U30958 ( .A(a[28]), .B(b[63]), .Z(n23426) );
  XOR U30959 ( .A(n23432), .B(n23433), .Z(n22890) );
  ANDN U30960 ( .B(n23434), .A(n23435), .Z(n23432) );
  AND U30961 ( .A(a[29]), .B(b[62]), .Z(n23431) );
  XOR U30962 ( .A(n23437), .B(n23438), .Z(n22895) );
  ANDN U30963 ( .B(n23439), .A(n23440), .Z(n23437) );
  AND U30964 ( .A(a[30]), .B(b[61]), .Z(n23436) );
  XOR U30965 ( .A(n23442), .B(n23443), .Z(n22900) );
  ANDN U30966 ( .B(n23444), .A(n23445), .Z(n23442) );
  AND U30967 ( .A(a[31]), .B(b[60]), .Z(n23441) );
  XOR U30968 ( .A(n23447), .B(n23448), .Z(n22905) );
  ANDN U30969 ( .B(n23449), .A(n23450), .Z(n23447) );
  AND U30970 ( .A(a[32]), .B(b[59]), .Z(n23446) );
  XOR U30971 ( .A(n23452), .B(n23453), .Z(n22910) );
  ANDN U30972 ( .B(n23454), .A(n23455), .Z(n23452) );
  AND U30973 ( .A(a[33]), .B(b[58]), .Z(n23451) );
  XOR U30974 ( .A(n23457), .B(n23458), .Z(n22915) );
  ANDN U30975 ( .B(n23459), .A(n23460), .Z(n23457) );
  AND U30976 ( .A(a[34]), .B(b[57]), .Z(n23456) );
  XOR U30977 ( .A(n23462), .B(n23463), .Z(n22920) );
  ANDN U30978 ( .B(n23464), .A(n23465), .Z(n23462) );
  AND U30979 ( .A(a[35]), .B(b[56]), .Z(n23461) );
  XOR U30980 ( .A(n23467), .B(n23468), .Z(n22925) );
  ANDN U30981 ( .B(n23469), .A(n23470), .Z(n23467) );
  AND U30982 ( .A(a[36]), .B(b[55]), .Z(n23466) );
  XOR U30983 ( .A(n23472), .B(n23473), .Z(n22930) );
  ANDN U30984 ( .B(n23474), .A(n23475), .Z(n23472) );
  AND U30985 ( .A(a[37]), .B(b[54]), .Z(n23471) );
  XOR U30986 ( .A(n23477), .B(n23478), .Z(n22935) );
  ANDN U30987 ( .B(n23479), .A(n23480), .Z(n23477) );
  AND U30988 ( .A(a[38]), .B(b[53]), .Z(n23476) );
  XOR U30989 ( .A(n23482), .B(n23483), .Z(n22940) );
  ANDN U30990 ( .B(n23484), .A(n23485), .Z(n23482) );
  AND U30991 ( .A(a[39]), .B(b[52]), .Z(n23481) );
  XOR U30992 ( .A(n23487), .B(n23488), .Z(n22945) );
  ANDN U30993 ( .B(n23489), .A(n23490), .Z(n23487) );
  AND U30994 ( .A(a[40]), .B(b[51]), .Z(n23486) );
  XOR U30995 ( .A(n23492), .B(n23493), .Z(n22950) );
  ANDN U30996 ( .B(n23494), .A(n23495), .Z(n23492) );
  AND U30997 ( .A(a[41]), .B(b[50]), .Z(n23491) );
  XOR U30998 ( .A(n23497), .B(n23498), .Z(n22955) );
  ANDN U30999 ( .B(n23499), .A(n23500), .Z(n23497) );
  AND U31000 ( .A(a[42]), .B(b[49]), .Z(n23496) );
  XOR U31001 ( .A(n23502), .B(n23503), .Z(n22960) );
  ANDN U31002 ( .B(n23504), .A(n23505), .Z(n23502) );
  AND U31003 ( .A(a[43]), .B(b[48]), .Z(n23501) );
  XOR U31004 ( .A(n23507), .B(n23508), .Z(n22965) );
  ANDN U31005 ( .B(n23509), .A(n23510), .Z(n23507) );
  AND U31006 ( .A(a[44]), .B(b[47]), .Z(n23506) );
  XOR U31007 ( .A(n23512), .B(n23513), .Z(n22970) );
  ANDN U31008 ( .B(n23514), .A(n23515), .Z(n23512) );
  AND U31009 ( .A(a[45]), .B(b[46]), .Z(n23511) );
  XOR U31010 ( .A(n23517), .B(n23518), .Z(n22975) );
  ANDN U31011 ( .B(n23519), .A(n23520), .Z(n23517) );
  AND U31012 ( .A(a[46]), .B(b[45]), .Z(n23516) );
  XOR U31013 ( .A(n23522), .B(n23523), .Z(n22980) );
  ANDN U31014 ( .B(n23524), .A(n23525), .Z(n23522) );
  AND U31015 ( .A(a[47]), .B(b[44]), .Z(n23521) );
  XOR U31016 ( .A(n23527), .B(n23528), .Z(n22985) );
  ANDN U31017 ( .B(n23529), .A(n23530), .Z(n23527) );
  AND U31018 ( .A(a[48]), .B(b[43]), .Z(n23526) );
  XOR U31019 ( .A(n23532), .B(n23533), .Z(n22990) );
  ANDN U31020 ( .B(n23534), .A(n23535), .Z(n23532) );
  AND U31021 ( .A(a[49]), .B(b[42]), .Z(n23531) );
  XOR U31022 ( .A(n23537), .B(n23538), .Z(n22995) );
  ANDN U31023 ( .B(n23539), .A(n23540), .Z(n23537) );
  AND U31024 ( .A(a[50]), .B(b[41]), .Z(n23536) );
  XOR U31025 ( .A(n23542), .B(n23543), .Z(n23000) );
  ANDN U31026 ( .B(n23544), .A(n23545), .Z(n23542) );
  AND U31027 ( .A(a[51]), .B(b[40]), .Z(n23541) );
  XOR U31028 ( .A(n23547), .B(n23548), .Z(n23005) );
  ANDN U31029 ( .B(n23549), .A(n23550), .Z(n23547) );
  AND U31030 ( .A(a[52]), .B(b[39]), .Z(n23546) );
  XOR U31031 ( .A(n23552), .B(n23553), .Z(n23010) );
  ANDN U31032 ( .B(n23554), .A(n23555), .Z(n23552) );
  AND U31033 ( .A(a[53]), .B(b[38]), .Z(n23551) );
  XOR U31034 ( .A(n23557), .B(n23558), .Z(n23015) );
  ANDN U31035 ( .B(n23559), .A(n23560), .Z(n23557) );
  AND U31036 ( .A(a[54]), .B(b[37]), .Z(n23556) );
  XOR U31037 ( .A(n23562), .B(n23563), .Z(n23020) );
  ANDN U31038 ( .B(n23564), .A(n23565), .Z(n23562) );
  AND U31039 ( .A(a[55]), .B(b[36]), .Z(n23561) );
  XOR U31040 ( .A(n23567), .B(n23568), .Z(n23025) );
  ANDN U31041 ( .B(n23569), .A(n23570), .Z(n23567) );
  AND U31042 ( .A(a[56]), .B(b[35]), .Z(n23566) );
  XOR U31043 ( .A(n23572), .B(n23573), .Z(n23030) );
  ANDN U31044 ( .B(n23574), .A(n23575), .Z(n23572) );
  AND U31045 ( .A(a[57]), .B(b[34]), .Z(n23571) );
  XOR U31046 ( .A(n23577), .B(n23578), .Z(n23035) );
  ANDN U31047 ( .B(n23579), .A(n23580), .Z(n23577) );
  AND U31048 ( .A(a[58]), .B(b[33]), .Z(n23576) );
  XOR U31049 ( .A(n23582), .B(n23583), .Z(n23040) );
  ANDN U31050 ( .B(n23584), .A(n23585), .Z(n23582) );
  AND U31051 ( .A(a[59]), .B(b[32]), .Z(n23581) );
  XOR U31052 ( .A(n23587), .B(n23588), .Z(n23045) );
  ANDN U31053 ( .B(n23589), .A(n23590), .Z(n23587) );
  AND U31054 ( .A(a[60]), .B(b[31]), .Z(n23586) );
  XOR U31055 ( .A(n23592), .B(n23593), .Z(n23050) );
  ANDN U31056 ( .B(n23594), .A(n23595), .Z(n23592) );
  AND U31057 ( .A(a[61]), .B(b[30]), .Z(n23591) );
  XOR U31058 ( .A(n23597), .B(n23598), .Z(n23055) );
  ANDN U31059 ( .B(n23599), .A(n23600), .Z(n23597) );
  AND U31060 ( .A(a[62]), .B(b[29]), .Z(n23596) );
  XOR U31061 ( .A(n23602), .B(n23603), .Z(n23060) );
  ANDN U31062 ( .B(n23604), .A(n23605), .Z(n23602) );
  AND U31063 ( .A(a[63]), .B(b[28]), .Z(n23601) );
  XOR U31064 ( .A(n23607), .B(n23608), .Z(n23065) );
  ANDN U31065 ( .B(n23609), .A(n23610), .Z(n23607) );
  AND U31066 ( .A(a[64]), .B(b[27]), .Z(n23606) );
  XOR U31067 ( .A(n23612), .B(n23613), .Z(n23070) );
  ANDN U31068 ( .B(n23614), .A(n23615), .Z(n23612) );
  AND U31069 ( .A(a[65]), .B(b[26]), .Z(n23611) );
  XOR U31070 ( .A(n23617), .B(n23618), .Z(n23075) );
  ANDN U31071 ( .B(n23619), .A(n23620), .Z(n23617) );
  AND U31072 ( .A(a[66]), .B(b[25]), .Z(n23616) );
  XOR U31073 ( .A(n23622), .B(n23623), .Z(n23080) );
  ANDN U31074 ( .B(n23624), .A(n23625), .Z(n23622) );
  AND U31075 ( .A(a[67]), .B(b[24]), .Z(n23621) );
  XOR U31076 ( .A(n23627), .B(n23628), .Z(n23085) );
  ANDN U31077 ( .B(n23629), .A(n23630), .Z(n23627) );
  AND U31078 ( .A(a[68]), .B(b[23]), .Z(n23626) );
  XOR U31079 ( .A(n23632), .B(n23633), .Z(n23090) );
  ANDN U31080 ( .B(n23634), .A(n23635), .Z(n23632) );
  AND U31081 ( .A(a[69]), .B(b[22]), .Z(n23631) );
  XOR U31082 ( .A(n23637), .B(n23638), .Z(n23095) );
  ANDN U31083 ( .B(n23639), .A(n23640), .Z(n23637) );
  AND U31084 ( .A(a[70]), .B(b[21]), .Z(n23636) );
  XOR U31085 ( .A(n23642), .B(n23643), .Z(n23100) );
  ANDN U31086 ( .B(n23644), .A(n23645), .Z(n23642) );
  AND U31087 ( .A(a[71]), .B(b[20]), .Z(n23641) );
  XOR U31088 ( .A(n23647), .B(n23648), .Z(n23105) );
  ANDN U31089 ( .B(n23649), .A(n23650), .Z(n23647) );
  AND U31090 ( .A(a[72]), .B(b[19]), .Z(n23646) );
  XOR U31091 ( .A(n23652), .B(n23653), .Z(n23110) );
  ANDN U31092 ( .B(n23654), .A(n23655), .Z(n23652) );
  AND U31093 ( .A(a[73]), .B(b[18]), .Z(n23651) );
  XOR U31094 ( .A(n23657), .B(n23658), .Z(n23115) );
  ANDN U31095 ( .B(n23659), .A(n23660), .Z(n23657) );
  AND U31096 ( .A(a[74]), .B(b[17]), .Z(n23656) );
  XOR U31097 ( .A(n23662), .B(n23663), .Z(n23120) );
  ANDN U31098 ( .B(n23664), .A(n23665), .Z(n23662) );
  AND U31099 ( .A(a[75]), .B(b[16]), .Z(n23661) );
  XOR U31100 ( .A(n23667), .B(n23668), .Z(n23125) );
  ANDN U31101 ( .B(n23669), .A(n23670), .Z(n23667) );
  AND U31102 ( .A(a[76]), .B(b[15]), .Z(n23666) );
  XOR U31103 ( .A(n23672), .B(n23673), .Z(n23130) );
  ANDN U31104 ( .B(n23674), .A(n23675), .Z(n23672) );
  AND U31105 ( .A(a[77]), .B(b[14]), .Z(n23671) );
  XOR U31106 ( .A(n23677), .B(n23678), .Z(n23135) );
  ANDN U31107 ( .B(n23679), .A(n23680), .Z(n23677) );
  AND U31108 ( .A(a[78]), .B(b[13]), .Z(n23676) );
  XOR U31109 ( .A(n23682), .B(n23683), .Z(n23140) );
  ANDN U31110 ( .B(n23684), .A(n23685), .Z(n23682) );
  AND U31111 ( .A(a[79]), .B(b[12]), .Z(n23681) );
  XOR U31112 ( .A(n23687), .B(n23688), .Z(n23145) );
  ANDN U31113 ( .B(n23689), .A(n23690), .Z(n23687) );
  AND U31114 ( .A(a[80]), .B(b[11]), .Z(n23686) );
  XOR U31115 ( .A(n23692), .B(n23693), .Z(n23150) );
  ANDN U31116 ( .B(n23694), .A(n23695), .Z(n23692) );
  AND U31117 ( .A(a[81]), .B(b[10]), .Z(n23691) );
  XOR U31118 ( .A(n23697), .B(n23698), .Z(n23155) );
  ANDN U31119 ( .B(n23699), .A(n23700), .Z(n23697) );
  AND U31120 ( .A(b[9]), .B(a[82]), .Z(n23696) );
  XOR U31121 ( .A(n23702), .B(n23703), .Z(n23160) );
  ANDN U31122 ( .B(n23704), .A(n23705), .Z(n23702) );
  AND U31123 ( .A(b[8]), .B(a[83]), .Z(n23701) );
  XOR U31124 ( .A(n23707), .B(n23708), .Z(n23165) );
  ANDN U31125 ( .B(n23709), .A(n23710), .Z(n23707) );
  AND U31126 ( .A(b[7]), .B(a[84]), .Z(n23706) );
  XOR U31127 ( .A(n23712), .B(n23713), .Z(n23170) );
  ANDN U31128 ( .B(n23714), .A(n23715), .Z(n23712) );
  AND U31129 ( .A(b[6]), .B(a[85]), .Z(n23711) );
  XOR U31130 ( .A(n23717), .B(n23718), .Z(n23175) );
  ANDN U31131 ( .B(n23719), .A(n23720), .Z(n23717) );
  AND U31132 ( .A(b[5]), .B(a[86]), .Z(n23716) );
  XOR U31133 ( .A(n23722), .B(n23723), .Z(n23180) );
  ANDN U31134 ( .B(n23724), .A(n23725), .Z(n23722) );
  AND U31135 ( .A(b[4]), .B(a[87]), .Z(n23721) );
  XOR U31136 ( .A(n23727), .B(n23728), .Z(n23185) );
  ANDN U31137 ( .B(n23197), .A(n23198), .Z(n23727) );
  AND U31138 ( .A(b[2]), .B(a[88]), .Z(n23729) );
  XNOR U31139 ( .A(n23724), .B(n23728), .Z(n23730) );
  XOR U31140 ( .A(n23731), .B(n23732), .Z(n23728) );
  OR U31141 ( .A(n23200), .B(n23201), .Z(n23732) );
  XNOR U31142 ( .A(n23734), .B(n23735), .Z(n23733) );
  XOR U31143 ( .A(n23734), .B(n23737), .Z(n23200) );
  NAND U31144 ( .A(b[1]), .B(a[88]), .Z(n23737) );
  IV U31145 ( .A(n23731), .Z(n23734) );
  NANDN U31146 ( .A(n27), .B(n28), .Z(n23731) );
  XOR U31147 ( .A(n23738), .B(n23739), .Z(n28) );
  NAND U31148 ( .A(a[88]), .B(b[0]), .Z(n27) );
  XNOR U31149 ( .A(n23719), .B(n23723), .Z(n23740) );
  XNOR U31150 ( .A(n23714), .B(n23718), .Z(n23741) );
  XNOR U31151 ( .A(n23709), .B(n23713), .Z(n23742) );
  XNOR U31152 ( .A(n23704), .B(n23708), .Z(n23743) );
  XNOR U31153 ( .A(n23699), .B(n23703), .Z(n23744) );
  XNOR U31154 ( .A(n23694), .B(n23698), .Z(n23745) );
  XNOR U31155 ( .A(n23689), .B(n23693), .Z(n23746) );
  XNOR U31156 ( .A(n23684), .B(n23688), .Z(n23747) );
  XNOR U31157 ( .A(n23679), .B(n23683), .Z(n23748) );
  XNOR U31158 ( .A(n23674), .B(n23678), .Z(n23749) );
  XNOR U31159 ( .A(n23669), .B(n23673), .Z(n23750) );
  XNOR U31160 ( .A(n23664), .B(n23668), .Z(n23751) );
  XNOR U31161 ( .A(n23659), .B(n23663), .Z(n23752) );
  XNOR U31162 ( .A(n23654), .B(n23658), .Z(n23753) );
  XNOR U31163 ( .A(n23649), .B(n23653), .Z(n23754) );
  XNOR U31164 ( .A(n23644), .B(n23648), .Z(n23755) );
  XNOR U31165 ( .A(n23639), .B(n23643), .Z(n23756) );
  XNOR U31166 ( .A(n23634), .B(n23638), .Z(n23757) );
  XNOR U31167 ( .A(n23629), .B(n23633), .Z(n23758) );
  XNOR U31168 ( .A(n23624), .B(n23628), .Z(n23759) );
  XNOR U31169 ( .A(n23619), .B(n23623), .Z(n23760) );
  XNOR U31170 ( .A(n23614), .B(n23618), .Z(n23761) );
  XNOR U31171 ( .A(n23609), .B(n23613), .Z(n23762) );
  XNOR U31172 ( .A(n23604), .B(n23608), .Z(n23763) );
  XNOR U31173 ( .A(n23599), .B(n23603), .Z(n23764) );
  XNOR U31174 ( .A(n23594), .B(n23598), .Z(n23765) );
  XNOR U31175 ( .A(n23589), .B(n23593), .Z(n23766) );
  XNOR U31176 ( .A(n23584), .B(n23588), .Z(n23767) );
  XNOR U31177 ( .A(n23579), .B(n23583), .Z(n23768) );
  XNOR U31178 ( .A(n23574), .B(n23578), .Z(n23769) );
  XNOR U31179 ( .A(n23569), .B(n23573), .Z(n23770) );
  XNOR U31180 ( .A(n23564), .B(n23568), .Z(n23771) );
  XNOR U31181 ( .A(n23559), .B(n23563), .Z(n23772) );
  XNOR U31182 ( .A(n23554), .B(n23558), .Z(n23773) );
  XNOR U31183 ( .A(n23549), .B(n23553), .Z(n23774) );
  XNOR U31184 ( .A(n23544), .B(n23548), .Z(n23775) );
  XNOR U31185 ( .A(n23539), .B(n23543), .Z(n23776) );
  XNOR U31186 ( .A(n23534), .B(n23538), .Z(n23777) );
  XNOR U31187 ( .A(n23529), .B(n23533), .Z(n23778) );
  XNOR U31188 ( .A(n23524), .B(n23528), .Z(n23779) );
  XNOR U31189 ( .A(n23519), .B(n23523), .Z(n23780) );
  XNOR U31190 ( .A(n23514), .B(n23518), .Z(n23781) );
  XNOR U31191 ( .A(n23509), .B(n23513), .Z(n23782) );
  XNOR U31192 ( .A(n23504), .B(n23508), .Z(n23783) );
  XNOR U31193 ( .A(n23499), .B(n23503), .Z(n23784) );
  XNOR U31194 ( .A(n23494), .B(n23498), .Z(n23785) );
  XNOR U31195 ( .A(n23489), .B(n23493), .Z(n23786) );
  XNOR U31196 ( .A(n23484), .B(n23488), .Z(n23787) );
  XNOR U31197 ( .A(n23479), .B(n23483), .Z(n23788) );
  XNOR U31198 ( .A(n23474), .B(n23478), .Z(n23789) );
  XNOR U31199 ( .A(n23469), .B(n23473), .Z(n23790) );
  XNOR U31200 ( .A(n23464), .B(n23468), .Z(n23791) );
  XNOR U31201 ( .A(n23459), .B(n23463), .Z(n23792) );
  XNOR U31202 ( .A(n23454), .B(n23458), .Z(n23793) );
  XNOR U31203 ( .A(n23449), .B(n23453), .Z(n23794) );
  XNOR U31204 ( .A(n23444), .B(n23448), .Z(n23795) );
  XNOR U31205 ( .A(n23439), .B(n23443), .Z(n23796) );
  XNOR U31206 ( .A(n23434), .B(n23438), .Z(n23797) );
  XNOR U31207 ( .A(n23429), .B(n23433), .Z(n23798) );
  XNOR U31208 ( .A(n23424), .B(n23428), .Z(n23799) );
  XNOR U31209 ( .A(n23419), .B(n23423), .Z(n23800) );
  XNOR U31210 ( .A(n23414), .B(n23418), .Z(n23801) );
  XNOR U31211 ( .A(n23409), .B(n23413), .Z(n23802) );
  XNOR U31212 ( .A(n23404), .B(n23408), .Z(n23803) );
  XNOR U31213 ( .A(n23399), .B(n23403), .Z(n23804) );
  XNOR U31214 ( .A(n23394), .B(n23398), .Z(n23805) );
  XNOR U31215 ( .A(n23389), .B(n23393), .Z(n23806) );
  XNOR U31216 ( .A(n23384), .B(n23388), .Z(n23807) );
  XNOR U31217 ( .A(n23379), .B(n23383), .Z(n23808) );
  XNOR U31218 ( .A(n23374), .B(n23378), .Z(n23809) );
  XNOR U31219 ( .A(n23369), .B(n23373), .Z(n23810) );
  XNOR U31220 ( .A(n23364), .B(n23368), .Z(n23811) );
  XNOR U31221 ( .A(n23359), .B(n23363), .Z(n23812) );
  XNOR U31222 ( .A(n23354), .B(n23358), .Z(n23813) );
  XNOR U31223 ( .A(n23349), .B(n23353), .Z(n23814) );
  XNOR U31224 ( .A(n23344), .B(n23348), .Z(n23815) );
  XNOR U31225 ( .A(n23339), .B(n23343), .Z(n23816) );
  XNOR U31226 ( .A(n23334), .B(n23338), .Z(n23817) );
  XNOR U31227 ( .A(n23329), .B(n23333), .Z(n23818) );
  XNOR U31228 ( .A(n23324), .B(n23328), .Z(n23819) );
  XNOR U31229 ( .A(n23319), .B(n23323), .Z(n23820) );
  XNOR U31230 ( .A(n23314), .B(n23318), .Z(n23821) );
  XNOR U31231 ( .A(n23309), .B(n23313), .Z(n23822) );
  XNOR U31232 ( .A(n23304), .B(n23308), .Z(n23823) );
  XNOR U31233 ( .A(n23299), .B(n23303), .Z(n23824) );
  XNOR U31234 ( .A(n23294), .B(n23298), .Z(n23825) );
  XOR U31235 ( .A(n23826), .B(n23293), .Z(n23294) );
  AND U31236 ( .A(a[0]), .B(b[90]), .Z(n23826) );
  XNOR U31237 ( .A(n23827), .B(n23293), .Z(n23295) );
  XNOR U31238 ( .A(n23828), .B(n23829), .Z(n23293) );
  ANDN U31239 ( .B(n23830), .A(n23831), .Z(n23828) );
  AND U31240 ( .A(a[1]), .B(b[89]), .Z(n23827) );
  XOR U31241 ( .A(n23833), .B(n23834), .Z(n23298) );
  ANDN U31242 ( .B(n23835), .A(n23836), .Z(n23833) );
  AND U31243 ( .A(a[2]), .B(b[88]), .Z(n23832) );
  XOR U31244 ( .A(n23838), .B(n23839), .Z(n23303) );
  ANDN U31245 ( .B(n23840), .A(n23841), .Z(n23838) );
  AND U31246 ( .A(a[3]), .B(b[87]), .Z(n23837) );
  XOR U31247 ( .A(n23843), .B(n23844), .Z(n23308) );
  ANDN U31248 ( .B(n23845), .A(n23846), .Z(n23843) );
  AND U31249 ( .A(a[4]), .B(b[86]), .Z(n23842) );
  XOR U31250 ( .A(n23848), .B(n23849), .Z(n23313) );
  ANDN U31251 ( .B(n23850), .A(n23851), .Z(n23848) );
  AND U31252 ( .A(a[5]), .B(b[85]), .Z(n23847) );
  XOR U31253 ( .A(n23853), .B(n23854), .Z(n23318) );
  ANDN U31254 ( .B(n23855), .A(n23856), .Z(n23853) );
  AND U31255 ( .A(a[6]), .B(b[84]), .Z(n23852) );
  XOR U31256 ( .A(n23858), .B(n23859), .Z(n23323) );
  ANDN U31257 ( .B(n23860), .A(n23861), .Z(n23858) );
  AND U31258 ( .A(a[7]), .B(b[83]), .Z(n23857) );
  XOR U31259 ( .A(n23863), .B(n23864), .Z(n23328) );
  ANDN U31260 ( .B(n23865), .A(n23866), .Z(n23863) );
  AND U31261 ( .A(a[8]), .B(b[82]), .Z(n23862) );
  XOR U31262 ( .A(n23868), .B(n23869), .Z(n23333) );
  ANDN U31263 ( .B(n23870), .A(n23871), .Z(n23868) );
  AND U31264 ( .A(a[9]), .B(b[81]), .Z(n23867) );
  XOR U31265 ( .A(n23873), .B(n23874), .Z(n23338) );
  ANDN U31266 ( .B(n23875), .A(n23876), .Z(n23873) );
  AND U31267 ( .A(a[10]), .B(b[80]), .Z(n23872) );
  XOR U31268 ( .A(n23878), .B(n23879), .Z(n23343) );
  ANDN U31269 ( .B(n23880), .A(n23881), .Z(n23878) );
  AND U31270 ( .A(a[11]), .B(b[79]), .Z(n23877) );
  XOR U31271 ( .A(n23883), .B(n23884), .Z(n23348) );
  ANDN U31272 ( .B(n23885), .A(n23886), .Z(n23883) );
  AND U31273 ( .A(a[12]), .B(b[78]), .Z(n23882) );
  XOR U31274 ( .A(n23888), .B(n23889), .Z(n23353) );
  ANDN U31275 ( .B(n23890), .A(n23891), .Z(n23888) );
  AND U31276 ( .A(a[13]), .B(b[77]), .Z(n23887) );
  XOR U31277 ( .A(n23893), .B(n23894), .Z(n23358) );
  ANDN U31278 ( .B(n23895), .A(n23896), .Z(n23893) );
  AND U31279 ( .A(a[14]), .B(b[76]), .Z(n23892) );
  XOR U31280 ( .A(n23898), .B(n23899), .Z(n23363) );
  ANDN U31281 ( .B(n23900), .A(n23901), .Z(n23898) );
  AND U31282 ( .A(a[15]), .B(b[75]), .Z(n23897) );
  XOR U31283 ( .A(n23903), .B(n23904), .Z(n23368) );
  ANDN U31284 ( .B(n23905), .A(n23906), .Z(n23903) );
  AND U31285 ( .A(a[16]), .B(b[74]), .Z(n23902) );
  XOR U31286 ( .A(n23908), .B(n23909), .Z(n23373) );
  ANDN U31287 ( .B(n23910), .A(n23911), .Z(n23908) );
  AND U31288 ( .A(a[17]), .B(b[73]), .Z(n23907) );
  XOR U31289 ( .A(n23913), .B(n23914), .Z(n23378) );
  ANDN U31290 ( .B(n23915), .A(n23916), .Z(n23913) );
  AND U31291 ( .A(a[18]), .B(b[72]), .Z(n23912) );
  XOR U31292 ( .A(n23918), .B(n23919), .Z(n23383) );
  ANDN U31293 ( .B(n23920), .A(n23921), .Z(n23918) );
  AND U31294 ( .A(a[19]), .B(b[71]), .Z(n23917) );
  XOR U31295 ( .A(n23923), .B(n23924), .Z(n23388) );
  ANDN U31296 ( .B(n23925), .A(n23926), .Z(n23923) );
  AND U31297 ( .A(a[20]), .B(b[70]), .Z(n23922) );
  XOR U31298 ( .A(n23928), .B(n23929), .Z(n23393) );
  ANDN U31299 ( .B(n23930), .A(n23931), .Z(n23928) );
  AND U31300 ( .A(a[21]), .B(b[69]), .Z(n23927) );
  XOR U31301 ( .A(n23933), .B(n23934), .Z(n23398) );
  ANDN U31302 ( .B(n23935), .A(n23936), .Z(n23933) );
  AND U31303 ( .A(a[22]), .B(b[68]), .Z(n23932) );
  XOR U31304 ( .A(n23938), .B(n23939), .Z(n23403) );
  ANDN U31305 ( .B(n23940), .A(n23941), .Z(n23938) );
  AND U31306 ( .A(a[23]), .B(b[67]), .Z(n23937) );
  XOR U31307 ( .A(n23943), .B(n23944), .Z(n23408) );
  ANDN U31308 ( .B(n23945), .A(n23946), .Z(n23943) );
  AND U31309 ( .A(a[24]), .B(b[66]), .Z(n23942) );
  XOR U31310 ( .A(n23948), .B(n23949), .Z(n23413) );
  ANDN U31311 ( .B(n23950), .A(n23951), .Z(n23948) );
  AND U31312 ( .A(a[25]), .B(b[65]), .Z(n23947) );
  XOR U31313 ( .A(n23953), .B(n23954), .Z(n23418) );
  ANDN U31314 ( .B(n23955), .A(n23956), .Z(n23953) );
  AND U31315 ( .A(a[26]), .B(b[64]), .Z(n23952) );
  XOR U31316 ( .A(n23958), .B(n23959), .Z(n23423) );
  ANDN U31317 ( .B(n23960), .A(n23961), .Z(n23958) );
  AND U31318 ( .A(a[27]), .B(b[63]), .Z(n23957) );
  XOR U31319 ( .A(n23963), .B(n23964), .Z(n23428) );
  ANDN U31320 ( .B(n23965), .A(n23966), .Z(n23963) );
  AND U31321 ( .A(a[28]), .B(b[62]), .Z(n23962) );
  XOR U31322 ( .A(n23968), .B(n23969), .Z(n23433) );
  ANDN U31323 ( .B(n23970), .A(n23971), .Z(n23968) );
  AND U31324 ( .A(a[29]), .B(b[61]), .Z(n23967) );
  XOR U31325 ( .A(n23973), .B(n23974), .Z(n23438) );
  ANDN U31326 ( .B(n23975), .A(n23976), .Z(n23973) );
  AND U31327 ( .A(a[30]), .B(b[60]), .Z(n23972) );
  XOR U31328 ( .A(n23978), .B(n23979), .Z(n23443) );
  ANDN U31329 ( .B(n23980), .A(n23981), .Z(n23978) );
  AND U31330 ( .A(a[31]), .B(b[59]), .Z(n23977) );
  XOR U31331 ( .A(n23983), .B(n23984), .Z(n23448) );
  ANDN U31332 ( .B(n23985), .A(n23986), .Z(n23983) );
  AND U31333 ( .A(a[32]), .B(b[58]), .Z(n23982) );
  XOR U31334 ( .A(n23988), .B(n23989), .Z(n23453) );
  ANDN U31335 ( .B(n23990), .A(n23991), .Z(n23988) );
  AND U31336 ( .A(a[33]), .B(b[57]), .Z(n23987) );
  XOR U31337 ( .A(n23993), .B(n23994), .Z(n23458) );
  ANDN U31338 ( .B(n23995), .A(n23996), .Z(n23993) );
  AND U31339 ( .A(a[34]), .B(b[56]), .Z(n23992) );
  XOR U31340 ( .A(n23998), .B(n23999), .Z(n23463) );
  ANDN U31341 ( .B(n24000), .A(n24001), .Z(n23998) );
  AND U31342 ( .A(a[35]), .B(b[55]), .Z(n23997) );
  XOR U31343 ( .A(n24003), .B(n24004), .Z(n23468) );
  ANDN U31344 ( .B(n24005), .A(n24006), .Z(n24003) );
  AND U31345 ( .A(a[36]), .B(b[54]), .Z(n24002) );
  XOR U31346 ( .A(n24008), .B(n24009), .Z(n23473) );
  ANDN U31347 ( .B(n24010), .A(n24011), .Z(n24008) );
  AND U31348 ( .A(a[37]), .B(b[53]), .Z(n24007) );
  XOR U31349 ( .A(n24013), .B(n24014), .Z(n23478) );
  ANDN U31350 ( .B(n24015), .A(n24016), .Z(n24013) );
  AND U31351 ( .A(a[38]), .B(b[52]), .Z(n24012) );
  XOR U31352 ( .A(n24018), .B(n24019), .Z(n23483) );
  ANDN U31353 ( .B(n24020), .A(n24021), .Z(n24018) );
  AND U31354 ( .A(a[39]), .B(b[51]), .Z(n24017) );
  XOR U31355 ( .A(n24023), .B(n24024), .Z(n23488) );
  ANDN U31356 ( .B(n24025), .A(n24026), .Z(n24023) );
  AND U31357 ( .A(a[40]), .B(b[50]), .Z(n24022) );
  XOR U31358 ( .A(n24028), .B(n24029), .Z(n23493) );
  ANDN U31359 ( .B(n24030), .A(n24031), .Z(n24028) );
  AND U31360 ( .A(a[41]), .B(b[49]), .Z(n24027) );
  XOR U31361 ( .A(n24033), .B(n24034), .Z(n23498) );
  ANDN U31362 ( .B(n24035), .A(n24036), .Z(n24033) );
  AND U31363 ( .A(a[42]), .B(b[48]), .Z(n24032) );
  XOR U31364 ( .A(n24038), .B(n24039), .Z(n23503) );
  ANDN U31365 ( .B(n24040), .A(n24041), .Z(n24038) );
  AND U31366 ( .A(a[43]), .B(b[47]), .Z(n24037) );
  XOR U31367 ( .A(n24043), .B(n24044), .Z(n23508) );
  ANDN U31368 ( .B(n24045), .A(n24046), .Z(n24043) );
  AND U31369 ( .A(a[44]), .B(b[46]), .Z(n24042) );
  XOR U31370 ( .A(n24048), .B(n24049), .Z(n23513) );
  ANDN U31371 ( .B(n24050), .A(n24051), .Z(n24048) );
  AND U31372 ( .A(a[45]), .B(b[45]), .Z(n24047) );
  XOR U31373 ( .A(n24053), .B(n24054), .Z(n23518) );
  ANDN U31374 ( .B(n24055), .A(n24056), .Z(n24053) );
  AND U31375 ( .A(a[46]), .B(b[44]), .Z(n24052) );
  XOR U31376 ( .A(n24058), .B(n24059), .Z(n23523) );
  ANDN U31377 ( .B(n24060), .A(n24061), .Z(n24058) );
  AND U31378 ( .A(a[47]), .B(b[43]), .Z(n24057) );
  XOR U31379 ( .A(n24063), .B(n24064), .Z(n23528) );
  ANDN U31380 ( .B(n24065), .A(n24066), .Z(n24063) );
  AND U31381 ( .A(a[48]), .B(b[42]), .Z(n24062) );
  XOR U31382 ( .A(n24068), .B(n24069), .Z(n23533) );
  ANDN U31383 ( .B(n24070), .A(n24071), .Z(n24068) );
  AND U31384 ( .A(a[49]), .B(b[41]), .Z(n24067) );
  XOR U31385 ( .A(n24073), .B(n24074), .Z(n23538) );
  ANDN U31386 ( .B(n24075), .A(n24076), .Z(n24073) );
  AND U31387 ( .A(a[50]), .B(b[40]), .Z(n24072) );
  XOR U31388 ( .A(n24078), .B(n24079), .Z(n23543) );
  ANDN U31389 ( .B(n24080), .A(n24081), .Z(n24078) );
  AND U31390 ( .A(a[51]), .B(b[39]), .Z(n24077) );
  XOR U31391 ( .A(n24083), .B(n24084), .Z(n23548) );
  ANDN U31392 ( .B(n24085), .A(n24086), .Z(n24083) );
  AND U31393 ( .A(a[52]), .B(b[38]), .Z(n24082) );
  XOR U31394 ( .A(n24088), .B(n24089), .Z(n23553) );
  ANDN U31395 ( .B(n24090), .A(n24091), .Z(n24088) );
  AND U31396 ( .A(a[53]), .B(b[37]), .Z(n24087) );
  XOR U31397 ( .A(n24093), .B(n24094), .Z(n23558) );
  ANDN U31398 ( .B(n24095), .A(n24096), .Z(n24093) );
  AND U31399 ( .A(a[54]), .B(b[36]), .Z(n24092) );
  XOR U31400 ( .A(n24098), .B(n24099), .Z(n23563) );
  ANDN U31401 ( .B(n24100), .A(n24101), .Z(n24098) );
  AND U31402 ( .A(a[55]), .B(b[35]), .Z(n24097) );
  XOR U31403 ( .A(n24103), .B(n24104), .Z(n23568) );
  ANDN U31404 ( .B(n24105), .A(n24106), .Z(n24103) );
  AND U31405 ( .A(a[56]), .B(b[34]), .Z(n24102) );
  XOR U31406 ( .A(n24108), .B(n24109), .Z(n23573) );
  ANDN U31407 ( .B(n24110), .A(n24111), .Z(n24108) );
  AND U31408 ( .A(a[57]), .B(b[33]), .Z(n24107) );
  XOR U31409 ( .A(n24113), .B(n24114), .Z(n23578) );
  ANDN U31410 ( .B(n24115), .A(n24116), .Z(n24113) );
  AND U31411 ( .A(a[58]), .B(b[32]), .Z(n24112) );
  XOR U31412 ( .A(n24118), .B(n24119), .Z(n23583) );
  ANDN U31413 ( .B(n24120), .A(n24121), .Z(n24118) );
  AND U31414 ( .A(a[59]), .B(b[31]), .Z(n24117) );
  XOR U31415 ( .A(n24123), .B(n24124), .Z(n23588) );
  ANDN U31416 ( .B(n24125), .A(n24126), .Z(n24123) );
  AND U31417 ( .A(a[60]), .B(b[30]), .Z(n24122) );
  XOR U31418 ( .A(n24128), .B(n24129), .Z(n23593) );
  ANDN U31419 ( .B(n24130), .A(n24131), .Z(n24128) );
  AND U31420 ( .A(a[61]), .B(b[29]), .Z(n24127) );
  XOR U31421 ( .A(n24133), .B(n24134), .Z(n23598) );
  ANDN U31422 ( .B(n24135), .A(n24136), .Z(n24133) );
  AND U31423 ( .A(a[62]), .B(b[28]), .Z(n24132) );
  XOR U31424 ( .A(n24138), .B(n24139), .Z(n23603) );
  ANDN U31425 ( .B(n24140), .A(n24141), .Z(n24138) );
  AND U31426 ( .A(a[63]), .B(b[27]), .Z(n24137) );
  XOR U31427 ( .A(n24143), .B(n24144), .Z(n23608) );
  ANDN U31428 ( .B(n24145), .A(n24146), .Z(n24143) );
  AND U31429 ( .A(a[64]), .B(b[26]), .Z(n24142) );
  XOR U31430 ( .A(n24148), .B(n24149), .Z(n23613) );
  ANDN U31431 ( .B(n24150), .A(n24151), .Z(n24148) );
  AND U31432 ( .A(a[65]), .B(b[25]), .Z(n24147) );
  XOR U31433 ( .A(n24153), .B(n24154), .Z(n23618) );
  ANDN U31434 ( .B(n24155), .A(n24156), .Z(n24153) );
  AND U31435 ( .A(a[66]), .B(b[24]), .Z(n24152) );
  XOR U31436 ( .A(n24158), .B(n24159), .Z(n23623) );
  ANDN U31437 ( .B(n24160), .A(n24161), .Z(n24158) );
  AND U31438 ( .A(a[67]), .B(b[23]), .Z(n24157) );
  XOR U31439 ( .A(n24163), .B(n24164), .Z(n23628) );
  ANDN U31440 ( .B(n24165), .A(n24166), .Z(n24163) );
  AND U31441 ( .A(a[68]), .B(b[22]), .Z(n24162) );
  XOR U31442 ( .A(n24168), .B(n24169), .Z(n23633) );
  ANDN U31443 ( .B(n24170), .A(n24171), .Z(n24168) );
  AND U31444 ( .A(a[69]), .B(b[21]), .Z(n24167) );
  XOR U31445 ( .A(n24173), .B(n24174), .Z(n23638) );
  ANDN U31446 ( .B(n24175), .A(n24176), .Z(n24173) );
  AND U31447 ( .A(a[70]), .B(b[20]), .Z(n24172) );
  XOR U31448 ( .A(n24178), .B(n24179), .Z(n23643) );
  ANDN U31449 ( .B(n24180), .A(n24181), .Z(n24178) );
  AND U31450 ( .A(a[71]), .B(b[19]), .Z(n24177) );
  XOR U31451 ( .A(n24183), .B(n24184), .Z(n23648) );
  ANDN U31452 ( .B(n24185), .A(n24186), .Z(n24183) );
  AND U31453 ( .A(a[72]), .B(b[18]), .Z(n24182) );
  XOR U31454 ( .A(n24188), .B(n24189), .Z(n23653) );
  ANDN U31455 ( .B(n24190), .A(n24191), .Z(n24188) );
  AND U31456 ( .A(a[73]), .B(b[17]), .Z(n24187) );
  XOR U31457 ( .A(n24193), .B(n24194), .Z(n23658) );
  ANDN U31458 ( .B(n24195), .A(n24196), .Z(n24193) );
  AND U31459 ( .A(a[74]), .B(b[16]), .Z(n24192) );
  XOR U31460 ( .A(n24198), .B(n24199), .Z(n23663) );
  ANDN U31461 ( .B(n24200), .A(n24201), .Z(n24198) );
  AND U31462 ( .A(a[75]), .B(b[15]), .Z(n24197) );
  XOR U31463 ( .A(n24203), .B(n24204), .Z(n23668) );
  ANDN U31464 ( .B(n24205), .A(n24206), .Z(n24203) );
  AND U31465 ( .A(a[76]), .B(b[14]), .Z(n24202) );
  XOR U31466 ( .A(n24208), .B(n24209), .Z(n23673) );
  ANDN U31467 ( .B(n24210), .A(n24211), .Z(n24208) );
  AND U31468 ( .A(a[77]), .B(b[13]), .Z(n24207) );
  XOR U31469 ( .A(n24213), .B(n24214), .Z(n23678) );
  ANDN U31470 ( .B(n24215), .A(n24216), .Z(n24213) );
  AND U31471 ( .A(a[78]), .B(b[12]), .Z(n24212) );
  XOR U31472 ( .A(n24218), .B(n24219), .Z(n23683) );
  ANDN U31473 ( .B(n24220), .A(n24221), .Z(n24218) );
  AND U31474 ( .A(a[79]), .B(b[11]), .Z(n24217) );
  XOR U31475 ( .A(n24223), .B(n24224), .Z(n23688) );
  ANDN U31476 ( .B(n24225), .A(n24226), .Z(n24223) );
  AND U31477 ( .A(a[80]), .B(b[10]), .Z(n24222) );
  XOR U31478 ( .A(n24228), .B(n24229), .Z(n23693) );
  ANDN U31479 ( .B(n24230), .A(n24231), .Z(n24228) );
  AND U31480 ( .A(b[9]), .B(a[81]), .Z(n24227) );
  XOR U31481 ( .A(n24233), .B(n24234), .Z(n23698) );
  ANDN U31482 ( .B(n24235), .A(n24236), .Z(n24233) );
  AND U31483 ( .A(b[8]), .B(a[82]), .Z(n24232) );
  XOR U31484 ( .A(n24238), .B(n24239), .Z(n23703) );
  ANDN U31485 ( .B(n24240), .A(n24241), .Z(n24238) );
  AND U31486 ( .A(b[7]), .B(a[83]), .Z(n24237) );
  XOR U31487 ( .A(n24243), .B(n24244), .Z(n23708) );
  ANDN U31488 ( .B(n24245), .A(n24246), .Z(n24243) );
  AND U31489 ( .A(b[6]), .B(a[84]), .Z(n24242) );
  XOR U31490 ( .A(n24248), .B(n24249), .Z(n23713) );
  ANDN U31491 ( .B(n24250), .A(n24251), .Z(n24248) );
  AND U31492 ( .A(b[5]), .B(a[85]), .Z(n24247) );
  XOR U31493 ( .A(n24253), .B(n24254), .Z(n23718) );
  ANDN U31494 ( .B(n24255), .A(n24256), .Z(n24253) );
  AND U31495 ( .A(b[4]), .B(a[86]), .Z(n24252) );
  XOR U31496 ( .A(n24258), .B(n24259), .Z(n23723) );
  ANDN U31497 ( .B(n23735), .A(n23736), .Z(n24258) );
  AND U31498 ( .A(b[2]), .B(a[87]), .Z(n24260) );
  XNOR U31499 ( .A(n24255), .B(n24259), .Z(n24261) );
  XOR U31500 ( .A(n24262), .B(n24263), .Z(n24259) );
  OR U31501 ( .A(n23738), .B(n23739), .Z(n24263) );
  XNOR U31502 ( .A(n24265), .B(n24266), .Z(n24264) );
  XOR U31503 ( .A(n24265), .B(n24268), .Z(n23738) );
  NAND U31504 ( .A(b[1]), .B(a[87]), .Z(n24268) );
  IV U31505 ( .A(n24262), .Z(n24265) );
  NANDN U31506 ( .A(n29), .B(n30), .Z(n24262) );
  XOR U31507 ( .A(n24269), .B(n24270), .Z(n30) );
  NAND U31508 ( .A(a[87]), .B(b[0]), .Z(n29) );
  XNOR U31509 ( .A(n24250), .B(n24254), .Z(n24271) );
  XNOR U31510 ( .A(n24245), .B(n24249), .Z(n24272) );
  XNOR U31511 ( .A(n24240), .B(n24244), .Z(n24273) );
  XNOR U31512 ( .A(n24235), .B(n24239), .Z(n24274) );
  XNOR U31513 ( .A(n24230), .B(n24234), .Z(n24275) );
  XNOR U31514 ( .A(n24225), .B(n24229), .Z(n24276) );
  XNOR U31515 ( .A(n24220), .B(n24224), .Z(n24277) );
  XNOR U31516 ( .A(n24215), .B(n24219), .Z(n24278) );
  XNOR U31517 ( .A(n24210), .B(n24214), .Z(n24279) );
  XNOR U31518 ( .A(n24205), .B(n24209), .Z(n24280) );
  XNOR U31519 ( .A(n24200), .B(n24204), .Z(n24281) );
  XNOR U31520 ( .A(n24195), .B(n24199), .Z(n24282) );
  XNOR U31521 ( .A(n24190), .B(n24194), .Z(n24283) );
  XNOR U31522 ( .A(n24185), .B(n24189), .Z(n24284) );
  XNOR U31523 ( .A(n24180), .B(n24184), .Z(n24285) );
  XNOR U31524 ( .A(n24175), .B(n24179), .Z(n24286) );
  XNOR U31525 ( .A(n24170), .B(n24174), .Z(n24287) );
  XNOR U31526 ( .A(n24165), .B(n24169), .Z(n24288) );
  XNOR U31527 ( .A(n24160), .B(n24164), .Z(n24289) );
  XNOR U31528 ( .A(n24155), .B(n24159), .Z(n24290) );
  XNOR U31529 ( .A(n24150), .B(n24154), .Z(n24291) );
  XNOR U31530 ( .A(n24145), .B(n24149), .Z(n24292) );
  XNOR U31531 ( .A(n24140), .B(n24144), .Z(n24293) );
  XNOR U31532 ( .A(n24135), .B(n24139), .Z(n24294) );
  XNOR U31533 ( .A(n24130), .B(n24134), .Z(n24295) );
  XNOR U31534 ( .A(n24125), .B(n24129), .Z(n24296) );
  XNOR U31535 ( .A(n24120), .B(n24124), .Z(n24297) );
  XNOR U31536 ( .A(n24115), .B(n24119), .Z(n24298) );
  XNOR U31537 ( .A(n24110), .B(n24114), .Z(n24299) );
  XNOR U31538 ( .A(n24105), .B(n24109), .Z(n24300) );
  XNOR U31539 ( .A(n24100), .B(n24104), .Z(n24301) );
  XNOR U31540 ( .A(n24095), .B(n24099), .Z(n24302) );
  XNOR U31541 ( .A(n24090), .B(n24094), .Z(n24303) );
  XNOR U31542 ( .A(n24085), .B(n24089), .Z(n24304) );
  XNOR U31543 ( .A(n24080), .B(n24084), .Z(n24305) );
  XNOR U31544 ( .A(n24075), .B(n24079), .Z(n24306) );
  XNOR U31545 ( .A(n24070), .B(n24074), .Z(n24307) );
  XNOR U31546 ( .A(n24065), .B(n24069), .Z(n24308) );
  XNOR U31547 ( .A(n24060), .B(n24064), .Z(n24309) );
  XNOR U31548 ( .A(n24055), .B(n24059), .Z(n24310) );
  XNOR U31549 ( .A(n24050), .B(n24054), .Z(n24311) );
  XNOR U31550 ( .A(n24045), .B(n24049), .Z(n24312) );
  XNOR U31551 ( .A(n24040), .B(n24044), .Z(n24313) );
  XNOR U31552 ( .A(n24035), .B(n24039), .Z(n24314) );
  XNOR U31553 ( .A(n24030), .B(n24034), .Z(n24315) );
  XNOR U31554 ( .A(n24025), .B(n24029), .Z(n24316) );
  XNOR U31555 ( .A(n24020), .B(n24024), .Z(n24317) );
  XNOR U31556 ( .A(n24015), .B(n24019), .Z(n24318) );
  XNOR U31557 ( .A(n24010), .B(n24014), .Z(n24319) );
  XNOR U31558 ( .A(n24005), .B(n24009), .Z(n24320) );
  XNOR U31559 ( .A(n24000), .B(n24004), .Z(n24321) );
  XNOR U31560 ( .A(n23995), .B(n23999), .Z(n24322) );
  XNOR U31561 ( .A(n23990), .B(n23994), .Z(n24323) );
  XNOR U31562 ( .A(n23985), .B(n23989), .Z(n24324) );
  XNOR U31563 ( .A(n23980), .B(n23984), .Z(n24325) );
  XNOR U31564 ( .A(n23975), .B(n23979), .Z(n24326) );
  XNOR U31565 ( .A(n23970), .B(n23974), .Z(n24327) );
  XNOR U31566 ( .A(n23965), .B(n23969), .Z(n24328) );
  XNOR U31567 ( .A(n23960), .B(n23964), .Z(n24329) );
  XNOR U31568 ( .A(n23955), .B(n23959), .Z(n24330) );
  XNOR U31569 ( .A(n23950), .B(n23954), .Z(n24331) );
  XNOR U31570 ( .A(n23945), .B(n23949), .Z(n24332) );
  XNOR U31571 ( .A(n23940), .B(n23944), .Z(n24333) );
  XNOR U31572 ( .A(n23935), .B(n23939), .Z(n24334) );
  XNOR U31573 ( .A(n23930), .B(n23934), .Z(n24335) );
  XNOR U31574 ( .A(n23925), .B(n23929), .Z(n24336) );
  XNOR U31575 ( .A(n23920), .B(n23924), .Z(n24337) );
  XNOR U31576 ( .A(n23915), .B(n23919), .Z(n24338) );
  XNOR U31577 ( .A(n23910), .B(n23914), .Z(n24339) );
  XNOR U31578 ( .A(n23905), .B(n23909), .Z(n24340) );
  XNOR U31579 ( .A(n23900), .B(n23904), .Z(n24341) );
  XNOR U31580 ( .A(n23895), .B(n23899), .Z(n24342) );
  XNOR U31581 ( .A(n23890), .B(n23894), .Z(n24343) );
  XNOR U31582 ( .A(n23885), .B(n23889), .Z(n24344) );
  XNOR U31583 ( .A(n23880), .B(n23884), .Z(n24345) );
  XNOR U31584 ( .A(n23875), .B(n23879), .Z(n24346) );
  XNOR U31585 ( .A(n23870), .B(n23874), .Z(n24347) );
  XNOR U31586 ( .A(n23865), .B(n23869), .Z(n24348) );
  XNOR U31587 ( .A(n23860), .B(n23864), .Z(n24349) );
  XNOR U31588 ( .A(n23855), .B(n23859), .Z(n24350) );
  XNOR U31589 ( .A(n23850), .B(n23854), .Z(n24351) );
  XNOR U31590 ( .A(n23845), .B(n23849), .Z(n24352) );
  XNOR U31591 ( .A(n23840), .B(n23844), .Z(n24353) );
  XNOR U31592 ( .A(n23835), .B(n23839), .Z(n24354) );
  XNOR U31593 ( .A(n23830), .B(n23834), .Z(n24355) );
  XNOR U31594 ( .A(n24356), .B(n23829), .Z(n23830) );
  AND U31595 ( .A(a[0]), .B(b[89]), .Z(n24356) );
  XOR U31596 ( .A(n24357), .B(n23829), .Z(n23831) );
  XNOR U31597 ( .A(n24358), .B(n24359), .Z(n23829) );
  ANDN U31598 ( .B(n24360), .A(n24361), .Z(n24358) );
  AND U31599 ( .A(a[1]), .B(b[88]), .Z(n24357) );
  XOR U31600 ( .A(n24363), .B(n24364), .Z(n23834) );
  ANDN U31601 ( .B(n24365), .A(n24366), .Z(n24363) );
  AND U31602 ( .A(a[2]), .B(b[87]), .Z(n24362) );
  XOR U31603 ( .A(n24368), .B(n24369), .Z(n23839) );
  ANDN U31604 ( .B(n24370), .A(n24371), .Z(n24368) );
  AND U31605 ( .A(a[3]), .B(b[86]), .Z(n24367) );
  XOR U31606 ( .A(n24373), .B(n24374), .Z(n23844) );
  ANDN U31607 ( .B(n24375), .A(n24376), .Z(n24373) );
  AND U31608 ( .A(a[4]), .B(b[85]), .Z(n24372) );
  XOR U31609 ( .A(n24378), .B(n24379), .Z(n23849) );
  ANDN U31610 ( .B(n24380), .A(n24381), .Z(n24378) );
  AND U31611 ( .A(a[5]), .B(b[84]), .Z(n24377) );
  XOR U31612 ( .A(n24383), .B(n24384), .Z(n23854) );
  ANDN U31613 ( .B(n24385), .A(n24386), .Z(n24383) );
  AND U31614 ( .A(a[6]), .B(b[83]), .Z(n24382) );
  XOR U31615 ( .A(n24388), .B(n24389), .Z(n23859) );
  ANDN U31616 ( .B(n24390), .A(n24391), .Z(n24388) );
  AND U31617 ( .A(a[7]), .B(b[82]), .Z(n24387) );
  XOR U31618 ( .A(n24393), .B(n24394), .Z(n23864) );
  ANDN U31619 ( .B(n24395), .A(n24396), .Z(n24393) );
  AND U31620 ( .A(a[8]), .B(b[81]), .Z(n24392) );
  XOR U31621 ( .A(n24398), .B(n24399), .Z(n23869) );
  ANDN U31622 ( .B(n24400), .A(n24401), .Z(n24398) );
  AND U31623 ( .A(a[9]), .B(b[80]), .Z(n24397) );
  XOR U31624 ( .A(n24403), .B(n24404), .Z(n23874) );
  ANDN U31625 ( .B(n24405), .A(n24406), .Z(n24403) );
  AND U31626 ( .A(a[10]), .B(b[79]), .Z(n24402) );
  XOR U31627 ( .A(n24408), .B(n24409), .Z(n23879) );
  ANDN U31628 ( .B(n24410), .A(n24411), .Z(n24408) );
  AND U31629 ( .A(a[11]), .B(b[78]), .Z(n24407) );
  XOR U31630 ( .A(n24413), .B(n24414), .Z(n23884) );
  ANDN U31631 ( .B(n24415), .A(n24416), .Z(n24413) );
  AND U31632 ( .A(a[12]), .B(b[77]), .Z(n24412) );
  XOR U31633 ( .A(n24418), .B(n24419), .Z(n23889) );
  ANDN U31634 ( .B(n24420), .A(n24421), .Z(n24418) );
  AND U31635 ( .A(a[13]), .B(b[76]), .Z(n24417) );
  XOR U31636 ( .A(n24423), .B(n24424), .Z(n23894) );
  ANDN U31637 ( .B(n24425), .A(n24426), .Z(n24423) );
  AND U31638 ( .A(a[14]), .B(b[75]), .Z(n24422) );
  XOR U31639 ( .A(n24428), .B(n24429), .Z(n23899) );
  ANDN U31640 ( .B(n24430), .A(n24431), .Z(n24428) );
  AND U31641 ( .A(a[15]), .B(b[74]), .Z(n24427) );
  XOR U31642 ( .A(n24433), .B(n24434), .Z(n23904) );
  ANDN U31643 ( .B(n24435), .A(n24436), .Z(n24433) );
  AND U31644 ( .A(a[16]), .B(b[73]), .Z(n24432) );
  XOR U31645 ( .A(n24438), .B(n24439), .Z(n23909) );
  ANDN U31646 ( .B(n24440), .A(n24441), .Z(n24438) );
  AND U31647 ( .A(a[17]), .B(b[72]), .Z(n24437) );
  XOR U31648 ( .A(n24443), .B(n24444), .Z(n23914) );
  ANDN U31649 ( .B(n24445), .A(n24446), .Z(n24443) );
  AND U31650 ( .A(a[18]), .B(b[71]), .Z(n24442) );
  XOR U31651 ( .A(n24448), .B(n24449), .Z(n23919) );
  ANDN U31652 ( .B(n24450), .A(n24451), .Z(n24448) );
  AND U31653 ( .A(a[19]), .B(b[70]), .Z(n24447) );
  XOR U31654 ( .A(n24453), .B(n24454), .Z(n23924) );
  ANDN U31655 ( .B(n24455), .A(n24456), .Z(n24453) );
  AND U31656 ( .A(a[20]), .B(b[69]), .Z(n24452) );
  XOR U31657 ( .A(n24458), .B(n24459), .Z(n23929) );
  ANDN U31658 ( .B(n24460), .A(n24461), .Z(n24458) );
  AND U31659 ( .A(a[21]), .B(b[68]), .Z(n24457) );
  XOR U31660 ( .A(n24463), .B(n24464), .Z(n23934) );
  ANDN U31661 ( .B(n24465), .A(n24466), .Z(n24463) );
  AND U31662 ( .A(a[22]), .B(b[67]), .Z(n24462) );
  XOR U31663 ( .A(n24468), .B(n24469), .Z(n23939) );
  ANDN U31664 ( .B(n24470), .A(n24471), .Z(n24468) );
  AND U31665 ( .A(a[23]), .B(b[66]), .Z(n24467) );
  XOR U31666 ( .A(n24473), .B(n24474), .Z(n23944) );
  ANDN U31667 ( .B(n24475), .A(n24476), .Z(n24473) );
  AND U31668 ( .A(a[24]), .B(b[65]), .Z(n24472) );
  XOR U31669 ( .A(n24478), .B(n24479), .Z(n23949) );
  ANDN U31670 ( .B(n24480), .A(n24481), .Z(n24478) );
  AND U31671 ( .A(a[25]), .B(b[64]), .Z(n24477) );
  XOR U31672 ( .A(n24483), .B(n24484), .Z(n23954) );
  ANDN U31673 ( .B(n24485), .A(n24486), .Z(n24483) );
  AND U31674 ( .A(a[26]), .B(b[63]), .Z(n24482) );
  XOR U31675 ( .A(n24488), .B(n24489), .Z(n23959) );
  ANDN U31676 ( .B(n24490), .A(n24491), .Z(n24488) );
  AND U31677 ( .A(a[27]), .B(b[62]), .Z(n24487) );
  XOR U31678 ( .A(n24493), .B(n24494), .Z(n23964) );
  ANDN U31679 ( .B(n24495), .A(n24496), .Z(n24493) );
  AND U31680 ( .A(a[28]), .B(b[61]), .Z(n24492) );
  XOR U31681 ( .A(n24498), .B(n24499), .Z(n23969) );
  ANDN U31682 ( .B(n24500), .A(n24501), .Z(n24498) );
  AND U31683 ( .A(a[29]), .B(b[60]), .Z(n24497) );
  XOR U31684 ( .A(n24503), .B(n24504), .Z(n23974) );
  ANDN U31685 ( .B(n24505), .A(n24506), .Z(n24503) );
  AND U31686 ( .A(a[30]), .B(b[59]), .Z(n24502) );
  XOR U31687 ( .A(n24508), .B(n24509), .Z(n23979) );
  ANDN U31688 ( .B(n24510), .A(n24511), .Z(n24508) );
  AND U31689 ( .A(a[31]), .B(b[58]), .Z(n24507) );
  XOR U31690 ( .A(n24513), .B(n24514), .Z(n23984) );
  ANDN U31691 ( .B(n24515), .A(n24516), .Z(n24513) );
  AND U31692 ( .A(a[32]), .B(b[57]), .Z(n24512) );
  XOR U31693 ( .A(n24518), .B(n24519), .Z(n23989) );
  ANDN U31694 ( .B(n24520), .A(n24521), .Z(n24518) );
  AND U31695 ( .A(a[33]), .B(b[56]), .Z(n24517) );
  XOR U31696 ( .A(n24523), .B(n24524), .Z(n23994) );
  ANDN U31697 ( .B(n24525), .A(n24526), .Z(n24523) );
  AND U31698 ( .A(a[34]), .B(b[55]), .Z(n24522) );
  XOR U31699 ( .A(n24528), .B(n24529), .Z(n23999) );
  ANDN U31700 ( .B(n24530), .A(n24531), .Z(n24528) );
  AND U31701 ( .A(a[35]), .B(b[54]), .Z(n24527) );
  XOR U31702 ( .A(n24533), .B(n24534), .Z(n24004) );
  ANDN U31703 ( .B(n24535), .A(n24536), .Z(n24533) );
  AND U31704 ( .A(a[36]), .B(b[53]), .Z(n24532) );
  XOR U31705 ( .A(n24538), .B(n24539), .Z(n24009) );
  ANDN U31706 ( .B(n24540), .A(n24541), .Z(n24538) );
  AND U31707 ( .A(a[37]), .B(b[52]), .Z(n24537) );
  XOR U31708 ( .A(n24543), .B(n24544), .Z(n24014) );
  ANDN U31709 ( .B(n24545), .A(n24546), .Z(n24543) );
  AND U31710 ( .A(a[38]), .B(b[51]), .Z(n24542) );
  XOR U31711 ( .A(n24548), .B(n24549), .Z(n24019) );
  ANDN U31712 ( .B(n24550), .A(n24551), .Z(n24548) );
  AND U31713 ( .A(a[39]), .B(b[50]), .Z(n24547) );
  XOR U31714 ( .A(n24553), .B(n24554), .Z(n24024) );
  ANDN U31715 ( .B(n24555), .A(n24556), .Z(n24553) );
  AND U31716 ( .A(a[40]), .B(b[49]), .Z(n24552) );
  XOR U31717 ( .A(n24558), .B(n24559), .Z(n24029) );
  ANDN U31718 ( .B(n24560), .A(n24561), .Z(n24558) );
  AND U31719 ( .A(a[41]), .B(b[48]), .Z(n24557) );
  XOR U31720 ( .A(n24563), .B(n24564), .Z(n24034) );
  ANDN U31721 ( .B(n24565), .A(n24566), .Z(n24563) );
  AND U31722 ( .A(a[42]), .B(b[47]), .Z(n24562) );
  XOR U31723 ( .A(n24568), .B(n24569), .Z(n24039) );
  ANDN U31724 ( .B(n24570), .A(n24571), .Z(n24568) );
  AND U31725 ( .A(a[43]), .B(b[46]), .Z(n24567) );
  XOR U31726 ( .A(n24573), .B(n24574), .Z(n24044) );
  ANDN U31727 ( .B(n24575), .A(n24576), .Z(n24573) );
  AND U31728 ( .A(a[44]), .B(b[45]), .Z(n24572) );
  XOR U31729 ( .A(n24578), .B(n24579), .Z(n24049) );
  ANDN U31730 ( .B(n24580), .A(n24581), .Z(n24578) );
  AND U31731 ( .A(a[45]), .B(b[44]), .Z(n24577) );
  XOR U31732 ( .A(n24583), .B(n24584), .Z(n24054) );
  ANDN U31733 ( .B(n24585), .A(n24586), .Z(n24583) );
  AND U31734 ( .A(a[46]), .B(b[43]), .Z(n24582) );
  XOR U31735 ( .A(n24588), .B(n24589), .Z(n24059) );
  ANDN U31736 ( .B(n24590), .A(n24591), .Z(n24588) );
  AND U31737 ( .A(a[47]), .B(b[42]), .Z(n24587) );
  XOR U31738 ( .A(n24593), .B(n24594), .Z(n24064) );
  ANDN U31739 ( .B(n24595), .A(n24596), .Z(n24593) );
  AND U31740 ( .A(a[48]), .B(b[41]), .Z(n24592) );
  XOR U31741 ( .A(n24598), .B(n24599), .Z(n24069) );
  ANDN U31742 ( .B(n24600), .A(n24601), .Z(n24598) );
  AND U31743 ( .A(a[49]), .B(b[40]), .Z(n24597) );
  XOR U31744 ( .A(n24603), .B(n24604), .Z(n24074) );
  ANDN U31745 ( .B(n24605), .A(n24606), .Z(n24603) );
  AND U31746 ( .A(a[50]), .B(b[39]), .Z(n24602) );
  XOR U31747 ( .A(n24608), .B(n24609), .Z(n24079) );
  ANDN U31748 ( .B(n24610), .A(n24611), .Z(n24608) );
  AND U31749 ( .A(a[51]), .B(b[38]), .Z(n24607) );
  XOR U31750 ( .A(n24613), .B(n24614), .Z(n24084) );
  ANDN U31751 ( .B(n24615), .A(n24616), .Z(n24613) );
  AND U31752 ( .A(a[52]), .B(b[37]), .Z(n24612) );
  XOR U31753 ( .A(n24618), .B(n24619), .Z(n24089) );
  ANDN U31754 ( .B(n24620), .A(n24621), .Z(n24618) );
  AND U31755 ( .A(a[53]), .B(b[36]), .Z(n24617) );
  XOR U31756 ( .A(n24623), .B(n24624), .Z(n24094) );
  ANDN U31757 ( .B(n24625), .A(n24626), .Z(n24623) );
  AND U31758 ( .A(a[54]), .B(b[35]), .Z(n24622) );
  XOR U31759 ( .A(n24628), .B(n24629), .Z(n24099) );
  ANDN U31760 ( .B(n24630), .A(n24631), .Z(n24628) );
  AND U31761 ( .A(a[55]), .B(b[34]), .Z(n24627) );
  XOR U31762 ( .A(n24633), .B(n24634), .Z(n24104) );
  ANDN U31763 ( .B(n24635), .A(n24636), .Z(n24633) );
  AND U31764 ( .A(a[56]), .B(b[33]), .Z(n24632) );
  XOR U31765 ( .A(n24638), .B(n24639), .Z(n24109) );
  ANDN U31766 ( .B(n24640), .A(n24641), .Z(n24638) );
  AND U31767 ( .A(a[57]), .B(b[32]), .Z(n24637) );
  XOR U31768 ( .A(n24643), .B(n24644), .Z(n24114) );
  ANDN U31769 ( .B(n24645), .A(n24646), .Z(n24643) );
  AND U31770 ( .A(a[58]), .B(b[31]), .Z(n24642) );
  XOR U31771 ( .A(n24648), .B(n24649), .Z(n24119) );
  ANDN U31772 ( .B(n24650), .A(n24651), .Z(n24648) );
  AND U31773 ( .A(a[59]), .B(b[30]), .Z(n24647) );
  XOR U31774 ( .A(n24653), .B(n24654), .Z(n24124) );
  ANDN U31775 ( .B(n24655), .A(n24656), .Z(n24653) );
  AND U31776 ( .A(a[60]), .B(b[29]), .Z(n24652) );
  XOR U31777 ( .A(n24658), .B(n24659), .Z(n24129) );
  ANDN U31778 ( .B(n24660), .A(n24661), .Z(n24658) );
  AND U31779 ( .A(a[61]), .B(b[28]), .Z(n24657) );
  XOR U31780 ( .A(n24663), .B(n24664), .Z(n24134) );
  ANDN U31781 ( .B(n24665), .A(n24666), .Z(n24663) );
  AND U31782 ( .A(a[62]), .B(b[27]), .Z(n24662) );
  XOR U31783 ( .A(n24668), .B(n24669), .Z(n24139) );
  ANDN U31784 ( .B(n24670), .A(n24671), .Z(n24668) );
  AND U31785 ( .A(a[63]), .B(b[26]), .Z(n24667) );
  XOR U31786 ( .A(n24673), .B(n24674), .Z(n24144) );
  ANDN U31787 ( .B(n24675), .A(n24676), .Z(n24673) );
  AND U31788 ( .A(a[64]), .B(b[25]), .Z(n24672) );
  XOR U31789 ( .A(n24678), .B(n24679), .Z(n24149) );
  ANDN U31790 ( .B(n24680), .A(n24681), .Z(n24678) );
  AND U31791 ( .A(a[65]), .B(b[24]), .Z(n24677) );
  XOR U31792 ( .A(n24683), .B(n24684), .Z(n24154) );
  ANDN U31793 ( .B(n24685), .A(n24686), .Z(n24683) );
  AND U31794 ( .A(a[66]), .B(b[23]), .Z(n24682) );
  XOR U31795 ( .A(n24688), .B(n24689), .Z(n24159) );
  ANDN U31796 ( .B(n24690), .A(n24691), .Z(n24688) );
  AND U31797 ( .A(a[67]), .B(b[22]), .Z(n24687) );
  XOR U31798 ( .A(n24693), .B(n24694), .Z(n24164) );
  ANDN U31799 ( .B(n24695), .A(n24696), .Z(n24693) );
  AND U31800 ( .A(a[68]), .B(b[21]), .Z(n24692) );
  XOR U31801 ( .A(n24698), .B(n24699), .Z(n24169) );
  ANDN U31802 ( .B(n24700), .A(n24701), .Z(n24698) );
  AND U31803 ( .A(a[69]), .B(b[20]), .Z(n24697) );
  XOR U31804 ( .A(n24703), .B(n24704), .Z(n24174) );
  ANDN U31805 ( .B(n24705), .A(n24706), .Z(n24703) );
  AND U31806 ( .A(a[70]), .B(b[19]), .Z(n24702) );
  XOR U31807 ( .A(n24708), .B(n24709), .Z(n24179) );
  ANDN U31808 ( .B(n24710), .A(n24711), .Z(n24708) );
  AND U31809 ( .A(a[71]), .B(b[18]), .Z(n24707) );
  XOR U31810 ( .A(n24713), .B(n24714), .Z(n24184) );
  ANDN U31811 ( .B(n24715), .A(n24716), .Z(n24713) );
  AND U31812 ( .A(a[72]), .B(b[17]), .Z(n24712) );
  XOR U31813 ( .A(n24718), .B(n24719), .Z(n24189) );
  ANDN U31814 ( .B(n24720), .A(n24721), .Z(n24718) );
  AND U31815 ( .A(a[73]), .B(b[16]), .Z(n24717) );
  XOR U31816 ( .A(n24723), .B(n24724), .Z(n24194) );
  ANDN U31817 ( .B(n24725), .A(n24726), .Z(n24723) );
  AND U31818 ( .A(a[74]), .B(b[15]), .Z(n24722) );
  XOR U31819 ( .A(n24728), .B(n24729), .Z(n24199) );
  ANDN U31820 ( .B(n24730), .A(n24731), .Z(n24728) );
  AND U31821 ( .A(a[75]), .B(b[14]), .Z(n24727) );
  XOR U31822 ( .A(n24733), .B(n24734), .Z(n24204) );
  ANDN U31823 ( .B(n24735), .A(n24736), .Z(n24733) );
  AND U31824 ( .A(a[76]), .B(b[13]), .Z(n24732) );
  XOR U31825 ( .A(n24738), .B(n24739), .Z(n24209) );
  ANDN U31826 ( .B(n24740), .A(n24741), .Z(n24738) );
  AND U31827 ( .A(a[77]), .B(b[12]), .Z(n24737) );
  XOR U31828 ( .A(n24743), .B(n24744), .Z(n24214) );
  ANDN U31829 ( .B(n24745), .A(n24746), .Z(n24743) );
  AND U31830 ( .A(a[78]), .B(b[11]), .Z(n24742) );
  XOR U31831 ( .A(n24748), .B(n24749), .Z(n24219) );
  ANDN U31832 ( .B(n24750), .A(n24751), .Z(n24748) );
  AND U31833 ( .A(a[79]), .B(b[10]), .Z(n24747) );
  XOR U31834 ( .A(n24753), .B(n24754), .Z(n24224) );
  ANDN U31835 ( .B(n24755), .A(n24756), .Z(n24753) );
  AND U31836 ( .A(b[9]), .B(a[80]), .Z(n24752) );
  XOR U31837 ( .A(n24758), .B(n24759), .Z(n24229) );
  ANDN U31838 ( .B(n24760), .A(n24761), .Z(n24758) );
  AND U31839 ( .A(b[8]), .B(a[81]), .Z(n24757) );
  XOR U31840 ( .A(n24763), .B(n24764), .Z(n24234) );
  ANDN U31841 ( .B(n24765), .A(n24766), .Z(n24763) );
  AND U31842 ( .A(b[7]), .B(a[82]), .Z(n24762) );
  XOR U31843 ( .A(n24768), .B(n24769), .Z(n24239) );
  ANDN U31844 ( .B(n24770), .A(n24771), .Z(n24768) );
  AND U31845 ( .A(b[6]), .B(a[83]), .Z(n24767) );
  XOR U31846 ( .A(n24773), .B(n24774), .Z(n24244) );
  ANDN U31847 ( .B(n24775), .A(n24776), .Z(n24773) );
  AND U31848 ( .A(b[5]), .B(a[84]), .Z(n24772) );
  XOR U31849 ( .A(n24778), .B(n24779), .Z(n24249) );
  ANDN U31850 ( .B(n24780), .A(n24781), .Z(n24778) );
  AND U31851 ( .A(b[4]), .B(a[85]), .Z(n24777) );
  XOR U31852 ( .A(n24783), .B(n24784), .Z(n24254) );
  ANDN U31853 ( .B(n24266), .A(n24267), .Z(n24783) );
  AND U31854 ( .A(b[2]), .B(a[86]), .Z(n24785) );
  XNOR U31855 ( .A(n24780), .B(n24784), .Z(n24786) );
  XOR U31856 ( .A(n24787), .B(n24788), .Z(n24784) );
  OR U31857 ( .A(n24269), .B(n24270), .Z(n24788) );
  XNOR U31858 ( .A(n24790), .B(n24791), .Z(n24789) );
  XOR U31859 ( .A(n24790), .B(n24793), .Z(n24269) );
  NAND U31860 ( .A(b[1]), .B(a[86]), .Z(n24793) );
  IV U31861 ( .A(n24787), .Z(n24790) );
  NANDN U31862 ( .A(n31), .B(n32), .Z(n24787) );
  XOR U31863 ( .A(n24794), .B(n24795), .Z(n32) );
  NAND U31864 ( .A(a[86]), .B(b[0]), .Z(n31) );
  XNOR U31865 ( .A(n24775), .B(n24779), .Z(n24796) );
  XNOR U31866 ( .A(n24770), .B(n24774), .Z(n24797) );
  XNOR U31867 ( .A(n24765), .B(n24769), .Z(n24798) );
  XNOR U31868 ( .A(n24760), .B(n24764), .Z(n24799) );
  XNOR U31869 ( .A(n24755), .B(n24759), .Z(n24800) );
  XNOR U31870 ( .A(n24750), .B(n24754), .Z(n24801) );
  XNOR U31871 ( .A(n24745), .B(n24749), .Z(n24802) );
  XNOR U31872 ( .A(n24740), .B(n24744), .Z(n24803) );
  XNOR U31873 ( .A(n24735), .B(n24739), .Z(n24804) );
  XNOR U31874 ( .A(n24730), .B(n24734), .Z(n24805) );
  XNOR U31875 ( .A(n24725), .B(n24729), .Z(n24806) );
  XNOR U31876 ( .A(n24720), .B(n24724), .Z(n24807) );
  XNOR U31877 ( .A(n24715), .B(n24719), .Z(n24808) );
  XNOR U31878 ( .A(n24710), .B(n24714), .Z(n24809) );
  XNOR U31879 ( .A(n24705), .B(n24709), .Z(n24810) );
  XNOR U31880 ( .A(n24700), .B(n24704), .Z(n24811) );
  XNOR U31881 ( .A(n24695), .B(n24699), .Z(n24812) );
  XNOR U31882 ( .A(n24690), .B(n24694), .Z(n24813) );
  XNOR U31883 ( .A(n24685), .B(n24689), .Z(n24814) );
  XNOR U31884 ( .A(n24680), .B(n24684), .Z(n24815) );
  XNOR U31885 ( .A(n24675), .B(n24679), .Z(n24816) );
  XNOR U31886 ( .A(n24670), .B(n24674), .Z(n24817) );
  XNOR U31887 ( .A(n24665), .B(n24669), .Z(n24818) );
  XNOR U31888 ( .A(n24660), .B(n24664), .Z(n24819) );
  XNOR U31889 ( .A(n24655), .B(n24659), .Z(n24820) );
  XNOR U31890 ( .A(n24650), .B(n24654), .Z(n24821) );
  XNOR U31891 ( .A(n24645), .B(n24649), .Z(n24822) );
  XNOR U31892 ( .A(n24640), .B(n24644), .Z(n24823) );
  XNOR U31893 ( .A(n24635), .B(n24639), .Z(n24824) );
  XNOR U31894 ( .A(n24630), .B(n24634), .Z(n24825) );
  XNOR U31895 ( .A(n24625), .B(n24629), .Z(n24826) );
  XNOR U31896 ( .A(n24620), .B(n24624), .Z(n24827) );
  XNOR U31897 ( .A(n24615), .B(n24619), .Z(n24828) );
  XNOR U31898 ( .A(n24610), .B(n24614), .Z(n24829) );
  XNOR U31899 ( .A(n24605), .B(n24609), .Z(n24830) );
  XNOR U31900 ( .A(n24600), .B(n24604), .Z(n24831) );
  XNOR U31901 ( .A(n24595), .B(n24599), .Z(n24832) );
  XNOR U31902 ( .A(n24590), .B(n24594), .Z(n24833) );
  XNOR U31903 ( .A(n24585), .B(n24589), .Z(n24834) );
  XNOR U31904 ( .A(n24580), .B(n24584), .Z(n24835) );
  XNOR U31905 ( .A(n24575), .B(n24579), .Z(n24836) );
  XNOR U31906 ( .A(n24570), .B(n24574), .Z(n24837) );
  XNOR U31907 ( .A(n24565), .B(n24569), .Z(n24838) );
  XNOR U31908 ( .A(n24560), .B(n24564), .Z(n24839) );
  XNOR U31909 ( .A(n24555), .B(n24559), .Z(n24840) );
  XNOR U31910 ( .A(n24550), .B(n24554), .Z(n24841) );
  XNOR U31911 ( .A(n24545), .B(n24549), .Z(n24842) );
  XNOR U31912 ( .A(n24540), .B(n24544), .Z(n24843) );
  XNOR U31913 ( .A(n24535), .B(n24539), .Z(n24844) );
  XNOR U31914 ( .A(n24530), .B(n24534), .Z(n24845) );
  XNOR U31915 ( .A(n24525), .B(n24529), .Z(n24846) );
  XNOR U31916 ( .A(n24520), .B(n24524), .Z(n24847) );
  XNOR U31917 ( .A(n24515), .B(n24519), .Z(n24848) );
  XNOR U31918 ( .A(n24510), .B(n24514), .Z(n24849) );
  XNOR U31919 ( .A(n24505), .B(n24509), .Z(n24850) );
  XNOR U31920 ( .A(n24500), .B(n24504), .Z(n24851) );
  XNOR U31921 ( .A(n24495), .B(n24499), .Z(n24852) );
  XNOR U31922 ( .A(n24490), .B(n24494), .Z(n24853) );
  XNOR U31923 ( .A(n24485), .B(n24489), .Z(n24854) );
  XNOR U31924 ( .A(n24480), .B(n24484), .Z(n24855) );
  XNOR U31925 ( .A(n24475), .B(n24479), .Z(n24856) );
  XNOR U31926 ( .A(n24470), .B(n24474), .Z(n24857) );
  XNOR U31927 ( .A(n24465), .B(n24469), .Z(n24858) );
  XNOR U31928 ( .A(n24859), .B(n24860), .Z(n24465) );
  XNOR U31929 ( .A(n24460), .B(n24464), .Z(n24860) );
  XNOR U31930 ( .A(n24455), .B(n24459), .Z(n24861) );
  XNOR U31931 ( .A(n24862), .B(n24863), .Z(n24455) );
  XNOR U31932 ( .A(n24450), .B(n24454), .Z(n24863) );
  XNOR U31933 ( .A(n24864), .B(n24865), .Z(n24450) );
  XNOR U31934 ( .A(n24445), .B(n24449), .Z(n24865) );
  XNOR U31935 ( .A(n24440), .B(n24444), .Z(n24866) );
  XNOR U31936 ( .A(n24435), .B(n24439), .Z(n24867) );
  XNOR U31937 ( .A(n24430), .B(n24434), .Z(n24868) );
  XNOR U31938 ( .A(n24425), .B(n24429), .Z(n24869) );
  XNOR U31939 ( .A(n24420), .B(n24424), .Z(n24870) );
  XNOR U31940 ( .A(n24415), .B(n24419), .Z(n24871) );
  XNOR U31941 ( .A(n24410), .B(n24414), .Z(n24872) );
  XNOR U31942 ( .A(n24405), .B(n24409), .Z(n24873) );
  XNOR U31943 ( .A(n24400), .B(n24404), .Z(n24874) );
  XNOR U31944 ( .A(n24395), .B(n24399), .Z(n24875) );
  XNOR U31945 ( .A(n24390), .B(n24394), .Z(n24876) );
  XNOR U31946 ( .A(n24385), .B(n24389), .Z(n24877) );
  XNOR U31947 ( .A(n24380), .B(n24384), .Z(n24878) );
  XNOR U31948 ( .A(n24375), .B(n24379), .Z(n24879) );
  XNOR U31949 ( .A(n24370), .B(n24374), .Z(n24880) );
  XNOR U31950 ( .A(n24365), .B(n24369), .Z(n24881) );
  XNOR U31951 ( .A(n24360), .B(n24364), .Z(n24882) );
  XOR U31952 ( .A(n24883), .B(n24359), .Z(n24360) );
  AND U31953 ( .A(a[0]), .B(b[88]), .Z(n24883) );
  XNOR U31954 ( .A(n24884), .B(n24359), .Z(n24361) );
  XNOR U31955 ( .A(n24885), .B(n24886), .Z(n24359) );
  ANDN U31956 ( .B(n24887), .A(n24888), .Z(n24885) );
  AND U31957 ( .A(a[1]), .B(b[87]), .Z(n24884) );
  XOR U31958 ( .A(n24890), .B(n24891), .Z(n24364) );
  ANDN U31959 ( .B(n24892), .A(n24893), .Z(n24890) );
  AND U31960 ( .A(a[2]), .B(b[86]), .Z(n24889) );
  XOR U31961 ( .A(n24895), .B(n24896), .Z(n24369) );
  ANDN U31962 ( .B(n24897), .A(n24898), .Z(n24895) );
  AND U31963 ( .A(a[3]), .B(b[85]), .Z(n24894) );
  XOR U31964 ( .A(n24900), .B(n24901), .Z(n24374) );
  ANDN U31965 ( .B(n24902), .A(n24903), .Z(n24900) );
  AND U31966 ( .A(a[4]), .B(b[84]), .Z(n24899) );
  XOR U31967 ( .A(n24905), .B(n24906), .Z(n24379) );
  ANDN U31968 ( .B(n24907), .A(n24908), .Z(n24905) );
  AND U31969 ( .A(a[5]), .B(b[83]), .Z(n24904) );
  XOR U31970 ( .A(n24910), .B(n24911), .Z(n24384) );
  ANDN U31971 ( .B(n24912), .A(n24913), .Z(n24910) );
  AND U31972 ( .A(a[6]), .B(b[82]), .Z(n24909) );
  XOR U31973 ( .A(n24915), .B(n24916), .Z(n24389) );
  ANDN U31974 ( .B(n24917), .A(n24918), .Z(n24915) );
  AND U31975 ( .A(a[7]), .B(b[81]), .Z(n24914) );
  XOR U31976 ( .A(n24920), .B(n24921), .Z(n24394) );
  ANDN U31977 ( .B(n24922), .A(n24923), .Z(n24920) );
  AND U31978 ( .A(a[8]), .B(b[80]), .Z(n24919) );
  XOR U31979 ( .A(n24925), .B(n24926), .Z(n24399) );
  ANDN U31980 ( .B(n24927), .A(n24928), .Z(n24925) );
  AND U31981 ( .A(a[9]), .B(b[79]), .Z(n24924) );
  XOR U31982 ( .A(n24930), .B(n24931), .Z(n24404) );
  ANDN U31983 ( .B(n24932), .A(n24933), .Z(n24930) );
  AND U31984 ( .A(a[10]), .B(b[78]), .Z(n24929) );
  XOR U31985 ( .A(n24935), .B(n24936), .Z(n24409) );
  ANDN U31986 ( .B(n24937), .A(n24938), .Z(n24935) );
  AND U31987 ( .A(a[11]), .B(b[77]), .Z(n24934) );
  XOR U31988 ( .A(n24940), .B(n24941), .Z(n24414) );
  ANDN U31989 ( .B(n24942), .A(n24943), .Z(n24940) );
  AND U31990 ( .A(a[12]), .B(b[76]), .Z(n24939) );
  XOR U31991 ( .A(n24945), .B(n24946), .Z(n24419) );
  ANDN U31992 ( .B(n24947), .A(n24948), .Z(n24945) );
  AND U31993 ( .A(a[13]), .B(b[75]), .Z(n24944) );
  XOR U31994 ( .A(n24950), .B(n24951), .Z(n24424) );
  ANDN U31995 ( .B(n24952), .A(n24953), .Z(n24950) );
  AND U31996 ( .A(a[14]), .B(b[74]), .Z(n24949) );
  XOR U31997 ( .A(n24955), .B(n24956), .Z(n24429) );
  ANDN U31998 ( .B(n24957), .A(n24958), .Z(n24955) );
  AND U31999 ( .A(a[15]), .B(b[73]), .Z(n24954) );
  XOR U32000 ( .A(n24960), .B(n24961), .Z(n24434) );
  ANDN U32001 ( .B(n24962), .A(n24963), .Z(n24960) );
  AND U32002 ( .A(a[16]), .B(b[72]), .Z(n24959) );
  XOR U32003 ( .A(n24965), .B(n24966), .Z(n24439) );
  ANDN U32004 ( .B(n24967), .A(n24968), .Z(n24965) );
  AND U32005 ( .A(a[17]), .B(b[71]), .Z(n24964) );
  IV U32006 ( .A(n24446), .Z(n24864) );
  XOR U32007 ( .A(n24970), .B(n24971), .Z(n24444) );
  ANDN U32008 ( .B(n24972), .A(n24973), .Z(n24970) );
  AND U32009 ( .A(a[18]), .B(b[70]), .Z(n24969) );
  IV U32010 ( .A(n24451), .Z(n24862) );
  XOR U32011 ( .A(n24975), .B(n24976), .Z(n24449) );
  ANDN U32012 ( .B(n24977), .A(n24978), .Z(n24975) );
  AND U32013 ( .A(a[19]), .B(b[69]), .Z(n24974) );
  XOR U32014 ( .A(n24980), .B(n24981), .Z(n24454) );
  ANDN U32015 ( .B(n24982), .A(n24983), .Z(n24980) );
  AND U32016 ( .A(a[20]), .B(b[68]), .Z(n24979) );
  IV U32017 ( .A(n24461), .Z(n24859) );
  XOR U32018 ( .A(n24985), .B(n24986), .Z(n24459) );
  ANDN U32019 ( .B(n24987), .A(n24988), .Z(n24985) );
  AND U32020 ( .A(a[21]), .B(b[67]), .Z(n24984) );
  XOR U32021 ( .A(n24989), .B(n24990), .Z(n24466) );
  IV U32022 ( .A(n24464), .Z(n24990) );
  XOR U32023 ( .A(n24991), .B(n24992), .Z(n24464) );
  ANDN U32024 ( .B(n24993), .A(n24994), .Z(n24991) );
  AND U32025 ( .A(a[22]), .B(b[66]), .Z(n24989) );
  XOR U32026 ( .A(n24996), .B(n24997), .Z(n24469) );
  ANDN U32027 ( .B(n24998), .A(n24999), .Z(n24996) );
  AND U32028 ( .A(a[23]), .B(b[65]), .Z(n24995) );
  XOR U32029 ( .A(n25001), .B(n25002), .Z(n24474) );
  ANDN U32030 ( .B(n25003), .A(n25004), .Z(n25001) );
  AND U32031 ( .A(a[24]), .B(b[64]), .Z(n25000) );
  XOR U32032 ( .A(n25006), .B(n25007), .Z(n24479) );
  ANDN U32033 ( .B(n25008), .A(n25009), .Z(n25006) );
  AND U32034 ( .A(a[25]), .B(b[63]), .Z(n25005) );
  XOR U32035 ( .A(n25011), .B(n25012), .Z(n24484) );
  ANDN U32036 ( .B(n25013), .A(n25014), .Z(n25011) );
  AND U32037 ( .A(a[26]), .B(b[62]), .Z(n25010) );
  XOR U32038 ( .A(n25016), .B(n25017), .Z(n24489) );
  ANDN U32039 ( .B(n25018), .A(n25019), .Z(n25016) );
  AND U32040 ( .A(a[27]), .B(b[61]), .Z(n25015) );
  XOR U32041 ( .A(n25021), .B(n25022), .Z(n24494) );
  ANDN U32042 ( .B(n25023), .A(n25024), .Z(n25021) );
  AND U32043 ( .A(a[28]), .B(b[60]), .Z(n25020) );
  XOR U32044 ( .A(n25026), .B(n25027), .Z(n24499) );
  ANDN U32045 ( .B(n25028), .A(n25029), .Z(n25026) );
  AND U32046 ( .A(a[29]), .B(b[59]), .Z(n25025) );
  XOR U32047 ( .A(n25031), .B(n25032), .Z(n24504) );
  ANDN U32048 ( .B(n25033), .A(n25034), .Z(n25031) );
  AND U32049 ( .A(a[30]), .B(b[58]), .Z(n25030) );
  XOR U32050 ( .A(n25036), .B(n25037), .Z(n24509) );
  ANDN U32051 ( .B(n25038), .A(n25039), .Z(n25036) );
  AND U32052 ( .A(a[31]), .B(b[57]), .Z(n25035) );
  XOR U32053 ( .A(n25041), .B(n25042), .Z(n24514) );
  ANDN U32054 ( .B(n25043), .A(n25044), .Z(n25041) );
  AND U32055 ( .A(a[32]), .B(b[56]), .Z(n25040) );
  XOR U32056 ( .A(n25046), .B(n25047), .Z(n24519) );
  ANDN U32057 ( .B(n25048), .A(n25049), .Z(n25046) );
  AND U32058 ( .A(a[33]), .B(b[55]), .Z(n25045) );
  XOR U32059 ( .A(n25051), .B(n25052), .Z(n24524) );
  ANDN U32060 ( .B(n25053), .A(n25054), .Z(n25051) );
  AND U32061 ( .A(a[34]), .B(b[54]), .Z(n25050) );
  XOR U32062 ( .A(n25056), .B(n25057), .Z(n24529) );
  ANDN U32063 ( .B(n25058), .A(n25059), .Z(n25056) );
  AND U32064 ( .A(a[35]), .B(b[53]), .Z(n25055) );
  XOR U32065 ( .A(n25061), .B(n25062), .Z(n24534) );
  ANDN U32066 ( .B(n25063), .A(n25064), .Z(n25061) );
  AND U32067 ( .A(a[36]), .B(b[52]), .Z(n25060) );
  XOR U32068 ( .A(n25066), .B(n25067), .Z(n24539) );
  ANDN U32069 ( .B(n25068), .A(n25069), .Z(n25066) );
  AND U32070 ( .A(a[37]), .B(b[51]), .Z(n25065) );
  XOR U32071 ( .A(n25071), .B(n25072), .Z(n24544) );
  ANDN U32072 ( .B(n25073), .A(n25074), .Z(n25071) );
  AND U32073 ( .A(a[38]), .B(b[50]), .Z(n25070) );
  XOR U32074 ( .A(n25076), .B(n25077), .Z(n24549) );
  ANDN U32075 ( .B(n25078), .A(n25079), .Z(n25076) );
  AND U32076 ( .A(a[39]), .B(b[49]), .Z(n25075) );
  XOR U32077 ( .A(n25081), .B(n25082), .Z(n24554) );
  ANDN U32078 ( .B(n25083), .A(n25084), .Z(n25081) );
  AND U32079 ( .A(a[40]), .B(b[48]), .Z(n25080) );
  XOR U32080 ( .A(n25086), .B(n25087), .Z(n24559) );
  ANDN U32081 ( .B(n25088), .A(n25089), .Z(n25086) );
  AND U32082 ( .A(a[41]), .B(b[47]), .Z(n25085) );
  XOR U32083 ( .A(n25091), .B(n25092), .Z(n24564) );
  ANDN U32084 ( .B(n25093), .A(n25094), .Z(n25091) );
  AND U32085 ( .A(a[42]), .B(b[46]), .Z(n25090) );
  XOR U32086 ( .A(n25096), .B(n25097), .Z(n24569) );
  ANDN U32087 ( .B(n25098), .A(n25099), .Z(n25096) );
  AND U32088 ( .A(a[43]), .B(b[45]), .Z(n25095) );
  XOR U32089 ( .A(n25101), .B(n25102), .Z(n24574) );
  ANDN U32090 ( .B(n25103), .A(n25104), .Z(n25101) );
  AND U32091 ( .A(a[44]), .B(b[44]), .Z(n25100) );
  XOR U32092 ( .A(n25106), .B(n25107), .Z(n24579) );
  ANDN U32093 ( .B(n25108), .A(n25109), .Z(n25106) );
  AND U32094 ( .A(a[45]), .B(b[43]), .Z(n25105) );
  XOR U32095 ( .A(n25111), .B(n25112), .Z(n24584) );
  ANDN U32096 ( .B(n25113), .A(n25114), .Z(n25111) );
  AND U32097 ( .A(a[46]), .B(b[42]), .Z(n25110) );
  XOR U32098 ( .A(n25116), .B(n25117), .Z(n24589) );
  ANDN U32099 ( .B(n25118), .A(n25119), .Z(n25116) );
  AND U32100 ( .A(a[47]), .B(b[41]), .Z(n25115) );
  XOR U32101 ( .A(n25121), .B(n25122), .Z(n24594) );
  ANDN U32102 ( .B(n25123), .A(n25124), .Z(n25121) );
  AND U32103 ( .A(a[48]), .B(b[40]), .Z(n25120) );
  XOR U32104 ( .A(n25126), .B(n25127), .Z(n24599) );
  ANDN U32105 ( .B(n25128), .A(n25129), .Z(n25126) );
  AND U32106 ( .A(a[49]), .B(b[39]), .Z(n25125) );
  XOR U32107 ( .A(n25131), .B(n25132), .Z(n24604) );
  ANDN U32108 ( .B(n25133), .A(n25134), .Z(n25131) );
  AND U32109 ( .A(a[50]), .B(b[38]), .Z(n25130) );
  XOR U32110 ( .A(n25136), .B(n25137), .Z(n24609) );
  ANDN U32111 ( .B(n25138), .A(n25139), .Z(n25136) );
  AND U32112 ( .A(a[51]), .B(b[37]), .Z(n25135) );
  XOR U32113 ( .A(n25141), .B(n25142), .Z(n24614) );
  ANDN U32114 ( .B(n25143), .A(n25144), .Z(n25141) );
  AND U32115 ( .A(a[52]), .B(b[36]), .Z(n25140) );
  XOR U32116 ( .A(n25146), .B(n25147), .Z(n24619) );
  ANDN U32117 ( .B(n25148), .A(n25149), .Z(n25146) );
  AND U32118 ( .A(a[53]), .B(b[35]), .Z(n25145) );
  XOR U32119 ( .A(n25151), .B(n25152), .Z(n24624) );
  ANDN U32120 ( .B(n25153), .A(n25154), .Z(n25151) );
  AND U32121 ( .A(a[54]), .B(b[34]), .Z(n25150) );
  XOR U32122 ( .A(n25156), .B(n25157), .Z(n24629) );
  ANDN U32123 ( .B(n25158), .A(n25159), .Z(n25156) );
  AND U32124 ( .A(a[55]), .B(b[33]), .Z(n25155) );
  XOR U32125 ( .A(n25161), .B(n25162), .Z(n24634) );
  ANDN U32126 ( .B(n25163), .A(n25164), .Z(n25161) );
  AND U32127 ( .A(a[56]), .B(b[32]), .Z(n25160) );
  XOR U32128 ( .A(n25166), .B(n25167), .Z(n24639) );
  ANDN U32129 ( .B(n25168), .A(n25169), .Z(n25166) );
  AND U32130 ( .A(a[57]), .B(b[31]), .Z(n25165) );
  XOR U32131 ( .A(n25171), .B(n25172), .Z(n24644) );
  ANDN U32132 ( .B(n25173), .A(n25174), .Z(n25171) );
  AND U32133 ( .A(a[58]), .B(b[30]), .Z(n25170) );
  XOR U32134 ( .A(n25176), .B(n25177), .Z(n24649) );
  ANDN U32135 ( .B(n25178), .A(n25179), .Z(n25176) );
  AND U32136 ( .A(a[59]), .B(b[29]), .Z(n25175) );
  XOR U32137 ( .A(n25181), .B(n25182), .Z(n24654) );
  ANDN U32138 ( .B(n25183), .A(n25184), .Z(n25181) );
  AND U32139 ( .A(a[60]), .B(b[28]), .Z(n25180) );
  XOR U32140 ( .A(n25186), .B(n25187), .Z(n24659) );
  ANDN U32141 ( .B(n25188), .A(n25189), .Z(n25186) );
  AND U32142 ( .A(a[61]), .B(b[27]), .Z(n25185) );
  XOR U32143 ( .A(n25191), .B(n25192), .Z(n24664) );
  ANDN U32144 ( .B(n25193), .A(n25194), .Z(n25191) );
  AND U32145 ( .A(a[62]), .B(b[26]), .Z(n25190) );
  XOR U32146 ( .A(n25196), .B(n25197), .Z(n24669) );
  ANDN U32147 ( .B(n25198), .A(n25199), .Z(n25196) );
  AND U32148 ( .A(a[63]), .B(b[25]), .Z(n25195) );
  XOR U32149 ( .A(n25201), .B(n25202), .Z(n24674) );
  ANDN U32150 ( .B(n25203), .A(n25204), .Z(n25201) );
  AND U32151 ( .A(a[64]), .B(b[24]), .Z(n25200) );
  XOR U32152 ( .A(n25206), .B(n25207), .Z(n24679) );
  ANDN U32153 ( .B(n25208), .A(n25209), .Z(n25206) );
  AND U32154 ( .A(a[65]), .B(b[23]), .Z(n25205) );
  XOR U32155 ( .A(n25211), .B(n25212), .Z(n24684) );
  ANDN U32156 ( .B(n25213), .A(n25214), .Z(n25211) );
  AND U32157 ( .A(a[66]), .B(b[22]), .Z(n25210) );
  XOR U32158 ( .A(n25216), .B(n25217), .Z(n24689) );
  ANDN U32159 ( .B(n25218), .A(n25219), .Z(n25216) );
  AND U32160 ( .A(a[67]), .B(b[21]), .Z(n25215) );
  XOR U32161 ( .A(n25221), .B(n25222), .Z(n24694) );
  ANDN U32162 ( .B(n25223), .A(n25224), .Z(n25221) );
  AND U32163 ( .A(a[68]), .B(b[20]), .Z(n25220) );
  XOR U32164 ( .A(n25226), .B(n25227), .Z(n24699) );
  ANDN U32165 ( .B(n25228), .A(n25229), .Z(n25226) );
  AND U32166 ( .A(a[69]), .B(b[19]), .Z(n25225) );
  XOR U32167 ( .A(n25231), .B(n25232), .Z(n24704) );
  ANDN U32168 ( .B(n25233), .A(n25234), .Z(n25231) );
  AND U32169 ( .A(a[70]), .B(b[18]), .Z(n25230) );
  XOR U32170 ( .A(n25236), .B(n25237), .Z(n24709) );
  ANDN U32171 ( .B(n25238), .A(n25239), .Z(n25236) );
  AND U32172 ( .A(a[71]), .B(b[17]), .Z(n25235) );
  XOR U32173 ( .A(n25241), .B(n25242), .Z(n24714) );
  ANDN U32174 ( .B(n25243), .A(n25244), .Z(n25241) );
  AND U32175 ( .A(a[72]), .B(b[16]), .Z(n25240) );
  XOR U32176 ( .A(n25246), .B(n25247), .Z(n24719) );
  ANDN U32177 ( .B(n25248), .A(n25249), .Z(n25246) );
  AND U32178 ( .A(a[73]), .B(b[15]), .Z(n25245) );
  XOR U32179 ( .A(n25251), .B(n25252), .Z(n24724) );
  ANDN U32180 ( .B(n25253), .A(n25254), .Z(n25251) );
  AND U32181 ( .A(a[74]), .B(b[14]), .Z(n25250) );
  XOR U32182 ( .A(n25256), .B(n25257), .Z(n24729) );
  ANDN U32183 ( .B(n25258), .A(n25259), .Z(n25256) );
  AND U32184 ( .A(a[75]), .B(b[13]), .Z(n25255) );
  XOR U32185 ( .A(n25261), .B(n25262), .Z(n24734) );
  ANDN U32186 ( .B(n25263), .A(n25264), .Z(n25261) );
  AND U32187 ( .A(a[76]), .B(b[12]), .Z(n25260) );
  XOR U32188 ( .A(n25266), .B(n25267), .Z(n24739) );
  ANDN U32189 ( .B(n25268), .A(n25269), .Z(n25266) );
  AND U32190 ( .A(a[77]), .B(b[11]), .Z(n25265) );
  XOR U32191 ( .A(n25271), .B(n25272), .Z(n24744) );
  ANDN U32192 ( .B(n25273), .A(n25274), .Z(n25271) );
  AND U32193 ( .A(a[78]), .B(b[10]), .Z(n25270) );
  XOR U32194 ( .A(n25276), .B(n25277), .Z(n24749) );
  ANDN U32195 ( .B(n25278), .A(n25279), .Z(n25276) );
  AND U32196 ( .A(b[9]), .B(a[79]), .Z(n25275) );
  XOR U32197 ( .A(n25281), .B(n25282), .Z(n24754) );
  ANDN U32198 ( .B(n25283), .A(n25284), .Z(n25281) );
  AND U32199 ( .A(b[8]), .B(a[80]), .Z(n25280) );
  XOR U32200 ( .A(n25286), .B(n25287), .Z(n24759) );
  ANDN U32201 ( .B(n25288), .A(n25289), .Z(n25286) );
  AND U32202 ( .A(b[7]), .B(a[81]), .Z(n25285) );
  XOR U32203 ( .A(n25291), .B(n25292), .Z(n24764) );
  ANDN U32204 ( .B(n25293), .A(n25294), .Z(n25291) );
  AND U32205 ( .A(b[6]), .B(a[82]), .Z(n25290) );
  XOR U32206 ( .A(n25296), .B(n25297), .Z(n24769) );
  ANDN U32207 ( .B(n25298), .A(n25299), .Z(n25296) );
  AND U32208 ( .A(b[5]), .B(a[83]), .Z(n25295) );
  XOR U32209 ( .A(n25301), .B(n25302), .Z(n24774) );
  ANDN U32210 ( .B(n25303), .A(n25304), .Z(n25301) );
  AND U32211 ( .A(b[4]), .B(a[84]), .Z(n25300) );
  XOR U32212 ( .A(n25306), .B(n25307), .Z(n24779) );
  ANDN U32213 ( .B(n24791), .A(n24792), .Z(n25306) );
  AND U32214 ( .A(b[2]), .B(a[85]), .Z(n25308) );
  XNOR U32215 ( .A(n25303), .B(n25307), .Z(n25309) );
  XOR U32216 ( .A(n25310), .B(n25311), .Z(n25307) );
  OR U32217 ( .A(n24794), .B(n24795), .Z(n25311) );
  XNOR U32218 ( .A(n25313), .B(n25314), .Z(n25312) );
  XOR U32219 ( .A(n25313), .B(n25316), .Z(n24794) );
  NAND U32220 ( .A(b[1]), .B(a[85]), .Z(n25316) );
  IV U32221 ( .A(n25310), .Z(n25313) );
  NANDN U32222 ( .A(n33), .B(n34), .Z(n25310) );
  XOR U32223 ( .A(n25317), .B(n25318), .Z(n34) );
  NAND U32224 ( .A(a[85]), .B(b[0]), .Z(n33) );
  XNOR U32225 ( .A(n25298), .B(n25302), .Z(n25319) );
  XNOR U32226 ( .A(n25293), .B(n25297), .Z(n25320) );
  XNOR U32227 ( .A(n25288), .B(n25292), .Z(n25321) );
  XNOR U32228 ( .A(n25283), .B(n25287), .Z(n25322) );
  XNOR U32229 ( .A(n25278), .B(n25282), .Z(n25323) );
  XNOR U32230 ( .A(n25273), .B(n25277), .Z(n25324) );
  XNOR U32231 ( .A(n25268), .B(n25272), .Z(n25325) );
  XNOR U32232 ( .A(n25263), .B(n25267), .Z(n25326) );
  XNOR U32233 ( .A(n25258), .B(n25262), .Z(n25327) );
  XNOR U32234 ( .A(n25253), .B(n25257), .Z(n25328) );
  XNOR U32235 ( .A(n25248), .B(n25252), .Z(n25329) );
  XNOR U32236 ( .A(n25243), .B(n25247), .Z(n25330) );
  XNOR U32237 ( .A(n25238), .B(n25242), .Z(n25331) );
  XNOR U32238 ( .A(n25233), .B(n25237), .Z(n25332) );
  XNOR U32239 ( .A(n25228), .B(n25232), .Z(n25333) );
  XNOR U32240 ( .A(n25223), .B(n25227), .Z(n25334) );
  XNOR U32241 ( .A(n25218), .B(n25222), .Z(n25335) );
  XNOR U32242 ( .A(n25213), .B(n25217), .Z(n25336) );
  XNOR U32243 ( .A(n25208), .B(n25212), .Z(n25337) );
  XNOR U32244 ( .A(n25203), .B(n25207), .Z(n25338) );
  XNOR U32245 ( .A(n25198), .B(n25202), .Z(n25339) );
  XNOR U32246 ( .A(n25193), .B(n25197), .Z(n25340) );
  XNOR U32247 ( .A(n25188), .B(n25192), .Z(n25341) );
  XNOR U32248 ( .A(n25183), .B(n25187), .Z(n25342) );
  XNOR U32249 ( .A(n25178), .B(n25182), .Z(n25343) );
  XNOR U32250 ( .A(n25173), .B(n25177), .Z(n25344) );
  XNOR U32251 ( .A(n25168), .B(n25172), .Z(n25345) );
  XNOR U32252 ( .A(n25163), .B(n25167), .Z(n25346) );
  XNOR U32253 ( .A(n25158), .B(n25162), .Z(n25347) );
  XNOR U32254 ( .A(n25153), .B(n25157), .Z(n25348) );
  XNOR U32255 ( .A(n25148), .B(n25152), .Z(n25349) );
  XNOR U32256 ( .A(n25143), .B(n25147), .Z(n25350) );
  XNOR U32257 ( .A(n25138), .B(n25142), .Z(n25351) );
  XNOR U32258 ( .A(n25133), .B(n25137), .Z(n25352) );
  XNOR U32259 ( .A(n25128), .B(n25132), .Z(n25353) );
  XNOR U32260 ( .A(n25123), .B(n25127), .Z(n25354) );
  XNOR U32261 ( .A(n25118), .B(n25122), .Z(n25355) );
  XNOR U32262 ( .A(n25113), .B(n25117), .Z(n25356) );
  XNOR U32263 ( .A(n25108), .B(n25112), .Z(n25357) );
  XNOR U32264 ( .A(n25103), .B(n25107), .Z(n25358) );
  XNOR U32265 ( .A(n25098), .B(n25102), .Z(n25359) );
  XNOR U32266 ( .A(n25093), .B(n25097), .Z(n25360) );
  XNOR U32267 ( .A(n25088), .B(n25092), .Z(n25361) );
  XNOR U32268 ( .A(n25083), .B(n25087), .Z(n25362) );
  XNOR U32269 ( .A(n25078), .B(n25082), .Z(n25363) );
  XNOR U32270 ( .A(n25073), .B(n25077), .Z(n25364) );
  XNOR U32271 ( .A(n25068), .B(n25072), .Z(n25365) );
  XNOR U32272 ( .A(n25063), .B(n25067), .Z(n25366) );
  XNOR U32273 ( .A(n25058), .B(n25062), .Z(n25367) );
  XNOR U32274 ( .A(n25053), .B(n25057), .Z(n25368) );
  XNOR U32275 ( .A(n25048), .B(n25052), .Z(n25369) );
  XNOR U32276 ( .A(n25043), .B(n25047), .Z(n25370) );
  XNOR U32277 ( .A(n25038), .B(n25042), .Z(n25371) );
  XNOR U32278 ( .A(n25033), .B(n25037), .Z(n25372) );
  XNOR U32279 ( .A(n25028), .B(n25032), .Z(n25373) );
  XNOR U32280 ( .A(n25023), .B(n25027), .Z(n25374) );
  XNOR U32281 ( .A(n25018), .B(n25022), .Z(n25375) );
  XNOR U32282 ( .A(n25013), .B(n25017), .Z(n25376) );
  XNOR U32283 ( .A(n25008), .B(n25012), .Z(n25377) );
  XNOR U32284 ( .A(n25003), .B(n25007), .Z(n25378) );
  XNOR U32285 ( .A(n24998), .B(n25002), .Z(n25379) );
  XNOR U32286 ( .A(n24993), .B(n24997), .Z(n25380) );
  XNOR U32287 ( .A(n24987), .B(n24992), .Z(n25381) );
  XNOR U32288 ( .A(n24982), .B(n24986), .Z(n25382) );
  XNOR U32289 ( .A(n24977), .B(n24981), .Z(n25383) );
  XNOR U32290 ( .A(n24972), .B(n24976), .Z(n25384) );
  XNOR U32291 ( .A(n24967), .B(n24971), .Z(n25385) );
  XNOR U32292 ( .A(n24962), .B(n24966), .Z(n25386) );
  XNOR U32293 ( .A(n25387), .B(n25388), .Z(n24962) );
  XNOR U32294 ( .A(n24957), .B(n24961), .Z(n25388) );
  XNOR U32295 ( .A(n24952), .B(n24956), .Z(n25389) );
  XNOR U32296 ( .A(n24947), .B(n24951), .Z(n25390) );
  XNOR U32297 ( .A(n24942), .B(n24946), .Z(n25391) );
  XNOR U32298 ( .A(n24937), .B(n24941), .Z(n25392) );
  XNOR U32299 ( .A(n24932), .B(n24936), .Z(n25393) );
  XNOR U32300 ( .A(n24927), .B(n24931), .Z(n25394) );
  XNOR U32301 ( .A(n24922), .B(n24926), .Z(n25395) );
  XNOR U32302 ( .A(n24917), .B(n24921), .Z(n25396) );
  XNOR U32303 ( .A(n24912), .B(n24916), .Z(n25397) );
  XNOR U32304 ( .A(n24907), .B(n24911), .Z(n25398) );
  XNOR U32305 ( .A(n24902), .B(n24906), .Z(n25399) );
  XNOR U32306 ( .A(n24897), .B(n24901), .Z(n25400) );
  XNOR U32307 ( .A(n24892), .B(n24896), .Z(n25401) );
  XNOR U32308 ( .A(n24887), .B(n24891), .Z(n25402) );
  XNOR U32309 ( .A(n25403), .B(n24886), .Z(n24887) );
  AND U32310 ( .A(a[0]), .B(b[87]), .Z(n25403) );
  XOR U32311 ( .A(n25404), .B(n24886), .Z(n24888) );
  XNOR U32312 ( .A(n25405), .B(n25406), .Z(n24886) );
  ANDN U32313 ( .B(n25407), .A(n25408), .Z(n25405) );
  AND U32314 ( .A(a[1]), .B(b[86]), .Z(n25404) );
  XOR U32315 ( .A(n25410), .B(n25411), .Z(n24891) );
  ANDN U32316 ( .B(n25412), .A(n25413), .Z(n25410) );
  AND U32317 ( .A(a[2]), .B(b[85]), .Z(n25409) );
  XOR U32318 ( .A(n25415), .B(n25416), .Z(n24896) );
  ANDN U32319 ( .B(n25417), .A(n25418), .Z(n25415) );
  AND U32320 ( .A(a[3]), .B(b[84]), .Z(n25414) );
  XOR U32321 ( .A(n25420), .B(n25421), .Z(n24901) );
  ANDN U32322 ( .B(n25422), .A(n25423), .Z(n25420) );
  AND U32323 ( .A(a[4]), .B(b[83]), .Z(n25419) );
  XOR U32324 ( .A(n25425), .B(n25426), .Z(n24906) );
  ANDN U32325 ( .B(n25427), .A(n25428), .Z(n25425) );
  AND U32326 ( .A(a[5]), .B(b[82]), .Z(n25424) );
  XOR U32327 ( .A(n25430), .B(n25431), .Z(n24911) );
  ANDN U32328 ( .B(n25432), .A(n25433), .Z(n25430) );
  AND U32329 ( .A(a[6]), .B(b[81]), .Z(n25429) );
  XOR U32330 ( .A(n25435), .B(n25436), .Z(n24916) );
  ANDN U32331 ( .B(n25437), .A(n25438), .Z(n25435) );
  AND U32332 ( .A(a[7]), .B(b[80]), .Z(n25434) );
  XOR U32333 ( .A(n25440), .B(n25441), .Z(n24921) );
  ANDN U32334 ( .B(n25442), .A(n25443), .Z(n25440) );
  AND U32335 ( .A(a[8]), .B(b[79]), .Z(n25439) );
  XOR U32336 ( .A(n25445), .B(n25446), .Z(n24926) );
  ANDN U32337 ( .B(n25447), .A(n25448), .Z(n25445) );
  AND U32338 ( .A(a[9]), .B(b[78]), .Z(n25444) );
  XOR U32339 ( .A(n25450), .B(n25451), .Z(n24931) );
  ANDN U32340 ( .B(n25452), .A(n25453), .Z(n25450) );
  AND U32341 ( .A(a[10]), .B(b[77]), .Z(n25449) );
  XOR U32342 ( .A(n25455), .B(n25456), .Z(n24936) );
  ANDN U32343 ( .B(n25457), .A(n25458), .Z(n25455) );
  AND U32344 ( .A(a[11]), .B(b[76]), .Z(n25454) );
  XOR U32345 ( .A(n25460), .B(n25461), .Z(n24941) );
  ANDN U32346 ( .B(n25462), .A(n25463), .Z(n25460) );
  AND U32347 ( .A(a[12]), .B(b[75]), .Z(n25459) );
  XOR U32348 ( .A(n25465), .B(n25466), .Z(n24946) );
  ANDN U32349 ( .B(n25467), .A(n25468), .Z(n25465) );
  AND U32350 ( .A(a[13]), .B(b[74]), .Z(n25464) );
  XOR U32351 ( .A(n25470), .B(n25471), .Z(n24951) );
  ANDN U32352 ( .B(n25472), .A(n25473), .Z(n25470) );
  AND U32353 ( .A(a[14]), .B(b[73]), .Z(n25469) );
  IV U32354 ( .A(n24958), .Z(n25387) );
  XOR U32355 ( .A(n25475), .B(n25476), .Z(n24956) );
  ANDN U32356 ( .B(n25477), .A(n25478), .Z(n25475) );
  AND U32357 ( .A(a[15]), .B(b[72]), .Z(n25474) );
  XOR U32358 ( .A(n25480), .B(n25481), .Z(n24961) );
  ANDN U32359 ( .B(n25482), .A(n25483), .Z(n25480) );
  AND U32360 ( .A(a[16]), .B(b[71]), .Z(n25479) );
  XOR U32361 ( .A(n25485), .B(n25486), .Z(n24966) );
  ANDN U32362 ( .B(n25487), .A(n25488), .Z(n25485) );
  AND U32363 ( .A(a[17]), .B(b[70]), .Z(n25484) );
  XOR U32364 ( .A(n25490), .B(n25491), .Z(n24971) );
  ANDN U32365 ( .B(n25492), .A(n25493), .Z(n25490) );
  AND U32366 ( .A(a[18]), .B(b[69]), .Z(n25489) );
  XOR U32367 ( .A(n25495), .B(n25496), .Z(n24976) );
  ANDN U32368 ( .B(n25497), .A(n25498), .Z(n25495) );
  AND U32369 ( .A(a[19]), .B(b[68]), .Z(n25494) );
  XOR U32370 ( .A(n25500), .B(n25501), .Z(n24981) );
  ANDN U32371 ( .B(n25502), .A(n25503), .Z(n25500) );
  AND U32372 ( .A(a[20]), .B(b[67]), .Z(n25499) );
  XOR U32373 ( .A(n25505), .B(n25506), .Z(n24986) );
  ANDN U32374 ( .B(n25507), .A(n25508), .Z(n25505) );
  AND U32375 ( .A(a[21]), .B(b[66]), .Z(n25504) );
  XOR U32376 ( .A(n25510), .B(n25511), .Z(n24992) );
  ANDN U32377 ( .B(n25512), .A(n25513), .Z(n25510) );
  AND U32378 ( .A(a[22]), .B(b[65]), .Z(n25509) );
  XOR U32379 ( .A(n25515), .B(n25516), .Z(n24997) );
  ANDN U32380 ( .B(n25517), .A(n25518), .Z(n25515) );
  AND U32381 ( .A(a[23]), .B(b[64]), .Z(n25514) );
  XOR U32382 ( .A(n25520), .B(n25521), .Z(n25002) );
  ANDN U32383 ( .B(n25522), .A(n25523), .Z(n25520) );
  AND U32384 ( .A(a[24]), .B(b[63]), .Z(n25519) );
  XOR U32385 ( .A(n25525), .B(n25526), .Z(n25007) );
  ANDN U32386 ( .B(n25527), .A(n25528), .Z(n25525) );
  AND U32387 ( .A(a[25]), .B(b[62]), .Z(n25524) );
  XOR U32388 ( .A(n25530), .B(n25531), .Z(n25012) );
  ANDN U32389 ( .B(n25532), .A(n25533), .Z(n25530) );
  AND U32390 ( .A(a[26]), .B(b[61]), .Z(n25529) );
  XOR U32391 ( .A(n25535), .B(n25536), .Z(n25017) );
  ANDN U32392 ( .B(n25537), .A(n25538), .Z(n25535) );
  AND U32393 ( .A(a[27]), .B(b[60]), .Z(n25534) );
  XOR U32394 ( .A(n25540), .B(n25541), .Z(n25022) );
  ANDN U32395 ( .B(n25542), .A(n25543), .Z(n25540) );
  AND U32396 ( .A(a[28]), .B(b[59]), .Z(n25539) );
  XOR U32397 ( .A(n25545), .B(n25546), .Z(n25027) );
  ANDN U32398 ( .B(n25547), .A(n25548), .Z(n25545) );
  AND U32399 ( .A(a[29]), .B(b[58]), .Z(n25544) );
  XOR U32400 ( .A(n25550), .B(n25551), .Z(n25032) );
  ANDN U32401 ( .B(n25552), .A(n25553), .Z(n25550) );
  AND U32402 ( .A(a[30]), .B(b[57]), .Z(n25549) );
  XOR U32403 ( .A(n25555), .B(n25556), .Z(n25037) );
  ANDN U32404 ( .B(n25557), .A(n25558), .Z(n25555) );
  AND U32405 ( .A(a[31]), .B(b[56]), .Z(n25554) );
  XOR U32406 ( .A(n25560), .B(n25561), .Z(n25042) );
  ANDN U32407 ( .B(n25562), .A(n25563), .Z(n25560) );
  AND U32408 ( .A(a[32]), .B(b[55]), .Z(n25559) );
  XOR U32409 ( .A(n25565), .B(n25566), .Z(n25047) );
  ANDN U32410 ( .B(n25567), .A(n25568), .Z(n25565) );
  AND U32411 ( .A(a[33]), .B(b[54]), .Z(n25564) );
  XOR U32412 ( .A(n25570), .B(n25571), .Z(n25052) );
  ANDN U32413 ( .B(n25572), .A(n25573), .Z(n25570) );
  AND U32414 ( .A(a[34]), .B(b[53]), .Z(n25569) );
  XOR U32415 ( .A(n25575), .B(n25576), .Z(n25057) );
  ANDN U32416 ( .B(n25577), .A(n25578), .Z(n25575) );
  AND U32417 ( .A(a[35]), .B(b[52]), .Z(n25574) );
  XOR U32418 ( .A(n25580), .B(n25581), .Z(n25062) );
  ANDN U32419 ( .B(n25582), .A(n25583), .Z(n25580) );
  AND U32420 ( .A(a[36]), .B(b[51]), .Z(n25579) );
  XOR U32421 ( .A(n25585), .B(n25586), .Z(n25067) );
  ANDN U32422 ( .B(n25587), .A(n25588), .Z(n25585) );
  AND U32423 ( .A(a[37]), .B(b[50]), .Z(n25584) );
  XOR U32424 ( .A(n25590), .B(n25591), .Z(n25072) );
  ANDN U32425 ( .B(n25592), .A(n25593), .Z(n25590) );
  AND U32426 ( .A(a[38]), .B(b[49]), .Z(n25589) );
  XOR U32427 ( .A(n25595), .B(n25596), .Z(n25077) );
  ANDN U32428 ( .B(n25597), .A(n25598), .Z(n25595) );
  AND U32429 ( .A(a[39]), .B(b[48]), .Z(n25594) );
  XOR U32430 ( .A(n25600), .B(n25601), .Z(n25082) );
  ANDN U32431 ( .B(n25602), .A(n25603), .Z(n25600) );
  AND U32432 ( .A(a[40]), .B(b[47]), .Z(n25599) );
  XOR U32433 ( .A(n25605), .B(n25606), .Z(n25087) );
  ANDN U32434 ( .B(n25607), .A(n25608), .Z(n25605) );
  AND U32435 ( .A(a[41]), .B(b[46]), .Z(n25604) );
  XOR U32436 ( .A(n25610), .B(n25611), .Z(n25092) );
  ANDN U32437 ( .B(n25612), .A(n25613), .Z(n25610) );
  AND U32438 ( .A(a[42]), .B(b[45]), .Z(n25609) );
  XOR U32439 ( .A(n25615), .B(n25616), .Z(n25097) );
  ANDN U32440 ( .B(n25617), .A(n25618), .Z(n25615) );
  AND U32441 ( .A(a[43]), .B(b[44]), .Z(n25614) );
  XOR U32442 ( .A(n25620), .B(n25621), .Z(n25102) );
  ANDN U32443 ( .B(n25622), .A(n25623), .Z(n25620) );
  AND U32444 ( .A(a[44]), .B(b[43]), .Z(n25619) );
  XOR U32445 ( .A(n25625), .B(n25626), .Z(n25107) );
  ANDN U32446 ( .B(n25627), .A(n25628), .Z(n25625) );
  AND U32447 ( .A(a[45]), .B(b[42]), .Z(n25624) );
  XOR U32448 ( .A(n25630), .B(n25631), .Z(n25112) );
  ANDN U32449 ( .B(n25632), .A(n25633), .Z(n25630) );
  AND U32450 ( .A(a[46]), .B(b[41]), .Z(n25629) );
  XOR U32451 ( .A(n25635), .B(n25636), .Z(n25117) );
  ANDN U32452 ( .B(n25637), .A(n25638), .Z(n25635) );
  AND U32453 ( .A(a[47]), .B(b[40]), .Z(n25634) );
  XOR U32454 ( .A(n25640), .B(n25641), .Z(n25122) );
  ANDN U32455 ( .B(n25642), .A(n25643), .Z(n25640) );
  AND U32456 ( .A(a[48]), .B(b[39]), .Z(n25639) );
  XOR U32457 ( .A(n25645), .B(n25646), .Z(n25127) );
  ANDN U32458 ( .B(n25647), .A(n25648), .Z(n25645) );
  AND U32459 ( .A(a[49]), .B(b[38]), .Z(n25644) );
  XOR U32460 ( .A(n25650), .B(n25651), .Z(n25132) );
  ANDN U32461 ( .B(n25652), .A(n25653), .Z(n25650) );
  AND U32462 ( .A(a[50]), .B(b[37]), .Z(n25649) );
  XOR U32463 ( .A(n25655), .B(n25656), .Z(n25137) );
  ANDN U32464 ( .B(n25657), .A(n25658), .Z(n25655) );
  AND U32465 ( .A(a[51]), .B(b[36]), .Z(n25654) );
  XOR U32466 ( .A(n25660), .B(n25661), .Z(n25142) );
  ANDN U32467 ( .B(n25662), .A(n25663), .Z(n25660) );
  AND U32468 ( .A(a[52]), .B(b[35]), .Z(n25659) );
  XOR U32469 ( .A(n25665), .B(n25666), .Z(n25147) );
  ANDN U32470 ( .B(n25667), .A(n25668), .Z(n25665) );
  AND U32471 ( .A(a[53]), .B(b[34]), .Z(n25664) );
  XOR U32472 ( .A(n25670), .B(n25671), .Z(n25152) );
  ANDN U32473 ( .B(n25672), .A(n25673), .Z(n25670) );
  AND U32474 ( .A(a[54]), .B(b[33]), .Z(n25669) );
  XOR U32475 ( .A(n25675), .B(n25676), .Z(n25157) );
  ANDN U32476 ( .B(n25677), .A(n25678), .Z(n25675) );
  AND U32477 ( .A(a[55]), .B(b[32]), .Z(n25674) );
  XOR U32478 ( .A(n25680), .B(n25681), .Z(n25162) );
  ANDN U32479 ( .B(n25682), .A(n25683), .Z(n25680) );
  AND U32480 ( .A(a[56]), .B(b[31]), .Z(n25679) );
  XOR U32481 ( .A(n25685), .B(n25686), .Z(n25167) );
  ANDN U32482 ( .B(n25687), .A(n25688), .Z(n25685) );
  AND U32483 ( .A(a[57]), .B(b[30]), .Z(n25684) );
  XOR U32484 ( .A(n25690), .B(n25691), .Z(n25172) );
  ANDN U32485 ( .B(n25692), .A(n25693), .Z(n25690) );
  AND U32486 ( .A(a[58]), .B(b[29]), .Z(n25689) );
  XOR U32487 ( .A(n25695), .B(n25696), .Z(n25177) );
  ANDN U32488 ( .B(n25697), .A(n25698), .Z(n25695) );
  AND U32489 ( .A(a[59]), .B(b[28]), .Z(n25694) );
  XOR U32490 ( .A(n25700), .B(n25701), .Z(n25182) );
  ANDN U32491 ( .B(n25702), .A(n25703), .Z(n25700) );
  AND U32492 ( .A(a[60]), .B(b[27]), .Z(n25699) );
  XOR U32493 ( .A(n25705), .B(n25706), .Z(n25187) );
  ANDN U32494 ( .B(n25707), .A(n25708), .Z(n25705) );
  AND U32495 ( .A(a[61]), .B(b[26]), .Z(n25704) );
  XOR U32496 ( .A(n25710), .B(n25711), .Z(n25192) );
  ANDN U32497 ( .B(n25712), .A(n25713), .Z(n25710) );
  AND U32498 ( .A(a[62]), .B(b[25]), .Z(n25709) );
  XOR U32499 ( .A(n25715), .B(n25716), .Z(n25197) );
  ANDN U32500 ( .B(n25717), .A(n25718), .Z(n25715) );
  AND U32501 ( .A(a[63]), .B(b[24]), .Z(n25714) );
  XOR U32502 ( .A(n25720), .B(n25721), .Z(n25202) );
  ANDN U32503 ( .B(n25722), .A(n25723), .Z(n25720) );
  AND U32504 ( .A(a[64]), .B(b[23]), .Z(n25719) );
  XOR U32505 ( .A(n25725), .B(n25726), .Z(n25207) );
  ANDN U32506 ( .B(n25727), .A(n25728), .Z(n25725) );
  AND U32507 ( .A(a[65]), .B(b[22]), .Z(n25724) );
  XOR U32508 ( .A(n25730), .B(n25731), .Z(n25212) );
  ANDN U32509 ( .B(n25732), .A(n25733), .Z(n25730) );
  AND U32510 ( .A(a[66]), .B(b[21]), .Z(n25729) );
  XOR U32511 ( .A(n25735), .B(n25736), .Z(n25217) );
  ANDN U32512 ( .B(n25737), .A(n25738), .Z(n25735) );
  AND U32513 ( .A(a[67]), .B(b[20]), .Z(n25734) );
  XOR U32514 ( .A(n25740), .B(n25741), .Z(n25222) );
  ANDN U32515 ( .B(n25742), .A(n25743), .Z(n25740) );
  AND U32516 ( .A(a[68]), .B(b[19]), .Z(n25739) );
  XOR U32517 ( .A(n25745), .B(n25746), .Z(n25227) );
  ANDN U32518 ( .B(n25747), .A(n25748), .Z(n25745) );
  AND U32519 ( .A(a[69]), .B(b[18]), .Z(n25744) );
  XOR U32520 ( .A(n25750), .B(n25751), .Z(n25232) );
  ANDN U32521 ( .B(n25752), .A(n25753), .Z(n25750) );
  AND U32522 ( .A(a[70]), .B(b[17]), .Z(n25749) );
  XOR U32523 ( .A(n25755), .B(n25756), .Z(n25237) );
  ANDN U32524 ( .B(n25757), .A(n25758), .Z(n25755) );
  AND U32525 ( .A(a[71]), .B(b[16]), .Z(n25754) );
  XOR U32526 ( .A(n25760), .B(n25761), .Z(n25242) );
  ANDN U32527 ( .B(n25762), .A(n25763), .Z(n25760) );
  AND U32528 ( .A(a[72]), .B(b[15]), .Z(n25759) );
  XOR U32529 ( .A(n25765), .B(n25766), .Z(n25247) );
  ANDN U32530 ( .B(n25767), .A(n25768), .Z(n25765) );
  AND U32531 ( .A(a[73]), .B(b[14]), .Z(n25764) );
  XOR U32532 ( .A(n25770), .B(n25771), .Z(n25252) );
  ANDN U32533 ( .B(n25772), .A(n25773), .Z(n25770) );
  AND U32534 ( .A(a[74]), .B(b[13]), .Z(n25769) );
  XOR U32535 ( .A(n25775), .B(n25776), .Z(n25257) );
  ANDN U32536 ( .B(n25777), .A(n25778), .Z(n25775) );
  AND U32537 ( .A(a[75]), .B(b[12]), .Z(n25774) );
  XOR U32538 ( .A(n25780), .B(n25781), .Z(n25262) );
  ANDN U32539 ( .B(n25782), .A(n25783), .Z(n25780) );
  AND U32540 ( .A(a[76]), .B(b[11]), .Z(n25779) );
  XOR U32541 ( .A(n25785), .B(n25786), .Z(n25267) );
  ANDN U32542 ( .B(n25787), .A(n25788), .Z(n25785) );
  AND U32543 ( .A(a[77]), .B(b[10]), .Z(n25784) );
  XOR U32544 ( .A(n25790), .B(n25791), .Z(n25272) );
  ANDN U32545 ( .B(n25792), .A(n25793), .Z(n25790) );
  AND U32546 ( .A(b[9]), .B(a[78]), .Z(n25789) );
  XOR U32547 ( .A(n25795), .B(n25796), .Z(n25277) );
  ANDN U32548 ( .B(n25797), .A(n25798), .Z(n25795) );
  AND U32549 ( .A(b[8]), .B(a[79]), .Z(n25794) );
  XOR U32550 ( .A(n25800), .B(n25801), .Z(n25282) );
  ANDN U32551 ( .B(n25802), .A(n25803), .Z(n25800) );
  AND U32552 ( .A(b[7]), .B(a[80]), .Z(n25799) );
  XOR U32553 ( .A(n25805), .B(n25806), .Z(n25287) );
  ANDN U32554 ( .B(n25807), .A(n25808), .Z(n25805) );
  AND U32555 ( .A(b[6]), .B(a[81]), .Z(n25804) );
  XOR U32556 ( .A(n25810), .B(n25811), .Z(n25292) );
  ANDN U32557 ( .B(n25812), .A(n25813), .Z(n25810) );
  AND U32558 ( .A(b[5]), .B(a[82]), .Z(n25809) );
  XOR U32559 ( .A(n25815), .B(n25816), .Z(n25297) );
  ANDN U32560 ( .B(n25817), .A(n25818), .Z(n25815) );
  AND U32561 ( .A(b[4]), .B(a[83]), .Z(n25814) );
  XOR U32562 ( .A(n25820), .B(n25821), .Z(n25302) );
  ANDN U32563 ( .B(n25314), .A(n25315), .Z(n25820) );
  AND U32564 ( .A(b[2]), .B(a[84]), .Z(n25822) );
  XNOR U32565 ( .A(n25817), .B(n25821), .Z(n25823) );
  XOR U32566 ( .A(n25824), .B(n25825), .Z(n25821) );
  OR U32567 ( .A(n25317), .B(n25318), .Z(n25825) );
  XNOR U32568 ( .A(n25827), .B(n25828), .Z(n25826) );
  XOR U32569 ( .A(n25827), .B(n25830), .Z(n25317) );
  NAND U32570 ( .A(b[1]), .B(a[84]), .Z(n25830) );
  IV U32571 ( .A(n25824), .Z(n25827) );
  NANDN U32572 ( .A(n35), .B(n36), .Z(n25824) );
  XOR U32573 ( .A(n25831), .B(n25832), .Z(n36) );
  NAND U32574 ( .A(a[84]), .B(b[0]), .Z(n35) );
  XNOR U32575 ( .A(n25812), .B(n25816), .Z(n25833) );
  XNOR U32576 ( .A(n25807), .B(n25811), .Z(n25834) );
  XNOR U32577 ( .A(n25802), .B(n25806), .Z(n25835) );
  XNOR U32578 ( .A(n25797), .B(n25801), .Z(n25836) );
  XNOR U32579 ( .A(n25792), .B(n25796), .Z(n25837) );
  XNOR U32580 ( .A(n25787), .B(n25791), .Z(n25838) );
  XNOR U32581 ( .A(n25782), .B(n25786), .Z(n25839) );
  XNOR U32582 ( .A(n25777), .B(n25781), .Z(n25840) );
  XNOR U32583 ( .A(n25772), .B(n25776), .Z(n25841) );
  XNOR U32584 ( .A(n25767), .B(n25771), .Z(n25842) );
  XNOR U32585 ( .A(n25762), .B(n25766), .Z(n25843) );
  XNOR U32586 ( .A(n25757), .B(n25761), .Z(n25844) );
  XNOR U32587 ( .A(n25752), .B(n25756), .Z(n25845) );
  XNOR U32588 ( .A(n25747), .B(n25751), .Z(n25846) );
  XNOR U32589 ( .A(n25742), .B(n25746), .Z(n25847) );
  XNOR U32590 ( .A(n25737), .B(n25741), .Z(n25848) );
  XNOR U32591 ( .A(n25732), .B(n25736), .Z(n25849) );
  XNOR U32592 ( .A(n25727), .B(n25731), .Z(n25850) );
  XNOR U32593 ( .A(n25722), .B(n25726), .Z(n25851) );
  XNOR U32594 ( .A(n25717), .B(n25721), .Z(n25852) );
  XNOR U32595 ( .A(n25712), .B(n25716), .Z(n25853) );
  XNOR U32596 ( .A(n25707), .B(n25711), .Z(n25854) );
  XNOR U32597 ( .A(n25702), .B(n25706), .Z(n25855) );
  XNOR U32598 ( .A(n25697), .B(n25701), .Z(n25856) );
  XNOR U32599 ( .A(n25692), .B(n25696), .Z(n25857) );
  XNOR U32600 ( .A(n25687), .B(n25691), .Z(n25858) );
  XNOR U32601 ( .A(n25682), .B(n25686), .Z(n25859) );
  XNOR U32602 ( .A(n25677), .B(n25681), .Z(n25860) );
  XNOR U32603 ( .A(n25672), .B(n25676), .Z(n25861) );
  XNOR U32604 ( .A(n25667), .B(n25671), .Z(n25862) );
  XNOR U32605 ( .A(n25662), .B(n25666), .Z(n25863) );
  XNOR U32606 ( .A(n25657), .B(n25661), .Z(n25864) );
  XNOR U32607 ( .A(n25652), .B(n25656), .Z(n25865) );
  XNOR U32608 ( .A(n25647), .B(n25651), .Z(n25866) );
  XNOR U32609 ( .A(n25642), .B(n25646), .Z(n25867) );
  XNOR U32610 ( .A(n25637), .B(n25641), .Z(n25868) );
  XNOR U32611 ( .A(n25632), .B(n25636), .Z(n25869) );
  XNOR U32612 ( .A(n25627), .B(n25631), .Z(n25870) );
  XNOR U32613 ( .A(n25622), .B(n25626), .Z(n25871) );
  XNOR U32614 ( .A(n25617), .B(n25621), .Z(n25872) );
  XNOR U32615 ( .A(n25612), .B(n25616), .Z(n25873) );
  XNOR U32616 ( .A(n25607), .B(n25611), .Z(n25874) );
  XNOR U32617 ( .A(n25602), .B(n25606), .Z(n25875) );
  XNOR U32618 ( .A(n25597), .B(n25601), .Z(n25876) );
  XNOR U32619 ( .A(n25592), .B(n25596), .Z(n25877) );
  XNOR U32620 ( .A(n25587), .B(n25591), .Z(n25878) );
  XNOR U32621 ( .A(n25582), .B(n25586), .Z(n25879) );
  XNOR U32622 ( .A(n25577), .B(n25581), .Z(n25880) );
  XNOR U32623 ( .A(n25572), .B(n25576), .Z(n25881) );
  XNOR U32624 ( .A(n25567), .B(n25571), .Z(n25882) );
  XNOR U32625 ( .A(n25562), .B(n25566), .Z(n25883) );
  XNOR U32626 ( .A(n25557), .B(n25561), .Z(n25884) );
  XNOR U32627 ( .A(n25552), .B(n25556), .Z(n25885) );
  XNOR U32628 ( .A(n25547), .B(n25551), .Z(n25886) );
  XNOR U32629 ( .A(n25542), .B(n25546), .Z(n25887) );
  XNOR U32630 ( .A(n25537), .B(n25541), .Z(n25888) );
  XNOR U32631 ( .A(n25532), .B(n25536), .Z(n25889) );
  XNOR U32632 ( .A(n25527), .B(n25531), .Z(n25890) );
  XNOR U32633 ( .A(n25522), .B(n25526), .Z(n25891) );
  XNOR U32634 ( .A(n25517), .B(n25521), .Z(n25892) );
  XNOR U32635 ( .A(n25512), .B(n25516), .Z(n25893) );
  XNOR U32636 ( .A(n25507), .B(n25511), .Z(n25894) );
  XNOR U32637 ( .A(n25502), .B(n25506), .Z(n25895) );
  XNOR U32638 ( .A(n25497), .B(n25501), .Z(n25896) );
  XNOR U32639 ( .A(n25492), .B(n25496), .Z(n25897) );
  XNOR U32640 ( .A(n25487), .B(n25491), .Z(n25898) );
  XNOR U32641 ( .A(n25482), .B(n25486), .Z(n25899) );
  XNOR U32642 ( .A(n25477), .B(n25481), .Z(n25900) );
  XNOR U32643 ( .A(n25472), .B(n25476), .Z(n25901) );
  XNOR U32644 ( .A(n25902), .B(n25903), .Z(n25472) );
  XNOR U32645 ( .A(n25467), .B(n25471), .Z(n25903) );
  XNOR U32646 ( .A(n25462), .B(n25466), .Z(n25904) );
  XNOR U32647 ( .A(n25457), .B(n25461), .Z(n25905) );
  XNOR U32648 ( .A(n25452), .B(n25456), .Z(n25906) );
  XNOR U32649 ( .A(n25447), .B(n25451), .Z(n25907) );
  XNOR U32650 ( .A(n25442), .B(n25446), .Z(n25908) );
  XNOR U32651 ( .A(n25437), .B(n25441), .Z(n25909) );
  XNOR U32652 ( .A(n25432), .B(n25436), .Z(n25910) );
  XNOR U32653 ( .A(n25427), .B(n25431), .Z(n25911) );
  XNOR U32654 ( .A(n25422), .B(n25426), .Z(n25912) );
  XNOR U32655 ( .A(n25417), .B(n25421), .Z(n25913) );
  XNOR U32656 ( .A(n25412), .B(n25416), .Z(n25914) );
  XNOR U32657 ( .A(n25407), .B(n25411), .Z(n25915) );
  XOR U32658 ( .A(n25916), .B(n25406), .Z(n25407) );
  AND U32659 ( .A(a[0]), .B(b[86]), .Z(n25916) );
  XNOR U32660 ( .A(n25917), .B(n25406), .Z(n25408) );
  XNOR U32661 ( .A(n25918), .B(n25919), .Z(n25406) );
  ANDN U32662 ( .B(n25920), .A(n25921), .Z(n25918) );
  AND U32663 ( .A(a[1]), .B(b[85]), .Z(n25917) );
  XOR U32664 ( .A(n25923), .B(n25924), .Z(n25411) );
  ANDN U32665 ( .B(n25925), .A(n25926), .Z(n25923) );
  AND U32666 ( .A(a[2]), .B(b[84]), .Z(n25922) );
  XOR U32667 ( .A(n25928), .B(n25929), .Z(n25416) );
  ANDN U32668 ( .B(n25930), .A(n25931), .Z(n25928) );
  AND U32669 ( .A(a[3]), .B(b[83]), .Z(n25927) );
  XOR U32670 ( .A(n25933), .B(n25934), .Z(n25421) );
  ANDN U32671 ( .B(n25935), .A(n25936), .Z(n25933) );
  AND U32672 ( .A(a[4]), .B(b[82]), .Z(n25932) );
  XOR U32673 ( .A(n25938), .B(n25939), .Z(n25426) );
  ANDN U32674 ( .B(n25940), .A(n25941), .Z(n25938) );
  AND U32675 ( .A(a[5]), .B(b[81]), .Z(n25937) );
  XOR U32676 ( .A(n25943), .B(n25944), .Z(n25431) );
  ANDN U32677 ( .B(n25945), .A(n25946), .Z(n25943) );
  AND U32678 ( .A(a[6]), .B(b[80]), .Z(n25942) );
  XOR U32679 ( .A(n25948), .B(n25949), .Z(n25436) );
  ANDN U32680 ( .B(n25950), .A(n25951), .Z(n25948) );
  AND U32681 ( .A(a[7]), .B(b[79]), .Z(n25947) );
  XOR U32682 ( .A(n25953), .B(n25954), .Z(n25441) );
  ANDN U32683 ( .B(n25955), .A(n25956), .Z(n25953) );
  AND U32684 ( .A(a[8]), .B(b[78]), .Z(n25952) );
  XOR U32685 ( .A(n25958), .B(n25959), .Z(n25446) );
  ANDN U32686 ( .B(n25960), .A(n25961), .Z(n25958) );
  AND U32687 ( .A(a[9]), .B(b[77]), .Z(n25957) );
  XOR U32688 ( .A(n25963), .B(n25964), .Z(n25451) );
  ANDN U32689 ( .B(n25965), .A(n25966), .Z(n25963) );
  AND U32690 ( .A(a[10]), .B(b[76]), .Z(n25962) );
  XOR U32691 ( .A(n25968), .B(n25969), .Z(n25456) );
  ANDN U32692 ( .B(n25970), .A(n25971), .Z(n25968) );
  AND U32693 ( .A(a[11]), .B(b[75]), .Z(n25967) );
  XOR U32694 ( .A(n25973), .B(n25974), .Z(n25461) );
  ANDN U32695 ( .B(n25975), .A(n25976), .Z(n25973) );
  AND U32696 ( .A(a[12]), .B(b[74]), .Z(n25972) );
  IV U32697 ( .A(n25468), .Z(n25902) );
  XOR U32698 ( .A(n25978), .B(n25979), .Z(n25466) );
  ANDN U32699 ( .B(n25980), .A(n25981), .Z(n25978) );
  AND U32700 ( .A(a[13]), .B(b[73]), .Z(n25977) );
  XOR U32701 ( .A(n25983), .B(n25984), .Z(n25471) );
  ANDN U32702 ( .B(n25985), .A(n25986), .Z(n25983) );
  AND U32703 ( .A(a[14]), .B(b[72]), .Z(n25982) );
  XOR U32704 ( .A(n25988), .B(n25989), .Z(n25476) );
  ANDN U32705 ( .B(n25990), .A(n25991), .Z(n25988) );
  AND U32706 ( .A(a[15]), .B(b[71]), .Z(n25987) );
  XOR U32707 ( .A(n25993), .B(n25994), .Z(n25481) );
  ANDN U32708 ( .B(n25995), .A(n25996), .Z(n25993) );
  AND U32709 ( .A(a[16]), .B(b[70]), .Z(n25992) );
  XOR U32710 ( .A(n25998), .B(n25999), .Z(n25486) );
  ANDN U32711 ( .B(n26000), .A(n26001), .Z(n25998) );
  AND U32712 ( .A(a[17]), .B(b[69]), .Z(n25997) );
  XOR U32713 ( .A(n26003), .B(n26004), .Z(n25491) );
  ANDN U32714 ( .B(n26005), .A(n26006), .Z(n26003) );
  AND U32715 ( .A(a[18]), .B(b[68]), .Z(n26002) );
  XOR U32716 ( .A(n26008), .B(n26009), .Z(n25496) );
  ANDN U32717 ( .B(n26010), .A(n26011), .Z(n26008) );
  AND U32718 ( .A(a[19]), .B(b[67]), .Z(n26007) );
  XOR U32719 ( .A(n26013), .B(n26014), .Z(n25501) );
  ANDN U32720 ( .B(n26015), .A(n26016), .Z(n26013) );
  AND U32721 ( .A(a[20]), .B(b[66]), .Z(n26012) );
  XOR U32722 ( .A(n26018), .B(n26019), .Z(n25506) );
  ANDN U32723 ( .B(n26020), .A(n26021), .Z(n26018) );
  AND U32724 ( .A(a[21]), .B(b[65]), .Z(n26017) );
  XOR U32725 ( .A(n26023), .B(n26024), .Z(n25511) );
  ANDN U32726 ( .B(n26025), .A(n26026), .Z(n26023) );
  AND U32727 ( .A(a[22]), .B(b[64]), .Z(n26022) );
  XOR U32728 ( .A(n26028), .B(n26029), .Z(n25516) );
  ANDN U32729 ( .B(n26030), .A(n26031), .Z(n26028) );
  AND U32730 ( .A(a[23]), .B(b[63]), .Z(n26027) );
  XOR U32731 ( .A(n26033), .B(n26034), .Z(n25521) );
  ANDN U32732 ( .B(n26035), .A(n26036), .Z(n26033) );
  AND U32733 ( .A(a[24]), .B(b[62]), .Z(n26032) );
  XOR U32734 ( .A(n26038), .B(n26039), .Z(n25526) );
  ANDN U32735 ( .B(n26040), .A(n26041), .Z(n26038) );
  AND U32736 ( .A(a[25]), .B(b[61]), .Z(n26037) );
  XOR U32737 ( .A(n26043), .B(n26044), .Z(n25531) );
  ANDN U32738 ( .B(n26045), .A(n26046), .Z(n26043) );
  AND U32739 ( .A(a[26]), .B(b[60]), .Z(n26042) );
  XOR U32740 ( .A(n26048), .B(n26049), .Z(n25536) );
  ANDN U32741 ( .B(n26050), .A(n26051), .Z(n26048) );
  AND U32742 ( .A(a[27]), .B(b[59]), .Z(n26047) );
  XOR U32743 ( .A(n26053), .B(n26054), .Z(n25541) );
  ANDN U32744 ( .B(n26055), .A(n26056), .Z(n26053) );
  AND U32745 ( .A(a[28]), .B(b[58]), .Z(n26052) );
  XOR U32746 ( .A(n26058), .B(n26059), .Z(n25546) );
  ANDN U32747 ( .B(n26060), .A(n26061), .Z(n26058) );
  AND U32748 ( .A(a[29]), .B(b[57]), .Z(n26057) );
  XOR U32749 ( .A(n26063), .B(n26064), .Z(n25551) );
  ANDN U32750 ( .B(n26065), .A(n26066), .Z(n26063) );
  AND U32751 ( .A(a[30]), .B(b[56]), .Z(n26062) );
  XOR U32752 ( .A(n26068), .B(n26069), .Z(n25556) );
  ANDN U32753 ( .B(n26070), .A(n26071), .Z(n26068) );
  AND U32754 ( .A(a[31]), .B(b[55]), .Z(n26067) );
  XOR U32755 ( .A(n26073), .B(n26074), .Z(n25561) );
  ANDN U32756 ( .B(n26075), .A(n26076), .Z(n26073) );
  AND U32757 ( .A(a[32]), .B(b[54]), .Z(n26072) );
  XOR U32758 ( .A(n26078), .B(n26079), .Z(n25566) );
  ANDN U32759 ( .B(n26080), .A(n26081), .Z(n26078) );
  AND U32760 ( .A(a[33]), .B(b[53]), .Z(n26077) );
  XOR U32761 ( .A(n26083), .B(n26084), .Z(n25571) );
  ANDN U32762 ( .B(n26085), .A(n26086), .Z(n26083) );
  AND U32763 ( .A(a[34]), .B(b[52]), .Z(n26082) );
  XOR U32764 ( .A(n26088), .B(n26089), .Z(n25576) );
  ANDN U32765 ( .B(n26090), .A(n26091), .Z(n26088) );
  AND U32766 ( .A(a[35]), .B(b[51]), .Z(n26087) );
  XOR U32767 ( .A(n26093), .B(n26094), .Z(n25581) );
  ANDN U32768 ( .B(n26095), .A(n26096), .Z(n26093) );
  AND U32769 ( .A(a[36]), .B(b[50]), .Z(n26092) );
  XOR U32770 ( .A(n26098), .B(n26099), .Z(n25586) );
  ANDN U32771 ( .B(n26100), .A(n26101), .Z(n26098) );
  AND U32772 ( .A(a[37]), .B(b[49]), .Z(n26097) );
  XOR U32773 ( .A(n26103), .B(n26104), .Z(n25591) );
  ANDN U32774 ( .B(n26105), .A(n26106), .Z(n26103) );
  AND U32775 ( .A(a[38]), .B(b[48]), .Z(n26102) );
  XOR U32776 ( .A(n26108), .B(n26109), .Z(n25596) );
  ANDN U32777 ( .B(n26110), .A(n26111), .Z(n26108) );
  AND U32778 ( .A(a[39]), .B(b[47]), .Z(n26107) );
  XOR U32779 ( .A(n26113), .B(n26114), .Z(n25601) );
  ANDN U32780 ( .B(n26115), .A(n26116), .Z(n26113) );
  AND U32781 ( .A(a[40]), .B(b[46]), .Z(n26112) );
  XOR U32782 ( .A(n26118), .B(n26119), .Z(n25606) );
  ANDN U32783 ( .B(n26120), .A(n26121), .Z(n26118) );
  AND U32784 ( .A(a[41]), .B(b[45]), .Z(n26117) );
  XOR U32785 ( .A(n26123), .B(n26124), .Z(n25611) );
  ANDN U32786 ( .B(n26125), .A(n26126), .Z(n26123) );
  AND U32787 ( .A(a[42]), .B(b[44]), .Z(n26122) );
  XOR U32788 ( .A(n26128), .B(n26129), .Z(n25616) );
  ANDN U32789 ( .B(n26130), .A(n26131), .Z(n26128) );
  AND U32790 ( .A(a[43]), .B(b[43]), .Z(n26127) );
  XOR U32791 ( .A(n26133), .B(n26134), .Z(n25621) );
  ANDN U32792 ( .B(n26135), .A(n26136), .Z(n26133) );
  AND U32793 ( .A(a[44]), .B(b[42]), .Z(n26132) );
  XOR U32794 ( .A(n26138), .B(n26139), .Z(n25626) );
  ANDN U32795 ( .B(n26140), .A(n26141), .Z(n26138) );
  AND U32796 ( .A(a[45]), .B(b[41]), .Z(n26137) );
  XOR U32797 ( .A(n26143), .B(n26144), .Z(n25631) );
  ANDN U32798 ( .B(n26145), .A(n26146), .Z(n26143) );
  AND U32799 ( .A(a[46]), .B(b[40]), .Z(n26142) );
  XOR U32800 ( .A(n26148), .B(n26149), .Z(n25636) );
  ANDN U32801 ( .B(n26150), .A(n26151), .Z(n26148) );
  AND U32802 ( .A(a[47]), .B(b[39]), .Z(n26147) );
  XOR U32803 ( .A(n26153), .B(n26154), .Z(n25641) );
  ANDN U32804 ( .B(n26155), .A(n26156), .Z(n26153) );
  AND U32805 ( .A(a[48]), .B(b[38]), .Z(n26152) );
  XOR U32806 ( .A(n26158), .B(n26159), .Z(n25646) );
  ANDN U32807 ( .B(n26160), .A(n26161), .Z(n26158) );
  AND U32808 ( .A(a[49]), .B(b[37]), .Z(n26157) );
  XOR U32809 ( .A(n26163), .B(n26164), .Z(n25651) );
  ANDN U32810 ( .B(n26165), .A(n26166), .Z(n26163) );
  AND U32811 ( .A(a[50]), .B(b[36]), .Z(n26162) );
  XOR U32812 ( .A(n26168), .B(n26169), .Z(n25656) );
  ANDN U32813 ( .B(n26170), .A(n26171), .Z(n26168) );
  AND U32814 ( .A(a[51]), .B(b[35]), .Z(n26167) );
  XOR U32815 ( .A(n26173), .B(n26174), .Z(n25661) );
  ANDN U32816 ( .B(n26175), .A(n26176), .Z(n26173) );
  AND U32817 ( .A(a[52]), .B(b[34]), .Z(n26172) );
  XOR U32818 ( .A(n26178), .B(n26179), .Z(n25666) );
  ANDN U32819 ( .B(n26180), .A(n26181), .Z(n26178) );
  AND U32820 ( .A(a[53]), .B(b[33]), .Z(n26177) );
  XOR U32821 ( .A(n26183), .B(n26184), .Z(n25671) );
  ANDN U32822 ( .B(n26185), .A(n26186), .Z(n26183) );
  AND U32823 ( .A(a[54]), .B(b[32]), .Z(n26182) );
  XOR U32824 ( .A(n26188), .B(n26189), .Z(n25676) );
  ANDN U32825 ( .B(n26190), .A(n26191), .Z(n26188) );
  AND U32826 ( .A(a[55]), .B(b[31]), .Z(n26187) );
  XOR U32827 ( .A(n26193), .B(n26194), .Z(n25681) );
  ANDN U32828 ( .B(n26195), .A(n26196), .Z(n26193) );
  AND U32829 ( .A(a[56]), .B(b[30]), .Z(n26192) );
  XOR U32830 ( .A(n26198), .B(n26199), .Z(n25686) );
  ANDN U32831 ( .B(n26200), .A(n26201), .Z(n26198) );
  AND U32832 ( .A(a[57]), .B(b[29]), .Z(n26197) );
  XOR U32833 ( .A(n26203), .B(n26204), .Z(n25691) );
  ANDN U32834 ( .B(n26205), .A(n26206), .Z(n26203) );
  AND U32835 ( .A(a[58]), .B(b[28]), .Z(n26202) );
  XOR U32836 ( .A(n26208), .B(n26209), .Z(n25696) );
  ANDN U32837 ( .B(n26210), .A(n26211), .Z(n26208) );
  AND U32838 ( .A(a[59]), .B(b[27]), .Z(n26207) );
  XOR U32839 ( .A(n26213), .B(n26214), .Z(n25701) );
  ANDN U32840 ( .B(n26215), .A(n26216), .Z(n26213) );
  AND U32841 ( .A(a[60]), .B(b[26]), .Z(n26212) );
  XOR U32842 ( .A(n26218), .B(n26219), .Z(n25706) );
  ANDN U32843 ( .B(n26220), .A(n26221), .Z(n26218) );
  AND U32844 ( .A(a[61]), .B(b[25]), .Z(n26217) );
  XOR U32845 ( .A(n26223), .B(n26224), .Z(n25711) );
  ANDN U32846 ( .B(n26225), .A(n26226), .Z(n26223) );
  AND U32847 ( .A(a[62]), .B(b[24]), .Z(n26222) );
  XOR U32848 ( .A(n26228), .B(n26229), .Z(n25716) );
  ANDN U32849 ( .B(n26230), .A(n26231), .Z(n26228) );
  AND U32850 ( .A(a[63]), .B(b[23]), .Z(n26227) );
  XOR U32851 ( .A(n26233), .B(n26234), .Z(n25721) );
  ANDN U32852 ( .B(n26235), .A(n26236), .Z(n26233) );
  AND U32853 ( .A(a[64]), .B(b[22]), .Z(n26232) );
  XOR U32854 ( .A(n26238), .B(n26239), .Z(n25726) );
  ANDN U32855 ( .B(n26240), .A(n26241), .Z(n26238) );
  AND U32856 ( .A(a[65]), .B(b[21]), .Z(n26237) );
  XOR U32857 ( .A(n26243), .B(n26244), .Z(n25731) );
  ANDN U32858 ( .B(n26245), .A(n26246), .Z(n26243) );
  AND U32859 ( .A(a[66]), .B(b[20]), .Z(n26242) );
  XOR U32860 ( .A(n26248), .B(n26249), .Z(n25736) );
  ANDN U32861 ( .B(n26250), .A(n26251), .Z(n26248) );
  AND U32862 ( .A(a[67]), .B(b[19]), .Z(n26247) );
  XOR U32863 ( .A(n26253), .B(n26254), .Z(n25741) );
  ANDN U32864 ( .B(n26255), .A(n26256), .Z(n26253) );
  AND U32865 ( .A(a[68]), .B(b[18]), .Z(n26252) );
  XOR U32866 ( .A(n26258), .B(n26259), .Z(n25746) );
  ANDN U32867 ( .B(n26260), .A(n26261), .Z(n26258) );
  AND U32868 ( .A(a[69]), .B(b[17]), .Z(n26257) );
  XOR U32869 ( .A(n26263), .B(n26264), .Z(n25751) );
  ANDN U32870 ( .B(n26265), .A(n26266), .Z(n26263) );
  AND U32871 ( .A(a[70]), .B(b[16]), .Z(n26262) );
  XOR U32872 ( .A(n26268), .B(n26269), .Z(n25756) );
  ANDN U32873 ( .B(n26270), .A(n26271), .Z(n26268) );
  AND U32874 ( .A(a[71]), .B(b[15]), .Z(n26267) );
  XOR U32875 ( .A(n26273), .B(n26274), .Z(n25761) );
  ANDN U32876 ( .B(n26275), .A(n26276), .Z(n26273) );
  AND U32877 ( .A(a[72]), .B(b[14]), .Z(n26272) );
  XOR U32878 ( .A(n26278), .B(n26279), .Z(n25766) );
  ANDN U32879 ( .B(n26280), .A(n26281), .Z(n26278) );
  AND U32880 ( .A(a[73]), .B(b[13]), .Z(n26277) );
  XOR U32881 ( .A(n26283), .B(n26284), .Z(n25771) );
  ANDN U32882 ( .B(n26285), .A(n26286), .Z(n26283) );
  AND U32883 ( .A(a[74]), .B(b[12]), .Z(n26282) );
  XOR U32884 ( .A(n26288), .B(n26289), .Z(n25776) );
  ANDN U32885 ( .B(n26290), .A(n26291), .Z(n26288) );
  AND U32886 ( .A(a[75]), .B(b[11]), .Z(n26287) );
  XOR U32887 ( .A(n26293), .B(n26294), .Z(n25781) );
  ANDN U32888 ( .B(n26295), .A(n26296), .Z(n26293) );
  AND U32889 ( .A(a[76]), .B(b[10]), .Z(n26292) );
  XOR U32890 ( .A(n26298), .B(n26299), .Z(n25786) );
  ANDN U32891 ( .B(n26300), .A(n26301), .Z(n26298) );
  AND U32892 ( .A(b[9]), .B(a[77]), .Z(n26297) );
  XOR U32893 ( .A(n26303), .B(n26304), .Z(n25791) );
  ANDN U32894 ( .B(n26305), .A(n26306), .Z(n26303) );
  AND U32895 ( .A(b[8]), .B(a[78]), .Z(n26302) );
  XOR U32896 ( .A(n26308), .B(n26309), .Z(n25796) );
  ANDN U32897 ( .B(n26310), .A(n26311), .Z(n26308) );
  AND U32898 ( .A(b[7]), .B(a[79]), .Z(n26307) );
  XOR U32899 ( .A(n26313), .B(n26314), .Z(n25801) );
  ANDN U32900 ( .B(n26315), .A(n26316), .Z(n26313) );
  AND U32901 ( .A(b[6]), .B(a[80]), .Z(n26312) );
  XOR U32902 ( .A(n26318), .B(n26319), .Z(n25806) );
  ANDN U32903 ( .B(n26320), .A(n26321), .Z(n26318) );
  AND U32904 ( .A(b[5]), .B(a[81]), .Z(n26317) );
  XOR U32905 ( .A(n26323), .B(n26324), .Z(n25811) );
  ANDN U32906 ( .B(n26325), .A(n26326), .Z(n26323) );
  AND U32907 ( .A(b[4]), .B(a[82]), .Z(n26322) );
  XOR U32908 ( .A(n26328), .B(n26329), .Z(n25816) );
  ANDN U32909 ( .B(n25828), .A(n25829), .Z(n26328) );
  AND U32910 ( .A(b[2]), .B(a[83]), .Z(n26330) );
  XNOR U32911 ( .A(n26325), .B(n26329), .Z(n26331) );
  XOR U32912 ( .A(n26332), .B(n26333), .Z(n26329) );
  OR U32913 ( .A(n25831), .B(n25832), .Z(n26333) );
  XNOR U32914 ( .A(n26335), .B(n26336), .Z(n26334) );
  XOR U32915 ( .A(n26335), .B(n26338), .Z(n25831) );
  NAND U32916 ( .A(b[1]), .B(a[83]), .Z(n26338) );
  IV U32917 ( .A(n26332), .Z(n26335) );
  NANDN U32918 ( .A(n37), .B(n38), .Z(n26332) );
  XOR U32919 ( .A(n26339), .B(n26340), .Z(n38) );
  NAND U32920 ( .A(a[83]), .B(b[0]), .Z(n37) );
  XNOR U32921 ( .A(n26320), .B(n26324), .Z(n26341) );
  XNOR U32922 ( .A(n26315), .B(n26319), .Z(n26342) );
  XNOR U32923 ( .A(n26310), .B(n26314), .Z(n26343) );
  XNOR U32924 ( .A(n26305), .B(n26309), .Z(n26344) );
  XNOR U32925 ( .A(n26300), .B(n26304), .Z(n26345) );
  XNOR U32926 ( .A(n26295), .B(n26299), .Z(n26346) );
  XNOR U32927 ( .A(n26290), .B(n26294), .Z(n26347) );
  XNOR U32928 ( .A(n26285), .B(n26289), .Z(n26348) );
  XNOR U32929 ( .A(n26280), .B(n26284), .Z(n26349) );
  XNOR U32930 ( .A(n26275), .B(n26279), .Z(n26350) );
  XNOR U32931 ( .A(n26270), .B(n26274), .Z(n26351) );
  XNOR U32932 ( .A(n26265), .B(n26269), .Z(n26352) );
  XNOR U32933 ( .A(n26260), .B(n26264), .Z(n26353) );
  XNOR U32934 ( .A(n26255), .B(n26259), .Z(n26354) );
  XNOR U32935 ( .A(n26250), .B(n26254), .Z(n26355) );
  XNOR U32936 ( .A(n26245), .B(n26249), .Z(n26356) );
  XNOR U32937 ( .A(n26240), .B(n26244), .Z(n26357) );
  XNOR U32938 ( .A(n26235), .B(n26239), .Z(n26358) );
  XNOR U32939 ( .A(n26230), .B(n26234), .Z(n26359) );
  XNOR U32940 ( .A(n26225), .B(n26229), .Z(n26360) );
  XNOR U32941 ( .A(n26220), .B(n26224), .Z(n26361) );
  XNOR U32942 ( .A(n26215), .B(n26219), .Z(n26362) );
  XNOR U32943 ( .A(n26210), .B(n26214), .Z(n26363) );
  XNOR U32944 ( .A(n26205), .B(n26209), .Z(n26364) );
  XNOR U32945 ( .A(n26200), .B(n26204), .Z(n26365) );
  XNOR U32946 ( .A(n26195), .B(n26199), .Z(n26366) );
  XNOR U32947 ( .A(n26190), .B(n26194), .Z(n26367) );
  XNOR U32948 ( .A(n26185), .B(n26189), .Z(n26368) );
  XNOR U32949 ( .A(n26180), .B(n26184), .Z(n26369) );
  XNOR U32950 ( .A(n26175), .B(n26179), .Z(n26370) );
  XNOR U32951 ( .A(n26170), .B(n26174), .Z(n26371) );
  XNOR U32952 ( .A(n26165), .B(n26169), .Z(n26372) );
  XNOR U32953 ( .A(n26160), .B(n26164), .Z(n26373) );
  XNOR U32954 ( .A(n26155), .B(n26159), .Z(n26374) );
  XNOR U32955 ( .A(n26150), .B(n26154), .Z(n26375) );
  XNOR U32956 ( .A(n26145), .B(n26149), .Z(n26376) );
  XNOR U32957 ( .A(n26140), .B(n26144), .Z(n26377) );
  XNOR U32958 ( .A(n26135), .B(n26139), .Z(n26378) );
  XNOR U32959 ( .A(n26130), .B(n26134), .Z(n26379) );
  XNOR U32960 ( .A(n26125), .B(n26129), .Z(n26380) );
  XNOR U32961 ( .A(n26120), .B(n26124), .Z(n26381) );
  XNOR U32962 ( .A(n26115), .B(n26119), .Z(n26382) );
  XNOR U32963 ( .A(n26110), .B(n26114), .Z(n26383) );
  XNOR U32964 ( .A(n26105), .B(n26109), .Z(n26384) );
  XNOR U32965 ( .A(n26100), .B(n26104), .Z(n26385) );
  XNOR U32966 ( .A(n26095), .B(n26099), .Z(n26386) );
  XNOR U32967 ( .A(n26090), .B(n26094), .Z(n26387) );
  XNOR U32968 ( .A(n26085), .B(n26089), .Z(n26388) );
  XNOR U32969 ( .A(n26080), .B(n26084), .Z(n26389) );
  XNOR U32970 ( .A(n26075), .B(n26079), .Z(n26390) );
  XNOR U32971 ( .A(n26070), .B(n26074), .Z(n26391) );
  XNOR U32972 ( .A(n26065), .B(n26069), .Z(n26392) );
  XNOR U32973 ( .A(n26060), .B(n26064), .Z(n26393) );
  XNOR U32974 ( .A(n26055), .B(n26059), .Z(n26394) );
  XNOR U32975 ( .A(n26050), .B(n26054), .Z(n26395) );
  XNOR U32976 ( .A(n26045), .B(n26049), .Z(n26396) );
  XNOR U32977 ( .A(n26040), .B(n26044), .Z(n26397) );
  XNOR U32978 ( .A(n26035), .B(n26039), .Z(n26398) );
  XNOR U32979 ( .A(n26030), .B(n26034), .Z(n26399) );
  XNOR U32980 ( .A(n26025), .B(n26029), .Z(n26400) );
  XNOR U32981 ( .A(n26020), .B(n26024), .Z(n26401) );
  XNOR U32982 ( .A(n26015), .B(n26019), .Z(n26402) );
  XNOR U32983 ( .A(n26010), .B(n26014), .Z(n26403) );
  XNOR U32984 ( .A(n26005), .B(n26009), .Z(n26404) );
  XNOR U32985 ( .A(n26000), .B(n26004), .Z(n26405) );
  XNOR U32986 ( .A(n25995), .B(n25999), .Z(n26406) );
  XNOR U32987 ( .A(n25990), .B(n25994), .Z(n26407) );
  XNOR U32988 ( .A(n25985), .B(n25989), .Z(n26408) );
  XNOR U32989 ( .A(n25980), .B(n25984), .Z(n26409) );
  XNOR U32990 ( .A(n25975), .B(n25979), .Z(n26410) );
  XNOR U32991 ( .A(n25970), .B(n25974), .Z(n26411) );
  XNOR U32992 ( .A(n25965), .B(n25969), .Z(n26412) );
  XNOR U32993 ( .A(n25960), .B(n25964), .Z(n26413) );
  XNOR U32994 ( .A(n25955), .B(n25959), .Z(n26414) );
  XNOR U32995 ( .A(n25950), .B(n25954), .Z(n26415) );
  XNOR U32996 ( .A(n25945), .B(n25949), .Z(n26416) );
  XNOR U32997 ( .A(n25940), .B(n25944), .Z(n26417) );
  XNOR U32998 ( .A(n25935), .B(n25939), .Z(n26418) );
  XNOR U32999 ( .A(n25930), .B(n25934), .Z(n26419) );
  XNOR U33000 ( .A(n25925), .B(n25929), .Z(n26420) );
  XNOR U33001 ( .A(n25920), .B(n25924), .Z(n26421) );
  XNOR U33002 ( .A(n26422), .B(n25919), .Z(n25920) );
  AND U33003 ( .A(a[0]), .B(b[85]), .Z(n26422) );
  XOR U33004 ( .A(n26423), .B(n25919), .Z(n25921) );
  XNOR U33005 ( .A(n26424), .B(n26425), .Z(n25919) );
  ANDN U33006 ( .B(n26426), .A(n26427), .Z(n26424) );
  AND U33007 ( .A(a[1]), .B(b[84]), .Z(n26423) );
  XOR U33008 ( .A(n26429), .B(n26430), .Z(n25924) );
  ANDN U33009 ( .B(n26431), .A(n26432), .Z(n26429) );
  AND U33010 ( .A(a[2]), .B(b[83]), .Z(n26428) );
  XOR U33011 ( .A(n26434), .B(n26435), .Z(n25929) );
  ANDN U33012 ( .B(n26436), .A(n26437), .Z(n26434) );
  AND U33013 ( .A(a[3]), .B(b[82]), .Z(n26433) );
  XOR U33014 ( .A(n26439), .B(n26440), .Z(n25934) );
  ANDN U33015 ( .B(n26441), .A(n26442), .Z(n26439) );
  AND U33016 ( .A(a[4]), .B(b[81]), .Z(n26438) );
  XOR U33017 ( .A(n26444), .B(n26445), .Z(n25939) );
  ANDN U33018 ( .B(n26446), .A(n26447), .Z(n26444) );
  AND U33019 ( .A(a[5]), .B(b[80]), .Z(n26443) );
  XOR U33020 ( .A(n26449), .B(n26450), .Z(n25944) );
  ANDN U33021 ( .B(n26451), .A(n26452), .Z(n26449) );
  AND U33022 ( .A(a[6]), .B(b[79]), .Z(n26448) );
  XOR U33023 ( .A(n26454), .B(n26455), .Z(n25949) );
  ANDN U33024 ( .B(n26456), .A(n26457), .Z(n26454) );
  AND U33025 ( .A(a[7]), .B(b[78]), .Z(n26453) );
  XOR U33026 ( .A(n26459), .B(n26460), .Z(n25954) );
  ANDN U33027 ( .B(n26461), .A(n26462), .Z(n26459) );
  AND U33028 ( .A(a[8]), .B(b[77]), .Z(n26458) );
  XOR U33029 ( .A(n26464), .B(n26465), .Z(n25959) );
  ANDN U33030 ( .B(n26466), .A(n26467), .Z(n26464) );
  AND U33031 ( .A(a[9]), .B(b[76]), .Z(n26463) );
  XOR U33032 ( .A(n26469), .B(n26470), .Z(n25964) );
  ANDN U33033 ( .B(n26471), .A(n26472), .Z(n26469) );
  AND U33034 ( .A(a[10]), .B(b[75]), .Z(n26468) );
  XOR U33035 ( .A(n26474), .B(n26475), .Z(n25969) );
  ANDN U33036 ( .B(n26476), .A(n26477), .Z(n26474) );
  AND U33037 ( .A(a[11]), .B(b[74]), .Z(n26473) );
  XOR U33038 ( .A(n26479), .B(n26480), .Z(n25974) );
  ANDN U33039 ( .B(n26481), .A(n26482), .Z(n26479) );
  AND U33040 ( .A(a[12]), .B(b[73]), .Z(n26478) );
  XOR U33041 ( .A(n26484), .B(n26485), .Z(n25979) );
  ANDN U33042 ( .B(n26486), .A(n26487), .Z(n26484) );
  AND U33043 ( .A(a[13]), .B(b[72]), .Z(n26483) );
  XOR U33044 ( .A(n26489), .B(n26490), .Z(n25984) );
  ANDN U33045 ( .B(n26491), .A(n26492), .Z(n26489) );
  AND U33046 ( .A(a[14]), .B(b[71]), .Z(n26488) );
  XOR U33047 ( .A(n26494), .B(n26495), .Z(n25989) );
  ANDN U33048 ( .B(n26496), .A(n26497), .Z(n26494) );
  AND U33049 ( .A(a[15]), .B(b[70]), .Z(n26493) );
  XOR U33050 ( .A(n26499), .B(n26500), .Z(n25994) );
  ANDN U33051 ( .B(n26501), .A(n26502), .Z(n26499) );
  AND U33052 ( .A(a[16]), .B(b[69]), .Z(n26498) );
  XOR U33053 ( .A(n26504), .B(n26505), .Z(n25999) );
  ANDN U33054 ( .B(n26506), .A(n26507), .Z(n26504) );
  AND U33055 ( .A(a[17]), .B(b[68]), .Z(n26503) );
  XOR U33056 ( .A(n26509), .B(n26510), .Z(n26004) );
  ANDN U33057 ( .B(n26511), .A(n26512), .Z(n26509) );
  AND U33058 ( .A(a[18]), .B(b[67]), .Z(n26508) );
  XOR U33059 ( .A(n26514), .B(n26515), .Z(n26009) );
  ANDN U33060 ( .B(n26516), .A(n26517), .Z(n26514) );
  AND U33061 ( .A(a[19]), .B(b[66]), .Z(n26513) );
  XOR U33062 ( .A(n26519), .B(n26520), .Z(n26014) );
  ANDN U33063 ( .B(n26521), .A(n26522), .Z(n26519) );
  AND U33064 ( .A(a[20]), .B(b[65]), .Z(n26518) );
  XOR U33065 ( .A(n26524), .B(n26525), .Z(n26019) );
  ANDN U33066 ( .B(n26526), .A(n26527), .Z(n26524) );
  AND U33067 ( .A(a[21]), .B(b[64]), .Z(n26523) );
  XOR U33068 ( .A(n26529), .B(n26530), .Z(n26024) );
  ANDN U33069 ( .B(n26531), .A(n26532), .Z(n26529) );
  AND U33070 ( .A(a[22]), .B(b[63]), .Z(n26528) );
  XOR U33071 ( .A(n26534), .B(n26535), .Z(n26029) );
  ANDN U33072 ( .B(n26536), .A(n26537), .Z(n26534) );
  AND U33073 ( .A(a[23]), .B(b[62]), .Z(n26533) );
  XOR U33074 ( .A(n26539), .B(n26540), .Z(n26034) );
  ANDN U33075 ( .B(n26541), .A(n26542), .Z(n26539) );
  AND U33076 ( .A(a[24]), .B(b[61]), .Z(n26538) );
  XOR U33077 ( .A(n26544), .B(n26545), .Z(n26039) );
  ANDN U33078 ( .B(n26546), .A(n26547), .Z(n26544) );
  AND U33079 ( .A(a[25]), .B(b[60]), .Z(n26543) );
  XOR U33080 ( .A(n26549), .B(n26550), .Z(n26044) );
  ANDN U33081 ( .B(n26551), .A(n26552), .Z(n26549) );
  AND U33082 ( .A(a[26]), .B(b[59]), .Z(n26548) );
  XOR U33083 ( .A(n26554), .B(n26555), .Z(n26049) );
  ANDN U33084 ( .B(n26556), .A(n26557), .Z(n26554) );
  AND U33085 ( .A(a[27]), .B(b[58]), .Z(n26553) );
  XOR U33086 ( .A(n26559), .B(n26560), .Z(n26054) );
  ANDN U33087 ( .B(n26561), .A(n26562), .Z(n26559) );
  AND U33088 ( .A(a[28]), .B(b[57]), .Z(n26558) );
  XOR U33089 ( .A(n26564), .B(n26565), .Z(n26059) );
  ANDN U33090 ( .B(n26566), .A(n26567), .Z(n26564) );
  AND U33091 ( .A(a[29]), .B(b[56]), .Z(n26563) );
  XOR U33092 ( .A(n26569), .B(n26570), .Z(n26064) );
  ANDN U33093 ( .B(n26571), .A(n26572), .Z(n26569) );
  AND U33094 ( .A(a[30]), .B(b[55]), .Z(n26568) );
  XOR U33095 ( .A(n26574), .B(n26575), .Z(n26069) );
  ANDN U33096 ( .B(n26576), .A(n26577), .Z(n26574) );
  AND U33097 ( .A(a[31]), .B(b[54]), .Z(n26573) );
  XOR U33098 ( .A(n26579), .B(n26580), .Z(n26074) );
  ANDN U33099 ( .B(n26581), .A(n26582), .Z(n26579) );
  AND U33100 ( .A(a[32]), .B(b[53]), .Z(n26578) );
  XOR U33101 ( .A(n26584), .B(n26585), .Z(n26079) );
  ANDN U33102 ( .B(n26586), .A(n26587), .Z(n26584) );
  AND U33103 ( .A(a[33]), .B(b[52]), .Z(n26583) );
  XOR U33104 ( .A(n26589), .B(n26590), .Z(n26084) );
  ANDN U33105 ( .B(n26591), .A(n26592), .Z(n26589) );
  AND U33106 ( .A(a[34]), .B(b[51]), .Z(n26588) );
  XOR U33107 ( .A(n26594), .B(n26595), .Z(n26089) );
  ANDN U33108 ( .B(n26596), .A(n26597), .Z(n26594) );
  AND U33109 ( .A(a[35]), .B(b[50]), .Z(n26593) );
  XOR U33110 ( .A(n26599), .B(n26600), .Z(n26094) );
  ANDN U33111 ( .B(n26601), .A(n26602), .Z(n26599) );
  AND U33112 ( .A(a[36]), .B(b[49]), .Z(n26598) );
  XOR U33113 ( .A(n26604), .B(n26605), .Z(n26099) );
  ANDN U33114 ( .B(n26606), .A(n26607), .Z(n26604) );
  AND U33115 ( .A(a[37]), .B(b[48]), .Z(n26603) );
  XOR U33116 ( .A(n26609), .B(n26610), .Z(n26104) );
  ANDN U33117 ( .B(n26611), .A(n26612), .Z(n26609) );
  AND U33118 ( .A(a[38]), .B(b[47]), .Z(n26608) );
  XOR U33119 ( .A(n26614), .B(n26615), .Z(n26109) );
  ANDN U33120 ( .B(n26616), .A(n26617), .Z(n26614) );
  AND U33121 ( .A(a[39]), .B(b[46]), .Z(n26613) );
  XOR U33122 ( .A(n26619), .B(n26620), .Z(n26114) );
  ANDN U33123 ( .B(n26621), .A(n26622), .Z(n26619) );
  AND U33124 ( .A(a[40]), .B(b[45]), .Z(n26618) );
  XOR U33125 ( .A(n26624), .B(n26625), .Z(n26119) );
  ANDN U33126 ( .B(n26626), .A(n26627), .Z(n26624) );
  AND U33127 ( .A(a[41]), .B(b[44]), .Z(n26623) );
  XOR U33128 ( .A(n26629), .B(n26630), .Z(n26124) );
  ANDN U33129 ( .B(n26631), .A(n26632), .Z(n26629) );
  AND U33130 ( .A(a[42]), .B(b[43]), .Z(n26628) );
  XOR U33131 ( .A(n26634), .B(n26635), .Z(n26129) );
  ANDN U33132 ( .B(n26636), .A(n26637), .Z(n26634) );
  AND U33133 ( .A(a[43]), .B(b[42]), .Z(n26633) );
  XOR U33134 ( .A(n26639), .B(n26640), .Z(n26134) );
  ANDN U33135 ( .B(n26641), .A(n26642), .Z(n26639) );
  AND U33136 ( .A(a[44]), .B(b[41]), .Z(n26638) );
  XOR U33137 ( .A(n26644), .B(n26645), .Z(n26139) );
  ANDN U33138 ( .B(n26646), .A(n26647), .Z(n26644) );
  AND U33139 ( .A(a[45]), .B(b[40]), .Z(n26643) );
  XOR U33140 ( .A(n26649), .B(n26650), .Z(n26144) );
  ANDN U33141 ( .B(n26651), .A(n26652), .Z(n26649) );
  AND U33142 ( .A(a[46]), .B(b[39]), .Z(n26648) );
  XOR U33143 ( .A(n26654), .B(n26655), .Z(n26149) );
  ANDN U33144 ( .B(n26656), .A(n26657), .Z(n26654) );
  AND U33145 ( .A(a[47]), .B(b[38]), .Z(n26653) );
  XOR U33146 ( .A(n26659), .B(n26660), .Z(n26154) );
  ANDN U33147 ( .B(n26661), .A(n26662), .Z(n26659) );
  AND U33148 ( .A(a[48]), .B(b[37]), .Z(n26658) );
  XOR U33149 ( .A(n26664), .B(n26665), .Z(n26159) );
  ANDN U33150 ( .B(n26666), .A(n26667), .Z(n26664) );
  AND U33151 ( .A(a[49]), .B(b[36]), .Z(n26663) );
  XOR U33152 ( .A(n26669), .B(n26670), .Z(n26164) );
  ANDN U33153 ( .B(n26671), .A(n26672), .Z(n26669) );
  AND U33154 ( .A(a[50]), .B(b[35]), .Z(n26668) );
  XOR U33155 ( .A(n26674), .B(n26675), .Z(n26169) );
  ANDN U33156 ( .B(n26676), .A(n26677), .Z(n26674) );
  AND U33157 ( .A(a[51]), .B(b[34]), .Z(n26673) );
  XOR U33158 ( .A(n26679), .B(n26680), .Z(n26174) );
  ANDN U33159 ( .B(n26681), .A(n26682), .Z(n26679) );
  AND U33160 ( .A(a[52]), .B(b[33]), .Z(n26678) );
  XOR U33161 ( .A(n26684), .B(n26685), .Z(n26179) );
  ANDN U33162 ( .B(n26686), .A(n26687), .Z(n26684) );
  AND U33163 ( .A(a[53]), .B(b[32]), .Z(n26683) );
  XOR U33164 ( .A(n26689), .B(n26690), .Z(n26184) );
  ANDN U33165 ( .B(n26691), .A(n26692), .Z(n26689) );
  AND U33166 ( .A(a[54]), .B(b[31]), .Z(n26688) );
  XOR U33167 ( .A(n26694), .B(n26695), .Z(n26189) );
  ANDN U33168 ( .B(n26696), .A(n26697), .Z(n26694) );
  AND U33169 ( .A(a[55]), .B(b[30]), .Z(n26693) );
  XOR U33170 ( .A(n26699), .B(n26700), .Z(n26194) );
  ANDN U33171 ( .B(n26701), .A(n26702), .Z(n26699) );
  AND U33172 ( .A(a[56]), .B(b[29]), .Z(n26698) );
  XOR U33173 ( .A(n26704), .B(n26705), .Z(n26199) );
  ANDN U33174 ( .B(n26706), .A(n26707), .Z(n26704) );
  AND U33175 ( .A(a[57]), .B(b[28]), .Z(n26703) );
  XOR U33176 ( .A(n26709), .B(n26710), .Z(n26204) );
  ANDN U33177 ( .B(n26711), .A(n26712), .Z(n26709) );
  AND U33178 ( .A(a[58]), .B(b[27]), .Z(n26708) );
  XOR U33179 ( .A(n26714), .B(n26715), .Z(n26209) );
  ANDN U33180 ( .B(n26716), .A(n26717), .Z(n26714) );
  AND U33181 ( .A(a[59]), .B(b[26]), .Z(n26713) );
  XOR U33182 ( .A(n26719), .B(n26720), .Z(n26214) );
  ANDN U33183 ( .B(n26721), .A(n26722), .Z(n26719) );
  AND U33184 ( .A(a[60]), .B(b[25]), .Z(n26718) );
  XOR U33185 ( .A(n26724), .B(n26725), .Z(n26219) );
  ANDN U33186 ( .B(n26726), .A(n26727), .Z(n26724) );
  AND U33187 ( .A(a[61]), .B(b[24]), .Z(n26723) );
  XOR U33188 ( .A(n26729), .B(n26730), .Z(n26224) );
  ANDN U33189 ( .B(n26731), .A(n26732), .Z(n26729) );
  AND U33190 ( .A(a[62]), .B(b[23]), .Z(n26728) );
  XOR U33191 ( .A(n26734), .B(n26735), .Z(n26229) );
  ANDN U33192 ( .B(n26736), .A(n26737), .Z(n26734) );
  AND U33193 ( .A(a[63]), .B(b[22]), .Z(n26733) );
  XOR U33194 ( .A(n26739), .B(n26740), .Z(n26234) );
  ANDN U33195 ( .B(n26741), .A(n26742), .Z(n26739) );
  AND U33196 ( .A(a[64]), .B(b[21]), .Z(n26738) );
  XOR U33197 ( .A(n26744), .B(n26745), .Z(n26239) );
  ANDN U33198 ( .B(n26746), .A(n26747), .Z(n26744) );
  AND U33199 ( .A(a[65]), .B(b[20]), .Z(n26743) );
  XOR U33200 ( .A(n26749), .B(n26750), .Z(n26244) );
  ANDN U33201 ( .B(n26751), .A(n26752), .Z(n26749) );
  AND U33202 ( .A(a[66]), .B(b[19]), .Z(n26748) );
  XOR U33203 ( .A(n26754), .B(n26755), .Z(n26249) );
  ANDN U33204 ( .B(n26756), .A(n26757), .Z(n26754) );
  AND U33205 ( .A(a[67]), .B(b[18]), .Z(n26753) );
  XOR U33206 ( .A(n26759), .B(n26760), .Z(n26254) );
  ANDN U33207 ( .B(n26761), .A(n26762), .Z(n26759) );
  AND U33208 ( .A(a[68]), .B(b[17]), .Z(n26758) );
  XOR U33209 ( .A(n26764), .B(n26765), .Z(n26259) );
  ANDN U33210 ( .B(n26766), .A(n26767), .Z(n26764) );
  AND U33211 ( .A(a[69]), .B(b[16]), .Z(n26763) );
  XOR U33212 ( .A(n26769), .B(n26770), .Z(n26264) );
  ANDN U33213 ( .B(n26771), .A(n26772), .Z(n26769) );
  AND U33214 ( .A(a[70]), .B(b[15]), .Z(n26768) );
  XOR U33215 ( .A(n26774), .B(n26775), .Z(n26269) );
  ANDN U33216 ( .B(n26776), .A(n26777), .Z(n26774) );
  AND U33217 ( .A(a[71]), .B(b[14]), .Z(n26773) );
  XOR U33218 ( .A(n26779), .B(n26780), .Z(n26274) );
  ANDN U33219 ( .B(n26781), .A(n26782), .Z(n26779) );
  AND U33220 ( .A(a[72]), .B(b[13]), .Z(n26778) );
  XOR U33221 ( .A(n26784), .B(n26785), .Z(n26279) );
  ANDN U33222 ( .B(n26786), .A(n26787), .Z(n26784) );
  AND U33223 ( .A(a[73]), .B(b[12]), .Z(n26783) );
  XOR U33224 ( .A(n26789), .B(n26790), .Z(n26284) );
  ANDN U33225 ( .B(n26791), .A(n26792), .Z(n26789) );
  AND U33226 ( .A(a[74]), .B(b[11]), .Z(n26788) );
  XOR U33227 ( .A(n26794), .B(n26795), .Z(n26289) );
  ANDN U33228 ( .B(n26796), .A(n26797), .Z(n26794) );
  AND U33229 ( .A(a[75]), .B(b[10]), .Z(n26793) );
  XOR U33230 ( .A(n26799), .B(n26800), .Z(n26294) );
  ANDN U33231 ( .B(n26801), .A(n26802), .Z(n26799) );
  AND U33232 ( .A(b[9]), .B(a[76]), .Z(n26798) );
  XOR U33233 ( .A(n26804), .B(n26805), .Z(n26299) );
  ANDN U33234 ( .B(n26806), .A(n26807), .Z(n26804) );
  AND U33235 ( .A(b[8]), .B(a[77]), .Z(n26803) );
  XOR U33236 ( .A(n26809), .B(n26810), .Z(n26304) );
  ANDN U33237 ( .B(n26811), .A(n26812), .Z(n26809) );
  AND U33238 ( .A(b[7]), .B(a[78]), .Z(n26808) );
  XOR U33239 ( .A(n26814), .B(n26815), .Z(n26309) );
  ANDN U33240 ( .B(n26816), .A(n26817), .Z(n26814) );
  AND U33241 ( .A(b[6]), .B(a[79]), .Z(n26813) );
  XOR U33242 ( .A(n26819), .B(n26820), .Z(n26314) );
  ANDN U33243 ( .B(n26821), .A(n26822), .Z(n26819) );
  AND U33244 ( .A(b[5]), .B(a[80]), .Z(n26818) );
  XOR U33245 ( .A(n26824), .B(n26825), .Z(n26319) );
  ANDN U33246 ( .B(n26826), .A(n26827), .Z(n26824) );
  AND U33247 ( .A(b[4]), .B(a[81]), .Z(n26823) );
  XOR U33248 ( .A(n26829), .B(n26830), .Z(n26324) );
  ANDN U33249 ( .B(n26336), .A(n26337), .Z(n26829) );
  AND U33250 ( .A(b[2]), .B(a[82]), .Z(n26831) );
  XNOR U33251 ( .A(n26826), .B(n26830), .Z(n26832) );
  XOR U33252 ( .A(n26833), .B(n26834), .Z(n26830) );
  OR U33253 ( .A(n26339), .B(n26340), .Z(n26834) );
  XNOR U33254 ( .A(n26836), .B(n26837), .Z(n26835) );
  XOR U33255 ( .A(n26836), .B(n26839), .Z(n26339) );
  NAND U33256 ( .A(b[1]), .B(a[82]), .Z(n26839) );
  IV U33257 ( .A(n26833), .Z(n26836) );
  NANDN U33258 ( .A(n39), .B(n40), .Z(n26833) );
  XOR U33259 ( .A(n26840), .B(n26841), .Z(n40) );
  NAND U33260 ( .A(a[82]), .B(b[0]), .Z(n39) );
  XNOR U33261 ( .A(n26821), .B(n26825), .Z(n26842) );
  XNOR U33262 ( .A(n26816), .B(n26820), .Z(n26843) );
  XNOR U33263 ( .A(n26811), .B(n26815), .Z(n26844) );
  XNOR U33264 ( .A(n26806), .B(n26810), .Z(n26845) );
  XNOR U33265 ( .A(n26801), .B(n26805), .Z(n26846) );
  XNOR U33266 ( .A(n26796), .B(n26800), .Z(n26847) );
  XNOR U33267 ( .A(n26791), .B(n26795), .Z(n26848) );
  XNOR U33268 ( .A(n26786), .B(n26790), .Z(n26849) );
  XNOR U33269 ( .A(n26781), .B(n26785), .Z(n26850) );
  XNOR U33270 ( .A(n26776), .B(n26780), .Z(n26851) );
  XNOR U33271 ( .A(n26771), .B(n26775), .Z(n26852) );
  XNOR U33272 ( .A(n26766), .B(n26770), .Z(n26853) );
  XNOR U33273 ( .A(n26761), .B(n26765), .Z(n26854) );
  XNOR U33274 ( .A(n26756), .B(n26760), .Z(n26855) );
  XNOR U33275 ( .A(n26751), .B(n26755), .Z(n26856) );
  XNOR U33276 ( .A(n26746), .B(n26750), .Z(n26857) );
  XNOR U33277 ( .A(n26741), .B(n26745), .Z(n26858) );
  XNOR U33278 ( .A(n26736), .B(n26740), .Z(n26859) );
  XNOR U33279 ( .A(n26731), .B(n26735), .Z(n26860) );
  XNOR U33280 ( .A(n26726), .B(n26730), .Z(n26861) );
  XNOR U33281 ( .A(n26721), .B(n26725), .Z(n26862) );
  XNOR U33282 ( .A(n26716), .B(n26720), .Z(n26863) );
  XNOR U33283 ( .A(n26711), .B(n26715), .Z(n26864) );
  XNOR U33284 ( .A(n26706), .B(n26710), .Z(n26865) );
  XNOR U33285 ( .A(n26701), .B(n26705), .Z(n26866) );
  XNOR U33286 ( .A(n26696), .B(n26700), .Z(n26867) );
  XNOR U33287 ( .A(n26691), .B(n26695), .Z(n26868) );
  XNOR U33288 ( .A(n26686), .B(n26690), .Z(n26869) );
  XNOR U33289 ( .A(n26681), .B(n26685), .Z(n26870) );
  XNOR U33290 ( .A(n26676), .B(n26680), .Z(n26871) );
  XNOR U33291 ( .A(n26671), .B(n26675), .Z(n26872) );
  XNOR U33292 ( .A(n26666), .B(n26670), .Z(n26873) );
  XNOR U33293 ( .A(n26661), .B(n26665), .Z(n26874) );
  XNOR U33294 ( .A(n26656), .B(n26660), .Z(n26875) );
  XNOR U33295 ( .A(n26651), .B(n26655), .Z(n26876) );
  XNOR U33296 ( .A(n26646), .B(n26650), .Z(n26877) );
  XNOR U33297 ( .A(n26641), .B(n26645), .Z(n26878) );
  XNOR U33298 ( .A(n26636), .B(n26640), .Z(n26879) );
  XNOR U33299 ( .A(n26631), .B(n26635), .Z(n26880) );
  XNOR U33300 ( .A(n26626), .B(n26630), .Z(n26881) );
  XNOR U33301 ( .A(n26621), .B(n26625), .Z(n26882) );
  XNOR U33302 ( .A(n26616), .B(n26620), .Z(n26883) );
  XNOR U33303 ( .A(n26611), .B(n26615), .Z(n26884) );
  XNOR U33304 ( .A(n26606), .B(n26610), .Z(n26885) );
  XNOR U33305 ( .A(n26601), .B(n26605), .Z(n26886) );
  XNOR U33306 ( .A(n26596), .B(n26600), .Z(n26887) );
  XNOR U33307 ( .A(n26591), .B(n26595), .Z(n26888) );
  XNOR U33308 ( .A(n26586), .B(n26590), .Z(n26889) );
  XNOR U33309 ( .A(n26581), .B(n26585), .Z(n26890) );
  XNOR U33310 ( .A(n26576), .B(n26580), .Z(n26891) );
  XNOR U33311 ( .A(n26571), .B(n26575), .Z(n26892) );
  XNOR U33312 ( .A(n26566), .B(n26570), .Z(n26893) );
  XNOR U33313 ( .A(n26561), .B(n26565), .Z(n26894) );
  XNOR U33314 ( .A(n26556), .B(n26560), .Z(n26895) );
  XNOR U33315 ( .A(n26551), .B(n26555), .Z(n26896) );
  XNOR U33316 ( .A(n26546), .B(n26550), .Z(n26897) );
  XNOR U33317 ( .A(n26541), .B(n26545), .Z(n26898) );
  XNOR U33318 ( .A(n26536), .B(n26540), .Z(n26899) );
  XNOR U33319 ( .A(n26531), .B(n26535), .Z(n26900) );
  XNOR U33320 ( .A(n26526), .B(n26530), .Z(n26901) );
  XNOR U33321 ( .A(n26521), .B(n26525), .Z(n26902) );
  XNOR U33322 ( .A(n26516), .B(n26520), .Z(n26903) );
  XNOR U33323 ( .A(n26511), .B(n26515), .Z(n26904) );
  XNOR U33324 ( .A(n26506), .B(n26510), .Z(n26905) );
  XNOR U33325 ( .A(n26501), .B(n26505), .Z(n26906) );
  XNOR U33326 ( .A(n26496), .B(n26500), .Z(n26907) );
  XNOR U33327 ( .A(n26491), .B(n26495), .Z(n26908) );
  XNOR U33328 ( .A(n26486), .B(n26490), .Z(n26909) );
  XNOR U33329 ( .A(n26481), .B(n26485), .Z(n26910) );
  XNOR U33330 ( .A(n26476), .B(n26480), .Z(n26911) );
  XNOR U33331 ( .A(n26471), .B(n26475), .Z(n26912) );
  XNOR U33332 ( .A(n26466), .B(n26470), .Z(n26913) );
  XNOR U33333 ( .A(n26914), .B(n26915), .Z(n26466) );
  XNOR U33334 ( .A(n26461), .B(n26465), .Z(n26915) );
  XNOR U33335 ( .A(n26456), .B(n26460), .Z(n26916) );
  XNOR U33336 ( .A(n26917), .B(n26918), .Z(n26456) );
  XNOR U33337 ( .A(n26451), .B(n26455), .Z(n26918) );
  XNOR U33338 ( .A(n26446), .B(n26450), .Z(n26919) );
  XNOR U33339 ( .A(n26441), .B(n26445), .Z(n26920) );
  XNOR U33340 ( .A(n26436), .B(n26440), .Z(n26921) );
  XNOR U33341 ( .A(n26431), .B(n26435), .Z(n26922) );
  XNOR U33342 ( .A(n26426), .B(n26430), .Z(n26923) );
  XOR U33343 ( .A(n26924), .B(n26425), .Z(n26426) );
  AND U33344 ( .A(a[0]), .B(b[84]), .Z(n26924) );
  XNOR U33345 ( .A(n26925), .B(n26425), .Z(n26427) );
  XNOR U33346 ( .A(n26926), .B(n26927), .Z(n26425) );
  ANDN U33347 ( .B(n26928), .A(n26929), .Z(n26926) );
  AND U33348 ( .A(a[1]), .B(b[83]), .Z(n26925) );
  XOR U33349 ( .A(n26931), .B(n26932), .Z(n26430) );
  ANDN U33350 ( .B(n26933), .A(n26934), .Z(n26931) );
  AND U33351 ( .A(a[2]), .B(b[82]), .Z(n26930) );
  XOR U33352 ( .A(n26936), .B(n26937), .Z(n26435) );
  ANDN U33353 ( .B(n26938), .A(n26939), .Z(n26936) );
  AND U33354 ( .A(a[3]), .B(b[81]), .Z(n26935) );
  XOR U33355 ( .A(n26941), .B(n26942), .Z(n26440) );
  ANDN U33356 ( .B(n26943), .A(n26944), .Z(n26941) );
  AND U33357 ( .A(a[4]), .B(b[80]), .Z(n26940) );
  XOR U33358 ( .A(n26946), .B(n26947), .Z(n26445) );
  ANDN U33359 ( .B(n26948), .A(n26949), .Z(n26946) );
  AND U33360 ( .A(a[5]), .B(b[79]), .Z(n26945) );
  IV U33361 ( .A(n26452), .Z(n26917) );
  XOR U33362 ( .A(n26951), .B(n26952), .Z(n26450) );
  ANDN U33363 ( .B(n26953), .A(n26954), .Z(n26951) );
  AND U33364 ( .A(a[6]), .B(b[78]), .Z(n26950) );
  XOR U33365 ( .A(n26956), .B(n26957), .Z(n26455) );
  ANDN U33366 ( .B(n26958), .A(n26959), .Z(n26956) );
  AND U33367 ( .A(a[7]), .B(b[77]), .Z(n26955) );
  IV U33368 ( .A(n26462), .Z(n26914) );
  XOR U33369 ( .A(n26961), .B(n26962), .Z(n26460) );
  ANDN U33370 ( .B(n26963), .A(n26964), .Z(n26961) );
  AND U33371 ( .A(a[8]), .B(b[76]), .Z(n26960) );
  XOR U33372 ( .A(n26966), .B(n26967), .Z(n26465) );
  ANDN U33373 ( .B(n26968), .A(n26969), .Z(n26966) );
  AND U33374 ( .A(a[9]), .B(b[75]), .Z(n26965) );
  XOR U33375 ( .A(n26971), .B(n26972), .Z(n26470) );
  ANDN U33376 ( .B(n26973), .A(n26974), .Z(n26971) );
  AND U33377 ( .A(a[10]), .B(b[74]), .Z(n26970) );
  XOR U33378 ( .A(n26976), .B(n26977), .Z(n26475) );
  ANDN U33379 ( .B(n26978), .A(n26979), .Z(n26976) );
  AND U33380 ( .A(a[11]), .B(b[73]), .Z(n26975) );
  XOR U33381 ( .A(n26981), .B(n26982), .Z(n26480) );
  ANDN U33382 ( .B(n26983), .A(n26984), .Z(n26981) );
  AND U33383 ( .A(a[12]), .B(b[72]), .Z(n26980) );
  XOR U33384 ( .A(n26986), .B(n26987), .Z(n26485) );
  ANDN U33385 ( .B(n26988), .A(n26989), .Z(n26986) );
  AND U33386 ( .A(a[13]), .B(b[71]), .Z(n26985) );
  XOR U33387 ( .A(n26991), .B(n26992), .Z(n26490) );
  ANDN U33388 ( .B(n26993), .A(n26994), .Z(n26991) );
  AND U33389 ( .A(a[14]), .B(b[70]), .Z(n26990) );
  XOR U33390 ( .A(n26996), .B(n26997), .Z(n26495) );
  ANDN U33391 ( .B(n26998), .A(n26999), .Z(n26996) );
  AND U33392 ( .A(a[15]), .B(b[69]), .Z(n26995) );
  XOR U33393 ( .A(n27001), .B(n27002), .Z(n26500) );
  ANDN U33394 ( .B(n27003), .A(n27004), .Z(n27001) );
  AND U33395 ( .A(a[16]), .B(b[68]), .Z(n27000) );
  XOR U33396 ( .A(n27006), .B(n27007), .Z(n26505) );
  ANDN U33397 ( .B(n27008), .A(n27009), .Z(n27006) );
  AND U33398 ( .A(a[17]), .B(b[67]), .Z(n27005) );
  XOR U33399 ( .A(n27011), .B(n27012), .Z(n26510) );
  ANDN U33400 ( .B(n27013), .A(n27014), .Z(n27011) );
  AND U33401 ( .A(a[18]), .B(b[66]), .Z(n27010) );
  XOR U33402 ( .A(n27016), .B(n27017), .Z(n26515) );
  ANDN U33403 ( .B(n27018), .A(n27019), .Z(n27016) );
  AND U33404 ( .A(a[19]), .B(b[65]), .Z(n27015) );
  XOR U33405 ( .A(n27021), .B(n27022), .Z(n26520) );
  ANDN U33406 ( .B(n27023), .A(n27024), .Z(n27021) );
  AND U33407 ( .A(a[20]), .B(b[64]), .Z(n27020) );
  XOR U33408 ( .A(n27026), .B(n27027), .Z(n26525) );
  ANDN U33409 ( .B(n27028), .A(n27029), .Z(n27026) );
  AND U33410 ( .A(a[21]), .B(b[63]), .Z(n27025) );
  XOR U33411 ( .A(n27031), .B(n27032), .Z(n26530) );
  ANDN U33412 ( .B(n27033), .A(n27034), .Z(n27031) );
  AND U33413 ( .A(a[22]), .B(b[62]), .Z(n27030) );
  XOR U33414 ( .A(n27036), .B(n27037), .Z(n26535) );
  ANDN U33415 ( .B(n27038), .A(n27039), .Z(n27036) );
  AND U33416 ( .A(a[23]), .B(b[61]), .Z(n27035) );
  XOR U33417 ( .A(n27041), .B(n27042), .Z(n26540) );
  ANDN U33418 ( .B(n27043), .A(n27044), .Z(n27041) );
  AND U33419 ( .A(a[24]), .B(b[60]), .Z(n27040) );
  XOR U33420 ( .A(n27046), .B(n27047), .Z(n26545) );
  ANDN U33421 ( .B(n27048), .A(n27049), .Z(n27046) );
  AND U33422 ( .A(a[25]), .B(b[59]), .Z(n27045) );
  XOR U33423 ( .A(n27051), .B(n27052), .Z(n26550) );
  ANDN U33424 ( .B(n27053), .A(n27054), .Z(n27051) );
  AND U33425 ( .A(a[26]), .B(b[58]), .Z(n27050) );
  XOR U33426 ( .A(n27056), .B(n27057), .Z(n26555) );
  ANDN U33427 ( .B(n27058), .A(n27059), .Z(n27056) );
  AND U33428 ( .A(a[27]), .B(b[57]), .Z(n27055) );
  XOR U33429 ( .A(n27061), .B(n27062), .Z(n26560) );
  ANDN U33430 ( .B(n27063), .A(n27064), .Z(n27061) );
  AND U33431 ( .A(a[28]), .B(b[56]), .Z(n27060) );
  XOR U33432 ( .A(n27066), .B(n27067), .Z(n26565) );
  ANDN U33433 ( .B(n27068), .A(n27069), .Z(n27066) );
  AND U33434 ( .A(a[29]), .B(b[55]), .Z(n27065) );
  XOR U33435 ( .A(n27071), .B(n27072), .Z(n26570) );
  ANDN U33436 ( .B(n27073), .A(n27074), .Z(n27071) );
  AND U33437 ( .A(a[30]), .B(b[54]), .Z(n27070) );
  XOR U33438 ( .A(n27076), .B(n27077), .Z(n26575) );
  ANDN U33439 ( .B(n27078), .A(n27079), .Z(n27076) );
  AND U33440 ( .A(a[31]), .B(b[53]), .Z(n27075) );
  XOR U33441 ( .A(n27081), .B(n27082), .Z(n26580) );
  ANDN U33442 ( .B(n27083), .A(n27084), .Z(n27081) );
  AND U33443 ( .A(a[32]), .B(b[52]), .Z(n27080) );
  XOR U33444 ( .A(n27086), .B(n27087), .Z(n26585) );
  ANDN U33445 ( .B(n27088), .A(n27089), .Z(n27086) );
  AND U33446 ( .A(a[33]), .B(b[51]), .Z(n27085) );
  XOR U33447 ( .A(n27091), .B(n27092), .Z(n26590) );
  ANDN U33448 ( .B(n27093), .A(n27094), .Z(n27091) );
  AND U33449 ( .A(a[34]), .B(b[50]), .Z(n27090) );
  XOR U33450 ( .A(n27096), .B(n27097), .Z(n26595) );
  ANDN U33451 ( .B(n27098), .A(n27099), .Z(n27096) );
  AND U33452 ( .A(a[35]), .B(b[49]), .Z(n27095) );
  XOR U33453 ( .A(n27101), .B(n27102), .Z(n26600) );
  ANDN U33454 ( .B(n27103), .A(n27104), .Z(n27101) );
  AND U33455 ( .A(a[36]), .B(b[48]), .Z(n27100) );
  XOR U33456 ( .A(n27106), .B(n27107), .Z(n26605) );
  ANDN U33457 ( .B(n27108), .A(n27109), .Z(n27106) );
  AND U33458 ( .A(a[37]), .B(b[47]), .Z(n27105) );
  XOR U33459 ( .A(n27111), .B(n27112), .Z(n26610) );
  ANDN U33460 ( .B(n27113), .A(n27114), .Z(n27111) );
  AND U33461 ( .A(a[38]), .B(b[46]), .Z(n27110) );
  XOR U33462 ( .A(n27116), .B(n27117), .Z(n26615) );
  ANDN U33463 ( .B(n27118), .A(n27119), .Z(n27116) );
  AND U33464 ( .A(a[39]), .B(b[45]), .Z(n27115) );
  XOR U33465 ( .A(n27121), .B(n27122), .Z(n26620) );
  ANDN U33466 ( .B(n27123), .A(n27124), .Z(n27121) );
  AND U33467 ( .A(a[40]), .B(b[44]), .Z(n27120) );
  XOR U33468 ( .A(n27126), .B(n27127), .Z(n26625) );
  ANDN U33469 ( .B(n27128), .A(n27129), .Z(n27126) );
  AND U33470 ( .A(a[41]), .B(b[43]), .Z(n27125) );
  XOR U33471 ( .A(n27131), .B(n27132), .Z(n26630) );
  ANDN U33472 ( .B(n27133), .A(n27134), .Z(n27131) );
  AND U33473 ( .A(a[42]), .B(b[42]), .Z(n27130) );
  XOR U33474 ( .A(n27136), .B(n27137), .Z(n26635) );
  ANDN U33475 ( .B(n27138), .A(n27139), .Z(n27136) );
  AND U33476 ( .A(a[43]), .B(b[41]), .Z(n27135) );
  XOR U33477 ( .A(n27141), .B(n27142), .Z(n26640) );
  ANDN U33478 ( .B(n27143), .A(n27144), .Z(n27141) );
  AND U33479 ( .A(a[44]), .B(b[40]), .Z(n27140) );
  XOR U33480 ( .A(n27146), .B(n27147), .Z(n26645) );
  ANDN U33481 ( .B(n27148), .A(n27149), .Z(n27146) );
  AND U33482 ( .A(a[45]), .B(b[39]), .Z(n27145) );
  XOR U33483 ( .A(n27151), .B(n27152), .Z(n26650) );
  ANDN U33484 ( .B(n27153), .A(n27154), .Z(n27151) );
  AND U33485 ( .A(a[46]), .B(b[38]), .Z(n27150) );
  XOR U33486 ( .A(n27156), .B(n27157), .Z(n26655) );
  ANDN U33487 ( .B(n27158), .A(n27159), .Z(n27156) );
  AND U33488 ( .A(a[47]), .B(b[37]), .Z(n27155) );
  XOR U33489 ( .A(n27161), .B(n27162), .Z(n26660) );
  ANDN U33490 ( .B(n27163), .A(n27164), .Z(n27161) );
  AND U33491 ( .A(a[48]), .B(b[36]), .Z(n27160) );
  XOR U33492 ( .A(n27166), .B(n27167), .Z(n26665) );
  ANDN U33493 ( .B(n27168), .A(n27169), .Z(n27166) );
  AND U33494 ( .A(a[49]), .B(b[35]), .Z(n27165) );
  XOR U33495 ( .A(n27171), .B(n27172), .Z(n26670) );
  ANDN U33496 ( .B(n27173), .A(n27174), .Z(n27171) );
  AND U33497 ( .A(a[50]), .B(b[34]), .Z(n27170) );
  XOR U33498 ( .A(n27176), .B(n27177), .Z(n26675) );
  ANDN U33499 ( .B(n27178), .A(n27179), .Z(n27176) );
  AND U33500 ( .A(a[51]), .B(b[33]), .Z(n27175) );
  XOR U33501 ( .A(n27181), .B(n27182), .Z(n26680) );
  ANDN U33502 ( .B(n27183), .A(n27184), .Z(n27181) );
  AND U33503 ( .A(a[52]), .B(b[32]), .Z(n27180) );
  XOR U33504 ( .A(n27186), .B(n27187), .Z(n26685) );
  ANDN U33505 ( .B(n27188), .A(n27189), .Z(n27186) );
  AND U33506 ( .A(a[53]), .B(b[31]), .Z(n27185) );
  XOR U33507 ( .A(n27191), .B(n27192), .Z(n26690) );
  ANDN U33508 ( .B(n27193), .A(n27194), .Z(n27191) );
  AND U33509 ( .A(a[54]), .B(b[30]), .Z(n27190) );
  XOR U33510 ( .A(n27196), .B(n27197), .Z(n26695) );
  ANDN U33511 ( .B(n27198), .A(n27199), .Z(n27196) );
  AND U33512 ( .A(a[55]), .B(b[29]), .Z(n27195) );
  XOR U33513 ( .A(n27201), .B(n27202), .Z(n26700) );
  ANDN U33514 ( .B(n27203), .A(n27204), .Z(n27201) );
  AND U33515 ( .A(a[56]), .B(b[28]), .Z(n27200) );
  XOR U33516 ( .A(n27206), .B(n27207), .Z(n26705) );
  ANDN U33517 ( .B(n27208), .A(n27209), .Z(n27206) );
  AND U33518 ( .A(a[57]), .B(b[27]), .Z(n27205) );
  XOR U33519 ( .A(n27211), .B(n27212), .Z(n26710) );
  ANDN U33520 ( .B(n27213), .A(n27214), .Z(n27211) );
  AND U33521 ( .A(a[58]), .B(b[26]), .Z(n27210) );
  XOR U33522 ( .A(n27216), .B(n27217), .Z(n26715) );
  ANDN U33523 ( .B(n27218), .A(n27219), .Z(n27216) );
  AND U33524 ( .A(a[59]), .B(b[25]), .Z(n27215) );
  XOR U33525 ( .A(n27221), .B(n27222), .Z(n26720) );
  ANDN U33526 ( .B(n27223), .A(n27224), .Z(n27221) );
  AND U33527 ( .A(a[60]), .B(b[24]), .Z(n27220) );
  XOR U33528 ( .A(n27226), .B(n27227), .Z(n26725) );
  ANDN U33529 ( .B(n27228), .A(n27229), .Z(n27226) );
  AND U33530 ( .A(a[61]), .B(b[23]), .Z(n27225) );
  XOR U33531 ( .A(n27231), .B(n27232), .Z(n26730) );
  ANDN U33532 ( .B(n27233), .A(n27234), .Z(n27231) );
  AND U33533 ( .A(a[62]), .B(b[22]), .Z(n27230) );
  XOR U33534 ( .A(n27236), .B(n27237), .Z(n26735) );
  ANDN U33535 ( .B(n27238), .A(n27239), .Z(n27236) );
  AND U33536 ( .A(a[63]), .B(b[21]), .Z(n27235) );
  XOR U33537 ( .A(n27241), .B(n27242), .Z(n26740) );
  ANDN U33538 ( .B(n27243), .A(n27244), .Z(n27241) );
  AND U33539 ( .A(a[64]), .B(b[20]), .Z(n27240) );
  XOR U33540 ( .A(n27246), .B(n27247), .Z(n26745) );
  ANDN U33541 ( .B(n27248), .A(n27249), .Z(n27246) );
  AND U33542 ( .A(a[65]), .B(b[19]), .Z(n27245) );
  XOR U33543 ( .A(n27251), .B(n27252), .Z(n26750) );
  ANDN U33544 ( .B(n27253), .A(n27254), .Z(n27251) );
  AND U33545 ( .A(a[66]), .B(b[18]), .Z(n27250) );
  XOR U33546 ( .A(n27256), .B(n27257), .Z(n26755) );
  ANDN U33547 ( .B(n27258), .A(n27259), .Z(n27256) );
  AND U33548 ( .A(a[67]), .B(b[17]), .Z(n27255) );
  XOR U33549 ( .A(n27261), .B(n27262), .Z(n26760) );
  ANDN U33550 ( .B(n27263), .A(n27264), .Z(n27261) );
  AND U33551 ( .A(a[68]), .B(b[16]), .Z(n27260) );
  XOR U33552 ( .A(n27266), .B(n27267), .Z(n26765) );
  ANDN U33553 ( .B(n27268), .A(n27269), .Z(n27266) );
  AND U33554 ( .A(a[69]), .B(b[15]), .Z(n27265) );
  XOR U33555 ( .A(n27271), .B(n27272), .Z(n26770) );
  ANDN U33556 ( .B(n27273), .A(n27274), .Z(n27271) );
  AND U33557 ( .A(a[70]), .B(b[14]), .Z(n27270) );
  XOR U33558 ( .A(n27276), .B(n27277), .Z(n26775) );
  ANDN U33559 ( .B(n27278), .A(n27279), .Z(n27276) );
  AND U33560 ( .A(a[71]), .B(b[13]), .Z(n27275) );
  XOR U33561 ( .A(n27281), .B(n27282), .Z(n26780) );
  ANDN U33562 ( .B(n27283), .A(n27284), .Z(n27281) );
  AND U33563 ( .A(a[72]), .B(b[12]), .Z(n27280) );
  XOR U33564 ( .A(n27286), .B(n27287), .Z(n26785) );
  ANDN U33565 ( .B(n27288), .A(n27289), .Z(n27286) );
  AND U33566 ( .A(a[73]), .B(b[11]), .Z(n27285) );
  XOR U33567 ( .A(n27291), .B(n27292), .Z(n26790) );
  ANDN U33568 ( .B(n27293), .A(n27294), .Z(n27291) );
  AND U33569 ( .A(a[74]), .B(b[10]), .Z(n27290) );
  XOR U33570 ( .A(n27296), .B(n27297), .Z(n26795) );
  ANDN U33571 ( .B(n27298), .A(n27299), .Z(n27296) );
  AND U33572 ( .A(b[9]), .B(a[75]), .Z(n27295) );
  XOR U33573 ( .A(n27301), .B(n27302), .Z(n26800) );
  ANDN U33574 ( .B(n27303), .A(n27304), .Z(n27301) );
  AND U33575 ( .A(b[8]), .B(a[76]), .Z(n27300) );
  XOR U33576 ( .A(n27306), .B(n27307), .Z(n26805) );
  ANDN U33577 ( .B(n27308), .A(n27309), .Z(n27306) );
  AND U33578 ( .A(b[7]), .B(a[77]), .Z(n27305) );
  XOR U33579 ( .A(n27311), .B(n27312), .Z(n26810) );
  ANDN U33580 ( .B(n27313), .A(n27314), .Z(n27311) );
  AND U33581 ( .A(b[6]), .B(a[78]), .Z(n27310) );
  XOR U33582 ( .A(n27316), .B(n27317), .Z(n26815) );
  ANDN U33583 ( .B(n27318), .A(n27319), .Z(n27316) );
  AND U33584 ( .A(b[5]), .B(a[79]), .Z(n27315) );
  XOR U33585 ( .A(n27321), .B(n27322), .Z(n26820) );
  ANDN U33586 ( .B(n27323), .A(n27324), .Z(n27321) );
  AND U33587 ( .A(b[4]), .B(a[80]), .Z(n27320) );
  XOR U33588 ( .A(n27326), .B(n27327), .Z(n26825) );
  ANDN U33589 ( .B(n26837), .A(n26838), .Z(n27326) );
  AND U33590 ( .A(b[2]), .B(a[81]), .Z(n27328) );
  XNOR U33591 ( .A(n27323), .B(n27327), .Z(n27329) );
  XOR U33592 ( .A(n27330), .B(n27331), .Z(n27327) );
  OR U33593 ( .A(n26840), .B(n26841), .Z(n27331) );
  XNOR U33594 ( .A(n27333), .B(n27334), .Z(n27332) );
  XOR U33595 ( .A(n27333), .B(n27336), .Z(n26840) );
  NAND U33596 ( .A(b[1]), .B(a[81]), .Z(n27336) );
  IV U33597 ( .A(n27330), .Z(n27333) );
  NANDN U33598 ( .A(n41), .B(n42), .Z(n27330) );
  XOR U33599 ( .A(n27337), .B(n27338), .Z(n42) );
  NAND U33600 ( .A(a[81]), .B(b[0]), .Z(n41) );
  XNOR U33601 ( .A(n27318), .B(n27322), .Z(n27339) );
  XNOR U33602 ( .A(n27313), .B(n27317), .Z(n27340) );
  XNOR U33603 ( .A(n27308), .B(n27312), .Z(n27341) );
  XNOR U33604 ( .A(n27303), .B(n27307), .Z(n27342) );
  XNOR U33605 ( .A(n27298), .B(n27302), .Z(n27343) );
  XNOR U33606 ( .A(n27293), .B(n27297), .Z(n27344) );
  XNOR U33607 ( .A(n27288), .B(n27292), .Z(n27345) );
  XNOR U33608 ( .A(n27283), .B(n27287), .Z(n27346) );
  XNOR U33609 ( .A(n27278), .B(n27282), .Z(n27347) );
  XNOR U33610 ( .A(n27273), .B(n27277), .Z(n27348) );
  XNOR U33611 ( .A(n27268), .B(n27272), .Z(n27349) );
  XNOR U33612 ( .A(n27263), .B(n27267), .Z(n27350) );
  XNOR U33613 ( .A(n27258), .B(n27262), .Z(n27351) );
  XNOR U33614 ( .A(n27253), .B(n27257), .Z(n27352) );
  XNOR U33615 ( .A(n27248), .B(n27252), .Z(n27353) );
  XNOR U33616 ( .A(n27243), .B(n27247), .Z(n27354) );
  XNOR U33617 ( .A(n27238), .B(n27242), .Z(n27355) );
  XNOR U33618 ( .A(n27233), .B(n27237), .Z(n27356) );
  XNOR U33619 ( .A(n27228), .B(n27232), .Z(n27357) );
  XNOR U33620 ( .A(n27223), .B(n27227), .Z(n27358) );
  XNOR U33621 ( .A(n27218), .B(n27222), .Z(n27359) );
  XNOR U33622 ( .A(n27213), .B(n27217), .Z(n27360) );
  XNOR U33623 ( .A(n27208), .B(n27212), .Z(n27361) );
  XNOR U33624 ( .A(n27203), .B(n27207), .Z(n27362) );
  XNOR U33625 ( .A(n27198), .B(n27202), .Z(n27363) );
  XNOR U33626 ( .A(n27193), .B(n27197), .Z(n27364) );
  XNOR U33627 ( .A(n27188), .B(n27192), .Z(n27365) );
  XNOR U33628 ( .A(n27183), .B(n27187), .Z(n27366) );
  XNOR U33629 ( .A(n27178), .B(n27182), .Z(n27367) );
  XNOR U33630 ( .A(n27173), .B(n27177), .Z(n27368) );
  XNOR U33631 ( .A(n27168), .B(n27172), .Z(n27369) );
  XNOR U33632 ( .A(n27163), .B(n27167), .Z(n27370) );
  XNOR U33633 ( .A(n27158), .B(n27162), .Z(n27371) );
  XNOR U33634 ( .A(n27153), .B(n27157), .Z(n27372) );
  XNOR U33635 ( .A(n27148), .B(n27152), .Z(n27373) );
  XNOR U33636 ( .A(n27143), .B(n27147), .Z(n27374) );
  XNOR U33637 ( .A(n27138), .B(n27142), .Z(n27375) );
  XNOR U33638 ( .A(n27133), .B(n27137), .Z(n27376) );
  XNOR U33639 ( .A(n27128), .B(n27132), .Z(n27377) );
  XNOR U33640 ( .A(n27123), .B(n27127), .Z(n27378) );
  XNOR U33641 ( .A(n27118), .B(n27122), .Z(n27379) );
  XNOR U33642 ( .A(n27113), .B(n27117), .Z(n27380) );
  XNOR U33643 ( .A(n27108), .B(n27112), .Z(n27381) );
  XNOR U33644 ( .A(n27103), .B(n27107), .Z(n27382) );
  XNOR U33645 ( .A(n27098), .B(n27102), .Z(n27383) );
  XNOR U33646 ( .A(n27093), .B(n27097), .Z(n27384) );
  XNOR U33647 ( .A(n27088), .B(n27092), .Z(n27385) );
  XNOR U33648 ( .A(n27083), .B(n27087), .Z(n27386) );
  XNOR U33649 ( .A(n27078), .B(n27082), .Z(n27387) );
  XNOR U33650 ( .A(n27073), .B(n27077), .Z(n27388) );
  XNOR U33651 ( .A(n27068), .B(n27072), .Z(n27389) );
  XNOR U33652 ( .A(n27063), .B(n27067), .Z(n27390) );
  XNOR U33653 ( .A(n27058), .B(n27062), .Z(n27391) );
  XNOR U33654 ( .A(n27053), .B(n27057), .Z(n27392) );
  XNOR U33655 ( .A(n27048), .B(n27052), .Z(n27393) );
  XNOR U33656 ( .A(n27043), .B(n27047), .Z(n27394) );
  XNOR U33657 ( .A(n27038), .B(n27042), .Z(n27395) );
  XNOR U33658 ( .A(n27033), .B(n27037), .Z(n27396) );
  XNOR U33659 ( .A(n27028), .B(n27032), .Z(n27397) );
  XNOR U33660 ( .A(n27023), .B(n27027), .Z(n27398) );
  XNOR U33661 ( .A(n27018), .B(n27022), .Z(n27399) );
  XNOR U33662 ( .A(n27013), .B(n27017), .Z(n27400) );
  XNOR U33663 ( .A(n27008), .B(n27012), .Z(n27401) );
  XNOR U33664 ( .A(n27003), .B(n27007), .Z(n27402) );
  XNOR U33665 ( .A(n26998), .B(n27002), .Z(n27403) );
  XNOR U33666 ( .A(n26993), .B(n26997), .Z(n27404) );
  XNOR U33667 ( .A(n26988), .B(n26992), .Z(n27405) );
  XNOR U33668 ( .A(n26983), .B(n26987), .Z(n27406) );
  XNOR U33669 ( .A(n26978), .B(n26982), .Z(n27407) );
  XNOR U33670 ( .A(n26973), .B(n26977), .Z(n27408) );
  XNOR U33671 ( .A(n26968), .B(n26972), .Z(n27409) );
  XNOR U33672 ( .A(n26963), .B(n26967), .Z(n27410) );
  XNOR U33673 ( .A(n26958), .B(n26962), .Z(n27411) );
  XNOR U33674 ( .A(n26953), .B(n26957), .Z(n27412) );
  XNOR U33675 ( .A(n26948), .B(n26952), .Z(n27413) );
  XNOR U33676 ( .A(n26943), .B(n26947), .Z(n27414) );
  XNOR U33677 ( .A(n26938), .B(n26942), .Z(n27415) );
  XNOR U33678 ( .A(n26933), .B(n26937), .Z(n27416) );
  XNOR U33679 ( .A(n26928), .B(n26932), .Z(n27417) );
  XNOR U33680 ( .A(n27418), .B(n26927), .Z(n26928) );
  AND U33681 ( .A(a[0]), .B(b[83]), .Z(n27418) );
  XOR U33682 ( .A(n27419), .B(n26927), .Z(n26929) );
  XNOR U33683 ( .A(n27420), .B(n27421), .Z(n26927) );
  ANDN U33684 ( .B(n27422), .A(n27423), .Z(n27420) );
  AND U33685 ( .A(a[1]), .B(b[82]), .Z(n27419) );
  XOR U33686 ( .A(n27425), .B(n27426), .Z(n26932) );
  ANDN U33687 ( .B(n27427), .A(n27428), .Z(n27425) );
  AND U33688 ( .A(a[2]), .B(b[81]), .Z(n27424) );
  XOR U33689 ( .A(n27430), .B(n27431), .Z(n26937) );
  ANDN U33690 ( .B(n27432), .A(n27433), .Z(n27430) );
  AND U33691 ( .A(a[3]), .B(b[80]), .Z(n27429) );
  XOR U33692 ( .A(n27435), .B(n27436), .Z(n26942) );
  ANDN U33693 ( .B(n27437), .A(n27438), .Z(n27435) );
  AND U33694 ( .A(a[4]), .B(b[79]), .Z(n27434) );
  XOR U33695 ( .A(n27440), .B(n27441), .Z(n26947) );
  ANDN U33696 ( .B(n27442), .A(n27443), .Z(n27440) );
  AND U33697 ( .A(a[5]), .B(b[78]), .Z(n27439) );
  XOR U33698 ( .A(n27445), .B(n27446), .Z(n26952) );
  ANDN U33699 ( .B(n27447), .A(n27448), .Z(n27445) );
  AND U33700 ( .A(a[6]), .B(b[77]), .Z(n27444) );
  XOR U33701 ( .A(n27450), .B(n27451), .Z(n26957) );
  ANDN U33702 ( .B(n27452), .A(n27453), .Z(n27450) );
  AND U33703 ( .A(a[7]), .B(b[76]), .Z(n27449) );
  XOR U33704 ( .A(n27455), .B(n27456), .Z(n26962) );
  ANDN U33705 ( .B(n27457), .A(n27458), .Z(n27455) );
  AND U33706 ( .A(a[8]), .B(b[75]), .Z(n27454) );
  XOR U33707 ( .A(n27460), .B(n27461), .Z(n26967) );
  ANDN U33708 ( .B(n27462), .A(n27463), .Z(n27460) );
  AND U33709 ( .A(a[9]), .B(b[74]), .Z(n27459) );
  XOR U33710 ( .A(n27465), .B(n27466), .Z(n26972) );
  ANDN U33711 ( .B(n27467), .A(n27468), .Z(n27465) );
  AND U33712 ( .A(a[10]), .B(b[73]), .Z(n27464) );
  XOR U33713 ( .A(n27470), .B(n27471), .Z(n26977) );
  ANDN U33714 ( .B(n27472), .A(n27473), .Z(n27470) );
  AND U33715 ( .A(a[11]), .B(b[72]), .Z(n27469) );
  XOR U33716 ( .A(n27475), .B(n27476), .Z(n26982) );
  ANDN U33717 ( .B(n27477), .A(n27478), .Z(n27475) );
  AND U33718 ( .A(a[12]), .B(b[71]), .Z(n27474) );
  XOR U33719 ( .A(n27480), .B(n27481), .Z(n26987) );
  ANDN U33720 ( .B(n27482), .A(n27483), .Z(n27480) );
  AND U33721 ( .A(a[13]), .B(b[70]), .Z(n27479) );
  XOR U33722 ( .A(n27485), .B(n27486), .Z(n26992) );
  ANDN U33723 ( .B(n27487), .A(n27488), .Z(n27485) );
  AND U33724 ( .A(a[14]), .B(b[69]), .Z(n27484) );
  XOR U33725 ( .A(n27490), .B(n27491), .Z(n26997) );
  ANDN U33726 ( .B(n27492), .A(n27493), .Z(n27490) );
  AND U33727 ( .A(a[15]), .B(b[68]), .Z(n27489) );
  XOR U33728 ( .A(n27495), .B(n27496), .Z(n27002) );
  ANDN U33729 ( .B(n27497), .A(n27498), .Z(n27495) );
  AND U33730 ( .A(a[16]), .B(b[67]), .Z(n27494) );
  XOR U33731 ( .A(n27500), .B(n27501), .Z(n27007) );
  ANDN U33732 ( .B(n27502), .A(n27503), .Z(n27500) );
  AND U33733 ( .A(a[17]), .B(b[66]), .Z(n27499) );
  XOR U33734 ( .A(n27505), .B(n27506), .Z(n27012) );
  ANDN U33735 ( .B(n27507), .A(n27508), .Z(n27505) );
  AND U33736 ( .A(a[18]), .B(b[65]), .Z(n27504) );
  XOR U33737 ( .A(n27510), .B(n27511), .Z(n27017) );
  ANDN U33738 ( .B(n27512), .A(n27513), .Z(n27510) );
  AND U33739 ( .A(a[19]), .B(b[64]), .Z(n27509) );
  XOR U33740 ( .A(n27515), .B(n27516), .Z(n27022) );
  ANDN U33741 ( .B(n27517), .A(n27518), .Z(n27515) );
  AND U33742 ( .A(a[20]), .B(b[63]), .Z(n27514) );
  XOR U33743 ( .A(n27520), .B(n27521), .Z(n27027) );
  ANDN U33744 ( .B(n27522), .A(n27523), .Z(n27520) );
  AND U33745 ( .A(a[21]), .B(b[62]), .Z(n27519) );
  XOR U33746 ( .A(n27525), .B(n27526), .Z(n27032) );
  ANDN U33747 ( .B(n27527), .A(n27528), .Z(n27525) );
  AND U33748 ( .A(a[22]), .B(b[61]), .Z(n27524) );
  XOR U33749 ( .A(n27530), .B(n27531), .Z(n27037) );
  ANDN U33750 ( .B(n27532), .A(n27533), .Z(n27530) );
  AND U33751 ( .A(a[23]), .B(b[60]), .Z(n27529) );
  XOR U33752 ( .A(n27535), .B(n27536), .Z(n27042) );
  ANDN U33753 ( .B(n27537), .A(n27538), .Z(n27535) );
  AND U33754 ( .A(a[24]), .B(b[59]), .Z(n27534) );
  XOR U33755 ( .A(n27540), .B(n27541), .Z(n27047) );
  ANDN U33756 ( .B(n27542), .A(n27543), .Z(n27540) );
  AND U33757 ( .A(a[25]), .B(b[58]), .Z(n27539) );
  XOR U33758 ( .A(n27545), .B(n27546), .Z(n27052) );
  ANDN U33759 ( .B(n27547), .A(n27548), .Z(n27545) );
  AND U33760 ( .A(a[26]), .B(b[57]), .Z(n27544) );
  XOR U33761 ( .A(n27550), .B(n27551), .Z(n27057) );
  ANDN U33762 ( .B(n27552), .A(n27553), .Z(n27550) );
  AND U33763 ( .A(a[27]), .B(b[56]), .Z(n27549) );
  XOR U33764 ( .A(n27555), .B(n27556), .Z(n27062) );
  ANDN U33765 ( .B(n27557), .A(n27558), .Z(n27555) );
  AND U33766 ( .A(a[28]), .B(b[55]), .Z(n27554) );
  XOR U33767 ( .A(n27560), .B(n27561), .Z(n27067) );
  ANDN U33768 ( .B(n27562), .A(n27563), .Z(n27560) );
  AND U33769 ( .A(a[29]), .B(b[54]), .Z(n27559) );
  XOR U33770 ( .A(n27565), .B(n27566), .Z(n27072) );
  ANDN U33771 ( .B(n27567), .A(n27568), .Z(n27565) );
  AND U33772 ( .A(a[30]), .B(b[53]), .Z(n27564) );
  XOR U33773 ( .A(n27570), .B(n27571), .Z(n27077) );
  ANDN U33774 ( .B(n27572), .A(n27573), .Z(n27570) );
  AND U33775 ( .A(a[31]), .B(b[52]), .Z(n27569) );
  XOR U33776 ( .A(n27575), .B(n27576), .Z(n27082) );
  ANDN U33777 ( .B(n27577), .A(n27578), .Z(n27575) );
  AND U33778 ( .A(a[32]), .B(b[51]), .Z(n27574) );
  XOR U33779 ( .A(n27580), .B(n27581), .Z(n27087) );
  ANDN U33780 ( .B(n27582), .A(n27583), .Z(n27580) );
  AND U33781 ( .A(a[33]), .B(b[50]), .Z(n27579) );
  XOR U33782 ( .A(n27585), .B(n27586), .Z(n27092) );
  ANDN U33783 ( .B(n27587), .A(n27588), .Z(n27585) );
  AND U33784 ( .A(a[34]), .B(b[49]), .Z(n27584) );
  XOR U33785 ( .A(n27590), .B(n27591), .Z(n27097) );
  ANDN U33786 ( .B(n27592), .A(n27593), .Z(n27590) );
  AND U33787 ( .A(a[35]), .B(b[48]), .Z(n27589) );
  XOR U33788 ( .A(n27595), .B(n27596), .Z(n27102) );
  ANDN U33789 ( .B(n27597), .A(n27598), .Z(n27595) );
  AND U33790 ( .A(a[36]), .B(b[47]), .Z(n27594) );
  XOR U33791 ( .A(n27600), .B(n27601), .Z(n27107) );
  ANDN U33792 ( .B(n27602), .A(n27603), .Z(n27600) );
  AND U33793 ( .A(a[37]), .B(b[46]), .Z(n27599) );
  XOR U33794 ( .A(n27605), .B(n27606), .Z(n27112) );
  ANDN U33795 ( .B(n27607), .A(n27608), .Z(n27605) );
  AND U33796 ( .A(a[38]), .B(b[45]), .Z(n27604) );
  XOR U33797 ( .A(n27610), .B(n27611), .Z(n27117) );
  ANDN U33798 ( .B(n27612), .A(n27613), .Z(n27610) );
  AND U33799 ( .A(a[39]), .B(b[44]), .Z(n27609) );
  XOR U33800 ( .A(n27615), .B(n27616), .Z(n27122) );
  ANDN U33801 ( .B(n27617), .A(n27618), .Z(n27615) );
  AND U33802 ( .A(a[40]), .B(b[43]), .Z(n27614) );
  XOR U33803 ( .A(n27620), .B(n27621), .Z(n27127) );
  ANDN U33804 ( .B(n27622), .A(n27623), .Z(n27620) );
  AND U33805 ( .A(a[41]), .B(b[42]), .Z(n27619) );
  XOR U33806 ( .A(n27625), .B(n27626), .Z(n27132) );
  ANDN U33807 ( .B(n27627), .A(n27628), .Z(n27625) );
  AND U33808 ( .A(a[42]), .B(b[41]), .Z(n27624) );
  XOR U33809 ( .A(n27630), .B(n27631), .Z(n27137) );
  ANDN U33810 ( .B(n27632), .A(n27633), .Z(n27630) );
  AND U33811 ( .A(a[43]), .B(b[40]), .Z(n27629) );
  XOR U33812 ( .A(n27635), .B(n27636), .Z(n27142) );
  ANDN U33813 ( .B(n27637), .A(n27638), .Z(n27635) );
  AND U33814 ( .A(a[44]), .B(b[39]), .Z(n27634) );
  XOR U33815 ( .A(n27640), .B(n27641), .Z(n27147) );
  ANDN U33816 ( .B(n27642), .A(n27643), .Z(n27640) );
  AND U33817 ( .A(a[45]), .B(b[38]), .Z(n27639) );
  XOR U33818 ( .A(n27645), .B(n27646), .Z(n27152) );
  ANDN U33819 ( .B(n27647), .A(n27648), .Z(n27645) );
  AND U33820 ( .A(a[46]), .B(b[37]), .Z(n27644) );
  XOR U33821 ( .A(n27650), .B(n27651), .Z(n27157) );
  ANDN U33822 ( .B(n27652), .A(n27653), .Z(n27650) );
  AND U33823 ( .A(a[47]), .B(b[36]), .Z(n27649) );
  XOR U33824 ( .A(n27655), .B(n27656), .Z(n27162) );
  ANDN U33825 ( .B(n27657), .A(n27658), .Z(n27655) );
  AND U33826 ( .A(a[48]), .B(b[35]), .Z(n27654) );
  XOR U33827 ( .A(n27660), .B(n27661), .Z(n27167) );
  ANDN U33828 ( .B(n27662), .A(n27663), .Z(n27660) );
  AND U33829 ( .A(a[49]), .B(b[34]), .Z(n27659) );
  XOR U33830 ( .A(n27665), .B(n27666), .Z(n27172) );
  ANDN U33831 ( .B(n27667), .A(n27668), .Z(n27665) );
  AND U33832 ( .A(a[50]), .B(b[33]), .Z(n27664) );
  XOR U33833 ( .A(n27670), .B(n27671), .Z(n27177) );
  ANDN U33834 ( .B(n27672), .A(n27673), .Z(n27670) );
  AND U33835 ( .A(a[51]), .B(b[32]), .Z(n27669) );
  XOR U33836 ( .A(n27675), .B(n27676), .Z(n27182) );
  ANDN U33837 ( .B(n27677), .A(n27678), .Z(n27675) );
  AND U33838 ( .A(a[52]), .B(b[31]), .Z(n27674) );
  XOR U33839 ( .A(n27680), .B(n27681), .Z(n27187) );
  ANDN U33840 ( .B(n27682), .A(n27683), .Z(n27680) );
  AND U33841 ( .A(a[53]), .B(b[30]), .Z(n27679) );
  XOR U33842 ( .A(n27685), .B(n27686), .Z(n27192) );
  ANDN U33843 ( .B(n27687), .A(n27688), .Z(n27685) );
  AND U33844 ( .A(a[54]), .B(b[29]), .Z(n27684) );
  XOR U33845 ( .A(n27690), .B(n27691), .Z(n27197) );
  ANDN U33846 ( .B(n27692), .A(n27693), .Z(n27690) );
  AND U33847 ( .A(a[55]), .B(b[28]), .Z(n27689) );
  XOR U33848 ( .A(n27695), .B(n27696), .Z(n27202) );
  ANDN U33849 ( .B(n27697), .A(n27698), .Z(n27695) );
  AND U33850 ( .A(a[56]), .B(b[27]), .Z(n27694) );
  XOR U33851 ( .A(n27700), .B(n27701), .Z(n27207) );
  ANDN U33852 ( .B(n27702), .A(n27703), .Z(n27700) );
  AND U33853 ( .A(a[57]), .B(b[26]), .Z(n27699) );
  XOR U33854 ( .A(n27705), .B(n27706), .Z(n27212) );
  ANDN U33855 ( .B(n27707), .A(n27708), .Z(n27705) );
  AND U33856 ( .A(a[58]), .B(b[25]), .Z(n27704) );
  XOR U33857 ( .A(n27710), .B(n27711), .Z(n27217) );
  ANDN U33858 ( .B(n27712), .A(n27713), .Z(n27710) );
  AND U33859 ( .A(a[59]), .B(b[24]), .Z(n27709) );
  XOR U33860 ( .A(n27715), .B(n27716), .Z(n27222) );
  ANDN U33861 ( .B(n27717), .A(n27718), .Z(n27715) );
  AND U33862 ( .A(a[60]), .B(b[23]), .Z(n27714) );
  XOR U33863 ( .A(n27720), .B(n27721), .Z(n27227) );
  ANDN U33864 ( .B(n27722), .A(n27723), .Z(n27720) );
  AND U33865 ( .A(a[61]), .B(b[22]), .Z(n27719) );
  XOR U33866 ( .A(n27725), .B(n27726), .Z(n27232) );
  ANDN U33867 ( .B(n27727), .A(n27728), .Z(n27725) );
  AND U33868 ( .A(a[62]), .B(b[21]), .Z(n27724) );
  XOR U33869 ( .A(n27730), .B(n27731), .Z(n27237) );
  ANDN U33870 ( .B(n27732), .A(n27733), .Z(n27730) );
  AND U33871 ( .A(a[63]), .B(b[20]), .Z(n27729) );
  XOR U33872 ( .A(n27735), .B(n27736), .Z(n27242) );
  ANDN U33873 ( .B(n27737), .A(n27738), .Z(n27735) );
  AND U33874 ( .A(a[64]), .B(b[19]), .Z(n27734) );
  XOR U33875 ( .A(n27740), .B(n27741), .Z(n27247) );
  ANDN U33876 ( .B(n27742), .A(n27743), .Z(n27740) );
  AND U33877 ( .A(a[65]), .B(b[18]), .Z(n27739) );
  XOR U33878 ( .A(n27745), .B(n27746), .Z(n27252) );
  ANDN U33879 ( .B(n27747), .A(n27748), .Z(n27745) );
  AND U33880 ( .A(a[66]), .B(b[17]), .Z(n27744) );
  XOR U33881 ( .A(n27750), .B(n27751), .Z(n27257) );
  ANDN U33882 ( .B(n27752), .A(n27753), .Z(n27750) );
  AND U33883 ( .A(a[67]), .B(b[16]), .Z(n27749) );
  XOR U33884 ( .A(n27755), .B(n27756), .Z(n27262) );
  ANDN U33885 ( .B(n27757), .A(n27758), .Z(n27755) );
  AND U33886 ( .A(a[68]), .B(b[15]), .Z(n27754) );
  XOR U33887 ( .A(n27760), .B(n27761), .Z(n27267) );
  ANDN U33888 ( .B(n27762), .A(n27763), .Z(n27760) );
  AND U33889 ( .A(a[69]), .B(b[14]), .Z(n27759) );
  XOR U33890 ( .A(n27765), .B(n27766), .Z(n27272) );
  ANDN U33891 ( .B(n27767), .A(n27768), .Z(n27765) );
  AND U33892 ( .A(a[70]), .B(b[13]), .Z(n27764) );
  XOR U33893 ( .A(n27770), .B(n27771), .Z(n27277) );
  ANDN U33894 ( .B(n27772), .A(n27773), .Z(n27770) );
  AND U33895 ( .A(a[71]), .B(b[12]), .Z(n27769) );
  XOR U33896 ( .A(n27775), .B(n27776), .Z(n27282) );
  ANDN U33897 ( .B(n27777), .A(n27778), .Z(n27775) );
  AND U33898 ( .A(a[72]), .B(b[11]), .Z(n27774) );
  XOR U33899 ( .A(n27780), .B(n27781), .Z(n27287) );
  ANDN U33900 ( .B(n27782), .A(n27783), .Z(n27780) );
  AND U33901 ( .A(a[73]), .B(b[10]), .Z(n27779) );
  XOR U33902 ( .A(n27785), .B(n27786), .Z(n27292) );
  ANDN U33903 ( .B(n27787), .A(n27788), .Z(n27785) );
  AND U33904 ( .A(b[9]), .B(a[74]), .Z(n27784) );
  XOR U33905 ( .A(n27790), .B(n27791), .Z(n27297) );
  ANDN U33906 ( .B(n27792), .A(n27793), .Z(n27790) );
  AND U33907 ( .A(b[8]), .B(a[75]), .Z(n27789) );
  XOR U33908 ( .A(n27795), .B(n27796), .Z(n27302) );
  ANDN U33909 ( .B(n27797), .A(n27798), .Z(n27795) );
  AND U33910 ( .A(b[7]), .B(a[76]), .Z(n27794) );
  XOR U33911 ( .A(n27800), .B(n27801), .Z(n27307) );
  ANDN U33912 ( .B(n27802), .A(n27803), .Z(n27800) );
  AND U33913 ( .A(b[6]), .B(a[77]), .Z(n27799) );
  XOR U33914 ( .A(n27805), .B(n27806), .Z(n27312) );
  ANDN U33915 ( .B(n27807), .A(n27808), .Z(n27805) );
  AND U33916 ( .A(b[5]), .B(a[78]), .Z(n27804) );
  XOR U33917 ( .A(n27810), .B(n27811), .Z(n27317) );
  ANDN U33918 ( .B(n27812), .A(n27813), .Z(n27810) );
  AND U33919 ( .A(b[4]), .B(a[79]), .Z(n27809) );
  XOR U33920 ( .A(n27815), .B(n27816), .Z(n27322) );
  ANDN U33921 ( .B(n27334), .A(n27335), .Z(n27815) );
  AND U33922 ( .A(b[2]), .B(a[80]), .Z(n27817) );
  XNOR U33923 ( .A(n27812), .B(n27816), .Z(n27818) );
  XOR U33924 ( .A(n27819), .B(n27820), .Z(n27816) );
  OR U33925 ( .A(n27337), .B(n27338), .Z(n27820) );
  XNOR U33926 ( .A(n27822), .B(n27823), .Z(n27821) );
  XOR U33927 ( .A(n27822), .B(n27825), .Z(n27337) );
  NAND U33928 ( .A(b[1]), .B(a[80]), .Z(n27825) );
  IV U33929 ( .A(n27819), .Z(n27822) );
  NANDN U33930 ( .A(n43), .B(n44), .Z(n27819) );
  XOR U33931 ( .A(n27826), .B(n27827), .Z(n44) );
  NAND U33932 ( .A(a[80]), .B(b[0]), .Z(n43) );
  XNOR U33933 ( .A(n27807), .B(n27811), .Z(n27828) );
  XNOR U33934 ( .A(n27802), .B(n27806), .Z(n27829) );
  XNOR U33935 ( .A(n27797), .B(n27801), .Z(n27830) );
  XNOR U33936 ( .A(n27792), .B(n27796), .Z(n27831) );
  XNOR U33937 ( .A(n27787), .B(n27791), .Z(n27832) );
  XNOR U33938 ( .A(n27782), .B(n27786), .Z(n27833) );
  XNOR U33939 ( .A(n27777), .B(n27781), .Z(n27834) );
  XNOR U33940 ( .A(n27772), .B(n27776), .Z(n27835) );
  XNOR U33941 ( .A(n27767), .B(n27771), .Z(n27836) );
  XNOR U33942 ( .A(n27762), .B(n27766), .Z(n27837) );
  XNOR U33943 ( .A(n27757), .B(n27761), .Z(n27838) );
  XNOR U33944 ( .A(n27752), .B(n27756), .Z(n27839) );
  XNOR U33945 ( .A(n27747), .B(n27751), .Z(n27840) );
  XNOR U33946 ( .A(n27742), .B(n27746), .Z(n27841) );
  XNOR U33947 ( .A(n27737), .B(n27741), .Z(n27842) );
  XNOR U33948 ( .A(n27732), .B(n27736), .Z(n27843) );
  XNOR U33949 ( .A(n27727), .B(n27731), .Z(n27844) );
  XNOR U33950 ( .A(n27722), .B(n27726), .Z(n27845) );
  XNOR U33951 ( .A(n27717), .B(n27721), .Z(n27846) );
  XNOR U33952 ( .A(n27712), .B(n27716), .Z(n27847) );
  XNOR U33953 ( .A(n27707), .B(n27711), .Z(n27848) );
  XNOR U33954 ( .A(n27702), .B(n27706), .Z(n27849) );
  XNOR U33955 ( .A(n27697), .B(n27701), .Z(n27850) );
  XNOR U33956 ( .A(n27692), .B(n27696), .Z(n27851) );
  XNOR U33957 ( .A(n27687), .B(n27691), .Z(n27852) );
  XNOR U33958 ( .A(n27682), .B(n27686), .Z(n27853) );
  XNOR U33959 ( .A(n27677), .B(n27681), .Z(n27854) );
  XNOR U33960 ( .A(n27672), .B(n27676), .Z(n27855) );
  XNOR U33961 ( .A(n27667), .B(n27671), .Z(n27856) );
  XNOR U33962 ( .A(n27662), .B(n27666), .Z(n27857) );
  XNOR U33963 ( .A(n27657), .B(n27661), .Z(n27858) );
  XNOR U33964 ( .A(n27652), .B(n27656), .Z(n27859) );
  XNOR U33965 ( .A(n27647), .B(n27651), .Z(n27860) );
  XNOR U33966 ( .A(n27642), .B(n27646), .Z(n27861) );
  XNOR U33967 ( .A(n27637), .B(n27641), .Z(n27862) );
  XNOR U33968 ( .A(n27632), .B(n27636), .Z(n27863) );
  XNOR U33969 ( .A(n27627), .B(n27631), .Z(n27864) );
  XNOR U33970 ( .A(n27622), .B(n27626), .Z(n27865) );
  XNOR U33971 ( .A(n27617), .B(n27621), .Z(n27866) );
  XNOR U33972 ( .A(n27612), .B(n27616), .Z(n27867) );
  XNOR U33973 ( .A(n27607), .B(n27611), .Z(n27868) );
  XNOR U33974 ( .A(n27602), .B(n27606), .Z(n27869) );
  XNOR U33975 ( .A(n27597), .B(n27601), .Z(n27870) );
  XNOR U33976 ( .A(n27592), .B(n27596), .Z(n27871) );
  XNOR U33977 ( .A(n27587), .B(n27591), .Z(n27872) );
  XNOR U33978 ( .A(n27582), .B(n27586), .Z(n27873) );
  XNOR U33979 ( .A(n27577), .B(n27581), .Z(n27874) );
  XNOR U33980 ( .A(n27572), .B(n27576), .Z(n27875) );
  XNOR U33981 ( .A(n27567), .B(n27571), .Z(n27876) );
  XNOR U33982 ( .A(n27562), .B(n27566), .Z(n27877) );
  XNOR U33983 ( .A(n27557), .B(n27561), .Z(n27878) );
  XNOR U33984 ( .A(n27552), .B(n27556), .Z(n27879) );
  XNOR U33985 ( .A(n27547), .B(n27551), .Z(n27880) );
  XNOR U33986 ( .A(n27542), .B(n27546), .Z(n27881) );
  XNOR U33987 ( .A(n27537), .B(n27541), .Z(n27882) );
  XNOR U33988 ( .A(n27532), .B(n27536), .Z(n27883) );
  XNOR U33989 ( .A(n27527), .B(n27531), .Z(n27884) );
  XNOR U33990 ( .A(n27522), .B(n27526), .Z(n27885) );
  XNOR U33991 ( .A(n27517), .B(n27521), .Z(n27886) );
  XNOR U33992 ( .A(n27512), .B(n27516), .Z(n27887) );
  XNOR U33993 ( .A(n27507), .B(n27511), .Z(n27888) );
  XNOR U33994 ( .A(n27502), .B(n27506), .Z(n27889) );
  XNOR U33995 ( .A(n27497), .B(n27501), .Z(n27890) );
  XNOR U33996 ( .A(n27492), .B(n27496), .Z(n27891) );
  XNOR U33997 ( .A(n27487), .B(n27491), .Z(n27892) );
  XNOR U33998 ( .A(n27482), .B(n27486), .Z(n27893) );
  XNOR U33999 ( .A(n27477), .B(n27481), .Z(n27894) );
  XNOR U34000 ( .A(n27472), .B(n27476), .Z(n27895) );
  XNOR U34001 ( .A(n27467), .B(n27471), .Z(n27896) );
  XNOR U34002 ( .A(n27462), .B(n27466), .Z(n27897) );
  XNOR U34003 ( .A(n27457), .B(n27461), .Z(n27898) );
  XNOR U34004 ( .A(n27452), .B(n27456), .Z(n27899) );
  XNOR U34005 ( .A(n27447), .B(n27451), .Z(n27900) );
  XNOR U34006 ( .A(n27442), .B(n27446), .Z(n27901) );
  XNOR U34007 ( .A(n27437), .B(n27441), .Z(n27902) );
  XNOR U34008 ( .A(n27432), .B(n27436), .Z(n27903) );
  XNOR U34009 ( .A(n27427), .B(n27431), .Z(n27904) );
  XNOR U34010 ( .A(n27422), .B(n27426), .Z(n27905) );
  XOR U34011 ( .A(n27906), .B(n27421), .Z(n27422) );
  AND U34012 ( .A(a[0]), .B(b[82]), .Z(n27906) );
  XNOR U34013 ( .A(n27907), .B(n27421), .Z(n27423) );
  XNOR U34014 ( .A(n27908), .B(n27909), .Z(n27421) );
  ANDN U34015 ( .B(n27910), .A(n27911), .Z(n27908) );
  AND U34016 ( .A(a[1]), .B(b[81]), .Z(n27907) );
  XOR U34017 ( .A(n27913), .B(n27914), .Z(n27426) );
  ANDN U34018 ( .B(n27915), .A(n27916), .Z(n27913) );
  AND U34019 ( .A(a[2]), .B(b[80]), .Z(n27912) );
  XOR U34020 ( .A(n27918), .B(n27919), .Z(n27431) );
  ANDN U34021 ( .B(n27920), .A(n27921), .Z(n27918) );
  AND U34022 ( .A(a[3]), .B(b[79]), .Z(n27917) );
  XOR U34023 ( .A(n27923), .B(n27924), .Z(n27436) );
  ANDN U34024 ( .B(n27925), .A(n27926), .Z(n27923) );
  AND U34025 ( .A(a[4]), .B(b[78]), .Z(n27922) );
  XOR U34026 ( .A(n27928), .B(n27929), .Z(n27441) );
  ANDN U34027 ( .B(n27930), .A(n27931), .Z(n27928) );
  AND U34028 ( .A(a[5]), .B(b[77]), .Z(n27927) );
  XOR U34029 ( .A(n27933), .B(n27934), .Z(n27446) );
  ANDN U34030 ( .B(n27935), .A(n27936), .Z(n27933) );
  AND U34031 ( .A(a[6]), .B(b[76]), .Z(n27932) );
  XOR U34032 ( .A(n27938), .B(n27939), .Z(n27451) );
  ANDN U34033 ( .B(n27940), .A(n27941), .Z(n27938) );
  AND U34034 ( .A(a[7]), .B(b[75]), .Z(n27937) );
  XOR U34035 ( .A(n27943), .B(n27944), .Z(n27456) );
  ANDN U34036 ( .B(n27945), .A(n27946), .Z(n27943) );
  AND U34037 ( .A(a[8]), .B(b[74]), .Z(n27942) );
  XOR U34038 ( .A(n27948), .B(n27949), .Z(n27461) );
  ANDN U34039 ( .B(n27950), .A(n27951), .Z(n27948) );
  AND U34040 ( .A(a[9]), .B(b[73]), .Z(n27947) );
  XOR U34041 ( .A(n27953), .B(n27954), .Z(n27466) );
  ANDN U34042 ( .B(n27955), .A(n27956), .Z(n27953) );
  AND U34043 ( .A(a[10]), .B(b[72]), .Z(n27952) );
  XOR U34044 ( .A(n27958), .B(n27959), .Z(n27471) );
  ANDN U34045 ( .B(n27960), .A(n27961), .Z(n27958) );
  AND U34046 ( .A(a[11]), .B(b[71]), .Z(n27957) );
  XOR U34047 ( .A(n27963), .B(n27964), .Z(n27476) );
  ANDN U34048 ( .B(n27965), .A(n27966), .Z(n27963) );
  AND U34049 ( .A(a[12]), .B(b[70]), .Z(n27962) );
  XOR U34050 ( .A(n27968), .B(n27969), .Z(n27481) );
  ANDN U34051 ( .B(n27970), .A(n27971), .Z(n27968) );
  AND U34052 ( .A(a[13]), .B(b[69]), .Z(n27967) );
  XOR U34053 ( .A(n27973), .B(n27974), .Z(n27486) );
  ANDN U34054 ( .B(n27975), .A(n27976), .Z(n27973) );
  AND U34055 ( .A(a[14]), .B(b[68]), .Z(n27972) );
  XOR U34056 ( .A(n27978), .B(n27979), .Z(n27491) );
  ANDN U34057 ( .B(n27980), .A(n27981), .Z(n27978) );
  AND U34058 ( .A(a[15]), .B(b[67]), .Z(n27977) );
  XOR U34059 ( .A(n27983), .B(n27984), .Z(n27496) );
  ANDN U34060 ( .B(n27985), .A(n27986), .Z(n27983) );
  AND U34061 ( .A(a[16]), .B(b[66]), .Z(n27982) );
  XOR U34062 ( .A(n27988), .B(n27989), .Z(n27501) );
  ANDN U34063 ( .B(n27990), .A(n27991), .Z(n27988) );
  AND U34064 ( .A(a[17]), .B(b[65]), .Z(n27987) );
  XOR U34065 ( .A(n27993), .B(n27994), .Z(n27506) );
  ANDN U34066 ( .B(n27995), .A(n27996), .Z(n27993) );
  AND U34067 ( .A(a[18]), .B(b[64]), .Z(n27992) );
  XOR U34068 ( .A(n27998), .B(n27999), .Z(n27511) );
  ANDN U34069 ( .B(n28000), .A(n28001), .Z(n27998) );
  AND U34070 ( .A(a[19]), .B(b[63]), .Z(n27997) );
  XOR U34071 ( .A(n28003), .B(n28004), .Z(n27516) );
  ANDN U34072 ( .B(n28005), .A(n28006), .Z(n28003) );
  AND U34073 ( .A(a[20]), .B(b[62]), .Z(n28002) );
  XOR U34074 ( .A(n28008), .B(n28009), .Z(n27521) );
  ANDN U34075 ( .B(n28010), .A(n28011), .Z(n28008) );
  AND U34076 ( .A(a[21]), .B(b[61]), .Z(n28007) );
  XOR U34077 ( .A(n28013), .B(n28014), .Z(n27526) );
  ANDN U34078 ( .B(n28015), .A(n28016), .Z(n28013) );
  AND U34079 ( .A(a[22]), .B(b[60]), .Z(n28012) );
  XOR U34080 ( .A(n28018), .B(n28019), .Z(n27531) );
  ANDN U34081 ( .B(n28020), .A(n28021), .Z(n28018) );
  AND U34082 ( .A(a[23]), .B(b[59]), .Z(n28017) );
  XOR U34083 ( .A(n28023), .B(n28024), .Z(n27536) );
  ANDN U34084 ( .B(n28025), .A(n28026), .Z(n28023) );
  AND U34085 ( .A(a[24]), .B(b[58]), .Z(n28022) );
  XOR U34086 ( .A(n28028), .B(n28029), .Z(n27541) );
  ANDN U34087 ( .B(n28030), .A(n28031), .Z(n28028) );
  AND U34088 ( .A(a[25]), .B(b[57]), .Z(n28027) );
  XOR U34089 ( .A(n28033), .B(n28034), .Z(n27546) );
  ANDN U34090 ( .B(n28035), .A(n28036), .Z(n28033) );
  AND U34091 ( .A(a[26]), .B(b[56]), .Z(n28032) );
  XOR U34092 ( .A(n28038), .B(n28039), .Z(n27551) );
  ANDN U34093 ( .B(n28040), .A(n28041), .Z(n28038) );
  AND U34094 ( .A(a[27]), .B(b[55]), .Z(n28037) );
  XOR U34095 ( .A(n28043), .B(n28044), .Z(n27556) );
  ANDN U34096 ( .B(n28045), .A(n28046), .Z(n28043) );
  AND U34097 ( .A(a[28]), .B(b[54]), .Z(n28042) );
  XOR U34098 ( .A(n28048), .B(n28049), .Z(n27561) );
  ANDN U34099 ( .B(n28050), .A(n28051), .Z(n28048) );
  AND U34100 ( .A(a[29]), .B(b[53]), .Z(n28047) );
  XOR U34101 ( .A(n28053), .B(n28054), .Z(n27566) );
  ANDN U34102 ( .B(n28055), .A(n28056), .Z(n28053) );
  AND U34103 ( .A(a[30]), .B(b[52]), .Z(n28052) );
  XOR U34104 ( .A(n28058), .B(n28059), .Z(n27571) );
  ANDN U34105 ( .B(n28060), .A(n28061), .Z(n28058) );
  AND U34106 ( .A(a[31]), .B(b[51]), .Z(n28057) );
  XOR U34107 ( .A(n28063), .B(n28064), .Z(n27576) );
  ANDN U34108 ( .B(n28065), .A(n28066), .Z(n28063) );
  AND U34109 ( .A(a[32]), .B(b[50]), .Z(n28062) );
  XOR U34110 ( .A(n28068), .B(n28069), .Z(n27581) );
  ANDN U34111 ( .B(n28070), .A(n28071), .Z(n28068) );
  AND U34112 ( .A(a[33]), .B(b[49]), .Z(n28067) );
  XOR U34113 ( .A(n28073), .B(n28074), .Z(n27586) );
  ANDN U34114 ( .B(n28075), .A(n28076), .Z(n28073) );
  AND U34115 ( .A(a[34]), .B(b[48]), .Z(n28072) );
  XOR U34116 ( .A(n28078), .B(n28079), .Z(n27591) );
  ANDN U34117 ( .B(n28080), .A(n28081), .Z(n28078) );
  AND U34118 ( .A(a[35]), .B(b[47]), .Z(n28077) );
  XOR U34119 ( .A(n28083), .B(n28084), .Z(n27596) );
  ANDN U34120 ( .B(n28085), .A(n28086), .Z(n28083) );
  AND U34121 ( .A(a[36]), .B(b[46]), .Z(n28082) );
  XOR U34122 ( .A(n28088), .B(n28089), .Z(n27601) );
  ANDN U34123 ( .B(n28090), .A(n28091), .Z(n28088) );
  AND U34124 ( .A(a[37]), .B(b[45]), .Z(n28087) );
  XOR U34125 ( .A(n28093), .B(n28094), .Z(n27606) );
  ANDN U34126 ( .B(n28095), .A(n28096), .Z(n28093) );
  AND U34127 ( .A(a[38]), .B(b[44]), .Z(n28092) );
  XOR U34128 ( .A(n28098), .B(n28099), .Z(n27611) );
  ANDN U34129 ( .B(n28100), .A(n28101), .Z(n28098) );
  AND U34130 ( .A(a[39]), .B(b[43]), .Z(n28097) );
  XOR U34131 ( .A(n28103), .B(n28104), .Z(n27616) );
  ANDN U34132 ( .B(n28105), .A(n28106), .Z(n28103) );
  AND U34133 ( .A(a[40]), .B(b[42]), .Z(n28102) );
  XOR U34134 ( .A(n28108), .B(n28109), .Z(n27621) );
  ANDN U34135 ( .B(n28110), .A(n28111), .Z(n28108) );
  AND U34136 ( .A(a[41]), .B(b[41]), .Z(n28107) );
  XOR U34137 ( .A(n28113), .B(n28114), .Z(n27626) );
  ANDN U34138 ( .B(n28115), .A(n28116), .Z(n28113) );
  AND U34139 ( .A(a[42]), .B(b[40]), .Z(n28112) );
  XOR U34140 ( .A(n28118), .B(n28119), .Z(n27631) );
  ANDN U34141 ( .B(n28120), .A(n28121), .Z(n28118) );
  AND U34142 ( .A(a[43]), .B(b[39]), .Z(n28117) );
  XOR U34143 ( .A(n28123), .B(n28124), .Z(n27636) );
  ANDN U34144 ( .B(n28125), .A(n28126), .Z(n28123) );
  AND U34145 ( .A(a[44]), .B(b[38]), .Z(n28122) );
  XOR U34146 ( .A(n28128), .B(n28129), .Z(n27641) );
  ANDN U34147 ( .B(n28130), .A(n28131), .Z(n28128) );
  AND U34148 ( .A(a[45]), .B(b[37]), .Z(n28127) );
  XOR U34149 ( .A(n28133), .B(n28134), .Z(n27646) );
  ANDN U34150 ( .B(n28135), .A(n28136), .Z(n28133) );
  AND U34151 ( .A(a[46]), .B(b[36]), .Z(n28132) );
  XOR U34152 ( .A(n28138), .B(n28139), .Z(n27651) );
  ANDN U34153 ( .B(n28140), .A(n28141), .Z(n28138) );
  AND U34154 ( .A(a[47]), .B(b[35]), .Z(n28137) );
  XOR U34155 ( .A(n28143), .B(n28144), .Z(n27656) );
  ANDN U34156 ( .B(n28145), .A(n28146), .Z(n28143) );
  AND U34157 ( .A(a[48]), .B(b[34]), .Z(n28142) );
  XOR U34158 ( .A(n28148), .B(n28149), .Z(n27661) );
  ANDN U34159 ( .B(n28150), .A(n28151), .Z(n28148) );
  AND U34160 ( .A(a[49]), .B(b[33]), .Z(n28147) );
  XOR U34161 ( .A(n28153), .B(n28154), .Z(n27666) );
  ANDN U34162 ( .B(n28155), .A(n28156), .Z(n28153) );
  AND U34163 ( .A(a[50]), .B(b[32]), .Z(n28152) );
  XOR U34164 ( .A(n28158), .B(n28159), .Z(n27671) );
  ANDN U34165 ( .B(n28160), .A(n28161), .Z(n28158) );
  AND U34166 ( .A(a[51]), .B(b[31]), .Z(n28157) );
  XOR U34167 ( .A(n28163), .B(n28164), .Z(n27676) );
  ANDN U34168 ( .B(n28165), .A(n28166), .Z(n28163) );
  AND U34169 ( .A(a[52]), .B(b[30]), .Z(n28162) );
  XOR U34170 ( .A(n28168), .B(n28169), .Z(n27681) );
  ANDN U34171 ( .B(n28170), .A(n28171), .Z(n28168) );
  AND U34172 ( .A(a[53]), .B(b[29]), .Z(n28167) );
  XOR U34173 ( .A(n28173), .B(n28174), .Z(n27686) );
  ANDN U34174 ( .B(n28175), .A(n28176), .Z(n28173) );
  AND U34175 ( .A(a[54]), .B(b[28]), .Z(n28172) );
  XOR U34176 ( .A(n28178), .B(n28179), .Z(n27691) );
  ANDN U34177 ( .B(n28180), .A(n28181), .Z(n28178) );
  AND U34178 ( .A(a[55]), .B(b[27]), .Z(n28177) );
  XOR U34179 ( .A(n28183), .B(n28184), .Z(n27696) );
  ANDN U34180 ( .B(n28185), .A(n28186), .Z(n28183) );
  AND U34181 ( .A(a[56]), .B(b[26]), .Z(n28182) );
  XOR U34182 ( .A(n28188), .B(n28189), .Z(n27701) );
  ANDN U34183 ( .B(n28190), .A(n28191), .Z(n28188) );
  AND U34184 ( .A(a[57]), .B(b[25]), .Z(n28187) );
  XOR U34185 ( .A(n28193), .B(n28194), .Z(n27706) );
  ANDN U34186 ( .B(n28195), .A(n28196), .Z(n28193) );
  AND U34187 ( .A(a[58]), .B(b[24]), .Z(n28192) );
  XOR U34188 ( .A(n28198), .B(n28199), .Z(n27711) );
  ANDN U34189 ( .B(n28200), .A(n28201), .Z(n28198) );
  AND U34190 ( .A(a[59]), .B(b[23]), .Z(n28197) );
  XOR U34191 ( .A(n28203), .B(n28204), .Z(n27716) );
  ANDN U34192 ( .B(n28205), .A(n28206), .Z(n28203) );
  AND U34193 ( .A(a[60]), .B(b[22]), .Z(n28202) );
  XOR U34194 ( .A(n28208), .B(n28209), .Z(n27721) );
  ANDN U34195 ( .B(n28210), .A(n28211), .Z(n28208) );
  AND U34196 ( .A(a[61]), .B(b[21]), .Z(n28207) );
  XOR U34197 ( .A(n28213), .B(n28214), .Z(n27726) );
  ANDN U34198 ( .B(n28215), .A(n28216), .Z(n28213) );
  AND U34199 ( .A(a[62]), .B(b[20]), .Z(n28212) );
  XOR U34200 ( .A(n28218), .B(n28219), .Z(n27731) );
  ANDN U34201 ( .B(n28220), .A(n28221), .Z(n28218) );
  AND U34202 ( .A(a[63]), .B(b[19]), .Z(n28217) );
  XOR U34203 ( .A(n28223), .B(n28224), .Z(n27736) );
  ANDN U34204 ( .B(n28225), .A(n28226), .Z(n28223) );
  AND U34205 ( .A(a[64]), .B(b[18]), .Z(n28222) );
  XOR U34206 ( .A(n28228), .B(n28229), .Z(n27741) );
  ANDN U34207 ( .B(n28230), .A(n28231), .Z(n28228) );
  AND U34208 ( .A(a[65]), .B(b[17]), .Z(n28227) );
  XOR U34209 ( .A(n28233), .B(n28234), .Z(n27746) );
  ANDN U34210 ( .B(n28235), .A(n28236), .Z(n28233) );
  AND U34211 ( .A(a[66]), .B(b[16]), .Z(n28232) );
  XOR U34212 ( .A(n28238), .B(n28239), .Z(n27751) );
  ANDN U34213 ( .B(n28240), .A(n28241), .Z(n28238) );
  AND U34214 ( .A(a[67]), .B(b[15]), .Z(n28237) );
  XOR U34215 ( .A(n28243), .B(n28244), .Z(n27756) );
  ANDN U34216 ( .B(n28245), .A(n28246), .Z(n28243) );
  AND U34217 ( .A(a[68]), .B(b[14]), .Z(n28242) );
  XOR U34218 ( .A(n28248), .B(n28249), .Z(n27761) );
  ANDN U34219 ( .B(n28250), .A(n28251), .Z(n28248) );
  AND U34220 ( .A(a[69]), .B(b[13]), .Z(n28247) );
  XOR U34221 ( .A(n28253), .B(n28254), .Z(n27766) );
  ANDN U34222 ( .B(n28255), .A(n28256), .Z(n28253) );
  AND U34223 ( .A(a[70]), .B(b[12]), .Z(n28252) );
  XOR U34224 ( .A(n28258), .B(n28259), .Z(n27771) );
  ANDN U34225 ( .B(n28260), .A(n28261), .Z(n28258) );
  AND U34226 ( .A(a[71]), .B(b[11]), .Z(n28257) );
  XOR U34227 ( .A(n28263), .B(n28264), .Z(n27776) );
  ANDN U34228 ( .B(n28265), .A(n28266), .Z(n28263) );
  AND U34229 ( .A(a[72]), .B(b[10]), .Z(n28262) );
  XOR U34230 ( .A(n28268), .B(n28269), .Z(n27781) );
  ANDN U34231 ( .B(n28270), .A(n28271), .Z(n28268) );
  AND U34232 ( .A(b[9]), .B(a[73]), .Z(n28267) );
  XOR U34233 ( .A(n28273), .B(n28274), .Z(n27786) );
  ANDN U34234 ( .B(n28275), .A(n28276), .Z(n28273) );
  AND U34235 ( .A(b[8]), .B(a[74]), .Z(n28272) );
  XOR U34236 ( .A(n28278), .B(n28279), .Z(n27791) );
  ANDN U34237 ( .B(n28280), .A(n28281), .Z(n28278) );
  AND U34238 ( .A(b[7]), .B(a[75]), .Z(n28277) );
  XOR U34239 ( .A(n28283), .B(n28284), .Z(n27796) );
  ANDN U34240 ( .B(n28285), .A(n28286), .Z(n28283) );
  AND U34241 ( .A(b[6]), .B(a[76]), .Z(n28282) );
  XOR U34242 ( .A(n28288), .B(n28289), .Z(n27801) );
  ANDN U34243 ( .B(n28290), .A(n28291), .Z(n28288) );
  AND U34244 ( .A(b[5]), .B(a[77]), .Z(n28287) );
  XOR U34245 ( .A(n28293), .B(n28294), .Z(n27806) );
  ANDN U34246 ( .B(n28295), .A(n28296), .Z(n28293) );
  AND U34247 ( .A(b[4]), .B(a[78]), .Z(n28292) );
  XOR U34248 ( .A(n28298), .B(n28299), .Z(n27811) );
  ANDN U34249 ( .B(n27823), .A(n27824), .Z(n28298) );
  AND U34250 ( .A(b[2]), .B(a[79]), .Z(n28300) );
  XNOR U34251 ( .A(n28295), .B(n28299), .Z(n28301) );
  XOR U34252 ( .A(n28302), .B(n28303), .Z(n28299) );
  OR U34253 ( .A(n27826), .B(n27827), .Z(n28303) );
  XNOR U34254 ( .A(n28305), .B(n28306), .Z(n28304) );
  XOR U34255 ( .A(n28305), .B(n28308), .Z(n27826) );
  NAND U34256 ( .A(b[1]), .B(a[79]), .Z(n28308) );
  IV U34257 ( .A(n28302), .Z(n28305) );
  NANDN U34258 ( .A(n47), .B(n48), .Z(n28302) );
  XOR U34259 ( .A(n28309), .B(n28310), .Z(n48) );
  NAND U34260 ( .A(a[79]), .B(b[0]), .Z(n47) );
  XNOR U34261 ( .A(n28290), .B(n28294), .Z(n28311) );
  XNOR U34262 ( .A(n28285), .B(n28289), .Z(n28312) );
  XNOR U34263 ( .A(n28280), .B(n28284), .Z(n28313) );
  XNOR U34264 ( .A(n28275), .B(n28279), .Z(n28314) );
  XNOR U34265 ( .A(n28270), .B(n28274), .Z(n28315) );
  XNOR U34266 ( .A(n28265), .B(n28269), .Z(n28316) );
  XNOR U34267 ( .A(n28260), .B(n28264), .Z(n28317) );
  XNOR U34268 ( .A(n28255), .B(n28259), .Z(n28318) );
  XNOR U34269 ( .A(n28250), .B(n28254), .Z(n28319) );
  XNOR U34270 ( .A(n28245), .B(n28249), .Z(n28320) );
  XNOR U34271 ( .A(n28240), .B(n28244), .Z(n28321) );
  XNOR U34272 ( .A(n28235), .B(n28239), .Z(n28322) );
  XNOR U34273 ( .A(n28230), .B(n28234), .Z(n28323) );
  XNOR U34274 ( .A(n28225), .B(n28229), .Z(n28324) );
  XNOR U34275 ( .A(n28220), .B(n28224), .Z(n28325) );
  XNOR U34276 ( .A(n28215), .B(n28219), .Z(n28326) );
  XNOR U34277 ( .A(n28210), .B(n28214), .Z(n28327) );
  XNOR U34278 ( .A(n28205), .B(n28209), .Z(n28328) );
  XNOR U34279 ( .A(n28200), .B(n28204), .Z(n28329) );
  XNOR U34280 ( .A(n28195), .B(n28199), .Z(n28330) );
  XNOR U34281 ( .A(n28190), .B(n28194), .Z(n28331) );
  XNOR U34282 ( .A(n28185), .B(n28189), .Z(n28332) );
  XNOR U34283 ( .A(n28180), .B(n28184), .Z(n28333) );
  XNOR U34284 ( .A(n28175), .B(n28179), .Z(n28334) );
  XNOR U34285 ( .A(n28170), .B(n28174), .Z(n28335) );
  XNOR U34286 ( .A(n28165), .B(n28169), .Z(n28336) );
  XNOR U34287 ( .A(n28160), .B(n28164), .Z(n28337) );
  XNOR U34288 ( .A(n28155), .B(n28159), .Z(n28338) );
  XNOR U34289 ( .A(n28150), .B(n28154), .Z(n28339) );
  XNOR U34290 ( .A(n28145), .B(n28149), .Z(n28340) );
  XNOR U34291 ( .A(n28140), .B(n28144), .Z(n28341) );
  XNOR U34292 ( .A(n28135), .B(n28139), .Z(n28342) );
  XNOR U34293 ( .A(n28130), .B(n28134), .Z(n28343) );
  XNOR U34294 ( .A(n28125), .B(n28129), .Z(n28344) );
  XNOR U34295 ( .A(n28120), .B(n28124), .Z(n28345) );
  XNOR U34296 ( .A(n28115), .B(n28119), .Z(n28346) );
  XNOR U34297 ( .A(n28110), .B(n28114), .Z(n28347) );
  XNOR U34298 ( .A(n28105), .B(n28109), .Z(n28348) );
  XNOR U34299 ( .A(n28100), .B(n28104), .Z(n28349) );
  XNOR U34300 ( .A(n28095), .B(n28099), .Z(n28350) );
  XNOR U34301 ( .A(n28090), .B(n28094), .Z(n28351) );
  XNOR U34302 ( .A(n28085), .B(n28089), .Z(n28352) );
  XNOR U34303 ( .A(n28080), .B(n28084), .Z(n28353) );
  XNOR U34304 ( .A(n28075), .B(n28079), .Z(n28354) );
  XNOR U34305 ( .A(n28070), .B(n28074), .Z(n28355) );
  XNOR U34306 ( .A(n28065), .B(n28069), .Z(n28356) );
  XNOR U34307 ( .A(n28060), .B(n28064), .Z(n28357) );
  XNOR U34308 ( .A(n28055), .B(n28059), .Z(n28358) );
  XNOR U34309 ( .A(n28050), .B(n28054), .Z(n28359) );
  XNOR U34310 ( .A(n28045), .B(n28049), .Z(n28360) );
  XNOR U34311 ( .A(n28040), .B(n28044), .Z(n28361) );
  XNOR U34312 ( .A(n28035), .B(n28039), .Z(n28362) );
  XNOR U34313 ( .A(n28030), .B(n28034), .Z(n28363) );
  XNOR U34314 ( .A(n28025), .B(n28029), .Z(n28364) );
  XNOR U34315 ( .A(n28020), .B(n28024), .Z(n28365) );
  XNOR U34316 ( .A(n28015), .B(n28019), .Z(n28366) );
  XNOR U34317 ( .A(n28010), .B(n28014), .Z(n28367) );
  XNOR U34318 ( .A(n28005), .B(n28009), .Z(n28368) );
  XNOR U34319 ( .A(n28000), .B(n28004), .Z(n28369) );
  XNOR U34320 ( .A(n27995), .B(n27999), .Z(n28370) );
  XNOR U34321 ( .A(n27990), .B(n27994), .Z(n28371) );
  XNOR U34322 ( .A(n27985), .B(n27989), .Z(n28372) );
  XNOR U34323 ( .A(n27980), .B(n27984), .Z(n28373) );
  XNOR U34324 ( .A(n27975), .B(n27979), .Z(n28374) );
  XNOR U34325 ( .A(n27970), .B(n27974), .Z(n28375) );
  XNOR U34326 ( .A(n27965), .B(n27969), .Z(n28376) );
  XNOR U34327 ( .A(n27960), .B(n27964), .Z(n28377) );
  XNOR U34328 ( .A(n27955), .B(n27959), .Z(n28378) );
  XNOR U34329 ( .A(n27950), .B(n27954), .Z(n28379) );
  XNOR U34330 ( .A(n27945), .B(n27949), .Z(n28380) );
  XNOR U34331 ( .A(n27940), .B(n27944), .Z(n28381) );
  XNOR U34332 ( .A(n27935), .B(n27939), .Z(n28382) );
  XNOR U34333 ( .A(n27930), .B(n27934), .Z(n28383) );
  XNOR U34334 ( .A(n27925), .B(n27929), .Z(n28384) );
  XNOR U34335 ( .A(n27920), .B(n27924), .Z(n28385) );
  XNOR U34336 ( .A(n27915), .B(n27919), .Z(n28386) );
  XNOR U34337 ( .A(n27910), .B(n27914), .Z(n28387) );
  XNOR U34338 ( .A(n28388), .B(n27909), .Z(n27910) );
  AND U34339 ( .A(a[0]), .B(b[81]), .Z(n28388) );
  XOR U34340 ( .A(n28389), .B(n27909), .Z(n27911) );
  XNOR U34341 ( .A(n28390), .B(n28391), .Z(n27909) );
  ANDN U34342 ( .B(n28392), .A(n28393), .Z(n28390) );
  AND U34343 ( .A(a[1]), .B(b[80]), .Z(n28389) );
  XOR U34344 ( .A(n28395), .B(n28396), .Z(n27914) );
  ANDN U34345 ( .B(n28397), .A(n28398), .Z(n28395) );
  AND U34346 ( .A(a[2]), .B(b[79]), .Z(n28394) );
  XOR U34347 ( .A(n28400), .B(n28401), .Z(n27919) );
  ANDN U34348 ( .B(n28402), .A(n28403), .Z(n28400) );
  AND U34349 ( .A(a[3]), .B(b[78]), .Z(n28399) );
  XOR U34350 ( .A(n28405), .B(n28406), .Z(n27924) );
  ANDN U34351 ( .B(n28407), .A(n28408), .Z(n28405) );
  AND U34352 ( .A(a[4]), .B(b[77]), .Z(n28404) );
  XOR U34353 ( .A(n28410), .B(n28411), .Z(n27929) );
  ANDN U34354 ( .B(n28412), .A(n28413), .Z(n28410) );
  AND U34355 ( .A(a[5]), .B(b[76]), .Z(n28409) );
  XOR U34356 ( .A(n28415), .B(n28416), .Z(n27934) );
  ANDN U34357 ( .B(n28417), .A(n28418), .Z(n28415) );
  AND U34358 ( .A(a[6]), .B(b[75]), .Z(n28414) );
  XOR U34359 ( .A(n28420), .B(n28421), .Z(n27939) );
  ANDN U34360 ( .B(n28422), .A(n28423), .Z(n28420) );
  AND U34361 ( .A(a[7]), .B(b[74]), .Z(n28419) );
  XOR U34362 ( .A(n28425), .B(n28426), .Z(n27944) );
  ANDN U34363 ( .B(n28427), .A(n28428), .Z(n28425) );
  AND U34364 ( .A(a[8]), .B(b[73]), .Z(n28424) );
  XOR U34365 ( .A(n28430), .B(n28431), .Z(n27949) );
  ANDN U34366 ( .B(n28432), .A(n28433), .Z(n28430) );
  AND U34367 ( .A(a[9]), .B(b[72]), .Z(n28429) );
  XOR U34368 ( .A(n28435), .B(n28436), .Z(n27954) );
  ANDN U34369 ( .B(n28437), .A(n28438), .Z(n28435) );
  AND U34370 ( .A(a[10]), .B(b[71]), .Z(n28434) );
  XOR U34371 ( .A(n28440), .B(n28441), .Z(n27959) );
  ANDN U34372 ( .B(n28442), .A(n28443), .Z(n28440) );
  AND U34373 ( .A(a[11]), .B(b[70]), .Z(n28439) );
  XOR U34374 ( .A(n28445), .B(n28446), .Z(n27964) );
  ANDN U34375 ( .B(n28447), .A(n28448), .Z(n28445) );
  AND U34376 ( .A(a[12]), .B(b[69]), .Z(n28444) );
  XOR U34377 ( .A(n28450), .B(n28451), .Z(n27969) );
  ANDN U34378 ( .B(n28452), .A(n28453), .Z(n28450) );
  AND U34379 ( .A(a[13]), .B(b[68]), .Z(n28449) );
  XOR U34380 ( .A(n28455), .B(n28456), .Z(n27974) );
  ANDN U34381 ( .B(n28457), .A(n28458), .Z(n28455) );
  AND U34382 ( .A(a[14]), .B(b[67]), .Z(n28454) );
  XOR U34383 ( .A(n28460), .B(n28461), .Z(n27979) );
  ANDN U34384 ( .B(n28462), .A(n28463), .Z(n28460) );
  AND U34385 ( .A(a[15]), .B(b[66]), .Z(n28459) );
  XOR U34386 ( .A(n28465), .B(n28466), .Z(n27984) );
  ANDN U34387 ( .B(n28467), .A(n28468), .Z(n28465) );
  AND U34388 ( .A(a[16]), .B(b[65]), .Z(n28464) );
  XOR U34389 ( .A(n28470), .B(n28471), .Z(n27989) );
  ANDN U34390 ( .B(n28472), .A(n28473), .Z(n28470) );
  AND U34391 ( .A(a[17]), .B(b[64]), .Z(n28469) );
  XOR U34392 ( .A(n28475), .B(n28476), .Z(n27994) );
  ANDN U34393 ( .B(n28477), .A(n28478), .Z(n28475) );
  AND U34394 ( .A(a[18]), .B(b[63]), .Z(n28474) );
  XOR U34395 ( .A(n28480), .B(n28481), .Z(n27999) );
  ANDN U34396 ( .B(n28482), .A(n28483), .Z(n28480) );
  AND U34397 ( .A(a[19]), .B(b[62]), .Z(n28479) );
  XOR U34398 ( .A(n28485), .B(n28486), .Z(n28004) );
  ANDN U34399 ( .B(n28487), .A(n28488), .Z(n28485) );
  AND U34400 ( .A(a[20]), .B(b[61]), .Z(n28484) );
  XOR U34401 ( .A(n28490), .B(n28491), .Z(n28009) );
  ANDN U34402 ( .B(n28492), .A(n28493), .Z(n28490) );
  AND U34403 ( .A(a[21]), .B(b[60]), .Z(n28489) );
  XOR U34404 ( .A(n28495), .B(n28496), .Z(n28014) );
  ANDN U34405 ( .B(n28497), .A(n28498), .Z(n28495) );
  AND U34406 ( .A(a[22]), .B(b[59]), .Z(n28494) );
  XOR U34407 ( .A(n28500), .B(n28501), .Z(n28019) );
  ANDN U34408 ( .B(n28502), .A(n28503), .Z(n28500) );
  AND U34409 ( .A(a[23]), .B(b[58]), .Z(n28499) );
  XOR U34410 ( .A(n28505), .B(n28506), .Z(n28024) );
  ANDN U34411 ( .B(n28507), .A(n28508), .Z(n28505) );
  AND U34412 ( .A(a[24]), .B(b[57]), .Z(n28504) );
  XOR U34413 ( .A(n28510), .B(n28511), .Z(n28029) );
  ANDN U34414 ( .B(n28512), .A(n28513), .Z(n28510) );
  AND U34415 ( .A(a[25]), .B(b[56]), .Z(n28509) );
  XOR U34416 ( .A(n28515), .B(n28516), .Z(n28034) );
  ANDN U34417 ( .B(n28517), .A(n28518), .Z(n28515) );
  AND U34418 ( .A(a[26]), .B(b[55]), .Z(n28514) );
  XOR U34419 ( .A(n28520), .B(n28521), .Z(n28039) );
  ANDN U34420 ( .B(n28522), .A(n28523), .Z(n28520) );
  AND U34421 ( .A(a[27]), .B(b[54]), .Z(n28519) );
  XOR U34422 ( .A(n28525), .B(n28526), .Z(n28044) );
  ANDN U34423 ( .B(n28527), .A(n28528), .Z(n28525) );
  AND U34424 ( .A(a[28]), .B(b[53]), .Z(n28524) );
  XOR U34425 ( .A(n28530), .B(n28531), .Z(n28049) );
  ANDN U34426 ( .B(n28532), .A(n28533), .Z(n28530) );
  AND U34427 ( .A(a[29]), .B(b[52]), .Z(n28529) );
  XOR U34428 ( .A(n28535), .B(n28536), .Z(n28054) );
  ANDN U34429 ( .B(n28537), .A(n28538), .Z(n28535) );
  AND U34430 ( .A(a[30]), .B(b[51]), .Z(n28534) );
  XOR U34431 ( .A(n28540), .B(n28541), .Z(n28059) );
  ANDN U34432 ( .B(n28542), .A(n28543), .Z(n28540) );
  AND U34433 ( .A(a[31]), .B(b[50]), .Z(n28539) );
  XOR U34434 ( .A(n28545), .B(n28546), .Z(n28064) );
  ANDN U34435 ( .B(n28547), .A(n28548), .Z(n28545) );
  AND U34436 ( .A(a[32]), .B(b[49]), .Z(n28544) );
  XOR U34437 ( .A(n28550), .B(n28551), .Z(n28069) );
  ANDN U34438 ( .B(n28552), .A(n28553), .Z(n28550) );
  AND U34439 ( .A(a[33]), .B(b[48]), .Z(n28549) );
  XOR U34440 ( .A(n28555), .B(n28556), .Z(n28074) );
  ANDN U34441 ( .B(n28557), .A(n28558), .Z(n28555) );
  AND U34442 ( .A(a[34]), .B(b[47]), .Z(n28554) );
  XOR U34443 ( .A(n28560), .B(n28561), .Z(n28079) );
  ANDN U34444 ( .B(n28562), .A(n28563), .Z(n28560) );
  AND U34445 ( .A(a[35]), .B(b[46]), .Z(n28559) );
  XOR U34446 ( .A(n28565), .B(n28566), .Z(n28084) );
  ANDN U34447 ( .B(n28567), .A(n28568), .Z(n28565) );
  AND U34448 ( .A(a[36]), .B(b[45]), .Z(n28564) );
  XOR U34449 ( .A(n28570), .B(n28571), .Z(n28089) );
  ANDN U34450 ( .B(n28572), .A(n28573), .Z(n28570) );
  AND U34451 ( .A(a[37]), .B(b[44]), .Z(n28569) );
  XOR U34452 ( .A(n28575), .B(n28576), .Z(n28094) );
  ANDN U34453 ( .B(n28577), .A(n28578), .Z(n28575) );
  AND U34454 ( .A(a[38]), .B(b[43]), .Z(n28574) );
  XOR U34455 ( .A(n28580), .B(n28581), .Z(n28099) );
  ANDN U34456 ( .B(n28582), .A(n28583), .Z(n28580) );
  AND U34457 ( .A(a[39]), .B(b[42]), .Z(n28579) );
  XOR U34458 ( .A(n28585), .B(n28586), .Z(n28104) );
  ANDN U34459 ( .B(n28587), .A(n28588), .Z(n28585) );
  AND U34460 ( .A(a[40]), .B(b[41]), .Z(n28584) );
  XOR U34461 ( .A(n28590), .B(n28591), .Z(n28109) );
  ANDN U34462 ( .B(n28592), .A(n28593), .Z(n28590) );
  AND U34463 ( .A(a[41]), .B(b[40]), .Z(n28589) );
  XOR U34464 ( .A(n28595), .B(n28596), .Z(n28114) );
  ANDN U34465 ( .B(n28597), .A(n28598), .Z(n28595) );
  AND U34466 ( .A(a[42]), .B(b[39]), .Z(n28594) );
  XOR U34467 ( .A(n28600), .B(n28601), .Z(n28119) );
  ANDN U34468 ( .B(n28602), .A(n28603), .Z(n28600) );
  AND U34469 ( .A(a[43]), .B(b[38]), .Z(n28599) );
  XOR U34470 ( .A(n28605), .B(n28606), .Z(n28124) );
  ANDN U34471 ( .B(n28607), .A(n28608), .Z(n28605) );
  AND U34472 ( .A(a[44]), .B(b[37]), .Z(n28604) );
  XOR U34473 ( .A(n28610), .B(n28611), .Z(n28129) );
  ANDN U34474 ( .B(n28612), .A(n28613), .Z(n28610) );
  AND U34475 ( .A(a[45]), .B(b[36]), .Z(n28609) );
  XOR U34476 ( .A(n28615), .B(n28616), .Z(n28134) );
  ANDN U34477 ( .B(n28617), .A(n28618), .Z(n28615) );
  AND U34478 ( .A(a[46]), .B(b[35]), .Z(n28614) );
  XOR U34479 ( .A(n28620), .B(n28621), .Z(n28139) );
  ANDN U34480 ( .B(n28622), .A(n28623), .Z(n28620) );
  AND U34481 ( .A(a[47]), .B(b[34]), .Z(n28619) );
  XOR U34482 ( .A(n28625), .B(n28626), .Z(n28144) );
  ANDN U34483 ( .B(n28627), .A(n28628), .Z(n28625) );
  AND U34484 ( .A(a[48]), .B(b[33]), .Z(n28624) );
  XOR U34485 ( .A(n28630), .B(n28631), .Z(n28149) );
  ANDN U34486 ( .B(n28632), .A(n28633), .Z(n28630) );
  AND U34487 ( .A(a[49]), .B(b[32]), .Z(n28629) );
  XOR U34488 ( .A(n28635), .B(n28636), .Z(n28154) );
  ANDN U34489 ( .B(n28637), .A(n28638), .Z(n28635) );
  AND U34490 ( .A(a[50]), .B(b[31]), .Z(n28634) );
  XOR U34491 ( .A(n28640), .B(n28641), .Z(n28159) );
  ANDN U34492 ( .B(n28642), .A(n28643), .Z(n28640) );
  AND U34493 ( .A(a[51]), .B(b[30]), .Z(n28639) );
  XOR U34494 ( .A(n28645), .B(n28646), .Z(n28164) );
  ANDN U34495 ( .B(n28647), .A(n28648), .Z(n28645) );
  AND U34496 ( .A(a[52]), .B(b[29]), .Z(n28644) );
  XOR U34497 ( .A(n28650), .B(n28651), .Z(n28169) );
  ANDN U34498 ( .B(n28652), .A(n28653), .Z(n28650) );
  AND U34499 ( .A(a[53]), .B(b[28]), .Z(n28649) );
  XOR U34500 ( .A(n28655), .B(n28656), .Z(n28174) );
  ANDN U34501 ( .B(n28657), .A(n28658), .Z(n28655) );
  AND U34502 ( .A(a[54]), .B(b[27]), .Z(n28654) );
  XOR U34503 ( .A(n28660), .B(n28661), .Z(n28179) );
  ANDN U34504 ( .B(n28662), .A(n28663), .Z(n28660) );
  AND U34505 ( .A(a[55]), .B(b[26]), .Z(n28659) );
  XOR U34506 ( .A(n28665), .B(n28666), .Z(n28184) );
  ANDN U34507 ( .B(n28667), .A(n28668), .Z(n28665) );
  AND U34508 ( .A(a[56]), .B(b[25]), .Z(n28664) );
  XOR U34509 ( .A(n28670), .B(n28671), .Z(n28189) );
  ANDN U34510 ( .B(n28672), .A(n28673), .Z(n28670) );
  AND U34511 ( .A(a[57]), .B(b[24]), .Z(n28669) );
  XOR U34512 ( .A(n28675), .B(n28676), .Z(n28194) );
  ANDN U34513 ( .B(n28677), .A(n28678), .Z(n28675) );
  AND U34514 ( .A(a[58]), .B(b[23]), .Z(n28674) );
  XOR U34515 ( .A(n28680), .B(n28681), .Z(n28199) );
  ANDN U34516 ( .B(n28682), .A(n28683), .Z(n28680) );
  AND U34517 ( .A(a[59]), .B(b[22]), .Z(n28679) );
  XOR U34518 ( .A(n28685), .B(n28686), .Z(n28204) );
  ANDN U34519 ( .B(n28687), .A(n28688), .Z(n28685) );
  AND U34520 ( .A(a[60]), .B(b[21]), .Z(n28684) );
  XOR U34521 ( .A(n28690), .B(n28691), .Z(n28209) );
  ANDN U34522 ( .B(n28692), .A(n28693), .Z(n28690) );
  AND U34523 ( .A(a[61]), .B(b[20]), .Z(n28689) );
  XOR U34524 ( .A(n28695), .B(n28696), .Z(n28214) );
  ANDN U34525 ( .B(n28697), .A(n28698), .Z(n28695) );
  AND U34526 ( .A(a[62]), .B(b[19]), .Z(n28694) );
  XOR U34527 ( .A(n28700), .B(n28701), .Z(n28219) );
  ANDN U34528 ( .B(n28702), .A(n28703), .Z(n28700) );
  AND U34529 ( .A(a[63]), .B(b[18]), .Z(n28699) );
  XOR U34530 ( .A(n28705), .B(n28706), .Z(n28224) );
  ANDN U34531 ( .B(n28707), .A(n28708), .Z(n28705) );
  AND U34532 ( .A(a[64]), .B(b[17]), .Z(n28704) );
  XOR U34533 ( .A(n28710), .B(n28711), .Z(n28229) );
  ANDN U34534 ( .B(n28712), .A(n28713), .Z(n28710) );
  AND U34535 ( .A(a[65]), .B(b[16]), .Z(n28709) );
  XOR U34536 ( .A(n28715), .B(n28716), .Z(n28234) );
  ANDN U34537 ( .B(n28717), .A(n28718), .Z(n28715) );
  AND U34538 ( .A(a[66]), .B(b[15]), .Z(n28714) );
  XOR U34539 ( .A(n28720), .B(n28721), .Z(n28239) );
  ANDN U34540 ( .B(n28722), .A(n28723), .Z(n28720) );
  AND U34541 ( .A(a[67]), .B(b[14]), .Z(n28719) );
  XOR U34542 ( .A(n28725), .B(n28726), .Z(n28244) );
  ANDN U34543 ( .B(n28727), .A(n28728), .Z(n28725) );
  AND U34544 ( .A(a[68]), .B(b[13]), .Z(n28724) );
  XOR U34545 ( .A(n28730), .B(n28731), .Z(n28249) );
  ANDN U34546 ( .B(n28732), .A(n28733), .Z(n28730) );
  AND U34547 ( .A(a[69]), .B(b[12]), .Z(n28729) );
  XOR U34548 ( .A(n28735), .B(n28736), .Z(n28254) );
  ANDN U34549 ( .B(n28737), .A(n28738), .Z(n28735) );
  AND U34550 ( .A(a[70]), .B(b[11]), .Z(n28734) );
  XOR U34551 ( .A(n28740), .B(n28741), .Z(n28259) );
  ANDN U34552 ( .B(n28742), .A(n28743), .Z(n28740) );
  AND U34553 ( .A(a[71]), .B(b[10]), .Z(n28739) );
  XOR U34554 ( .A(n28745), .B(n28746), .Z(n28264) );
  ANDN U34555 ( .B(n28747), .A(n28748), .Z(n28745) );
  AND U34556 ( .A(b[9]), .B(a[72]), .Z(n28744) );
  XOR U34557 ( .A(n28750), .B(n28751), .Z(n28269) );
  ANDN U34558 ( .B(n28752), .A(n28753), .Z(n28750) );
  AND U34559 ( .A(b[8]), .B(a[73]), .Z(n28749) );
  XOR U34560 ( .A(n28755), .B(n28756), .Z(n28274) );
  ANDN U34561 ( .B(n28757), .A(n28758), .Z(n28755) );
  AND U34562 ( .A(b[7]), .B(a[74]), .Z(n28754) );
  XOR U34563 ( .A(n28760), .B(n28761), .Z(n28279) );
  ANDN U34564 ( .B(n28762), .A(n28763), .Z(n28760) );
  AND U34565 ( .A(b[6]), .B(a[75]), .Z(n28759) );
  XOR U34566 ( .A(n28765), .B(n28766), .Z(n28284) );
  ANDN U34567 ( .B(n28767), .A(n28768), .Z(n28765) );
  AND U34568 ( .A(b[5]), .B(a[76]), .Z(n28764) );
  XOR U34569 ( .A(n28770), .B(n28771), .Z(n28289) );
  ANDN U34570 ( .B(n28772), .A(n28773), .Z(n28770) );
  AND U34571 ( .A(b[4]), .B(a[77]), .Z(n28769) );
  XOR U34572 ( .A(n28775), .B(n28776), .Z(n28294) );
  ANDN U34573 ( .B(n28306), .A(n28307), .Z(n28775) );
  AND U34574 ( .A(b[2]), .B(a[78]), .Z(n28777) );
  XNOR U34575 ( .A(n28772), .B(n28776), .Z(n28778) );
  XOR U34576 ( .A(n28779), .B(n28780), .Z(n28776) );
  OR U34577 ( .A(n28309), .B(n28310), .Z(n28780) );
  XNOR U34578 ( .A(n28782), .B(n28783), .Z(n28781) );
  XOR U34579 ( .A(n28782), .B(n28785), .Z(n28309) );
  NAND U34580 ( .A(b[1]), .B(a[78]), .Z(n28785) );
  IV U34581 ( .A(n28779), .Z(n28782) );
  NANDN U34582 ( .A(n49), .B(n50), .Z(n28779) );
  XOR U34583 ( .A(n28786), .B(n28787), .Z(n50) );
  NAND U34584 ( .A(a[78]), .B(b[0]), .Z(n49) );
  XNOR U34585 ( .A(n28767), .B(n28771), .Z(n28788) );
  XNOR U34586 ( .A(n28762), .B(n28766), .Z(n28789) );
  XNOR U34587 ( .A(n28757), .B(n28761), .Z(n28790) );
  XNOR U34588 ( .A(n28752), .B(n28756), .Z(n28791) );
  XNOR U34589 ( .A(n28747), .B(n28751), .Z(n28792) );
  XNOR U34590 ( .A(n28742), .B(n28746), .Z(n28793) );
  XNOR U34591 ( .A(n28737), .B(n28741), .Z(n28794) );
  XNOR U34592 ( .A(n28732), .B(n28736), .Z(n28795) );
  XNOR U34593 ( .A(n28727), .B(n28731), .Z(n28796) );
  XNOR U34594 ( .A(n28722), .B(n28726), .Z(n28797) );
  XNOR U34595 ( .A(n28717), .B(n28721), .Z(n28798) );
  XNOR U34596 ( .A(n28712), .B(n28716), .Z(n28799) );
  XNOR U34597 ( .A(n28707), .B(n28711), .Z(n28800) );
  XNOR U34598 ( .A(n28702), .B(n28706), .Z(n28801) );
  XNOR U34599 ( .A(n28697), .B(n28701), .Z(n28802) );
  XNOR U34600 ( .A(n28692), .B(n28696), .Z(n28803) );
  XNOR U34601 ( .A(n28687), .B(n28691), .Z(n28804) );
  XNOR U34602 ( .A(n28682), .B(n28686), .Z(n28805) );
  XNOR U34603 ( .A(n28677), .B(n28681), .Z(n28806) );
  XNOR U34604 ( .A(n28672), .B(n28676), .Z(n28807) );
  XNOR U34605 ( .A(n28667), .B(n28671), .Z(n28808) );
  XNOR U34606 ( .A(n28662), .B(n28666), .Z(n28809) );
  XNOR U34607 ( .A(n28657), .B(n28661), .Z(n28810) );
  XNOR U34608 ( .A(n28652), .B(n28656), .Z(n28811) );
  XNOR U34609 ( .A(n28647), .B(n28651), .Z(n28812) );
  XNOR U34610 ( .A(n28642), .B(n28646), .Z(n28813) );
  XNOR U34611 ( .A(n28637), .B(n28641), .Z(n28814) );
  XNOR U34612 ( .A(n28632), .B(n28636), .Z(n28815) );
  XNOR U34613 ( .A(n28627), .B(n28631), .Z(n28816) );
  XNOR U34614 ( .A(n28622), .B(n28626), .Z(n28817) );
  XNOR U34615 ( .A(n28617), .B(n28621), .Z(n28818) );
  XNOR U34616 ( .A(n28612), .B(n28616), .Z(n28819) );
  XNOR U34617 ( .A(n28607), .B(n28611), .Z(n28820) );
  XNOR U34618 ( .A(n28602), .B(n28606), .Z(n28821) );
  XNOR U34619 ( .A(n28597), .B(n28601), .Z(n28822) );
  XNOR U34620 ( .A(n28592), .B(n28596), .Z(n28823) );
  XNOR U34621 ( .A(n28587), .B(n28591), .Z(n28824) );
  XNOR U34622 ( .A(n28582), .B(n28586), .Z(n28825) );
  XNOR U34623 ( .A(n28577), .B(n28581), .Z(n28826) );
  XNOR U34624 ( .A(n28572), .B(n28576), .Z(n28827) );
  XNOR U34625 ( .A(n28567), .B(n28571), .Z(n28828) );
  XNOR U34626 ( .A(n28562), .B(n28566), .Z(n28829) );
  XNOR U34627 ( .A(n28557), .B(n28561), .Z(n28830) );
  XNOR U34628 ( .A(n28552), .B(n28556), .Z(n28831) );
  XNOR U34629 ( .A(n28547), .B(n28551), .Z(n28832) );
  XNOR U34630 ( .A(n28542), .B(n28546), .Z(n28833) );
  XNOR U34631 ( .A(n28537), .B(n28541), .Z(n28834) );
  XNOR U34632 ( .A(n28532), .B(n28536), .Z(n28835) );
  XNOR U34633 ( .A(n28527), .B(n28531), .Z(n28836) );
  XNOR U34634 ( .A(n28522), .B(n28526), .Z(n28837) );
  XNOR U34635 ( .A(n28517), .B(n28521), .Z(n28838) );
  XNOR U34636 ( .A(n28512), .B(n28516), .Z(n28839) );
  XNOR U34637 ( .A(n28507), .B(n28511), .Z(n28840) );
  XNOR U34638 ( .A(n28502), .B(n28506), .Z(n28841) );
  XNOR U34639 ( .A(n28497), .B(n28501), .Z(n28842) );
  XNOR U34640 ( .A(n28492), .B(n28496), .Z(n28843) );
  XNOR U34641 ( .A(n28487), .B(n28491), .Z(n28844) );
  XNOR U34642 ( .A(n28482), .B(n28486), .Z(n28845) );
  XNOR U34643 ( .A(n28477), .B(n28481), .Z(n28846) );
  XNOR U34644 ( .A(n28472), .B(n28476), .Z(n28847) );
  XNOR U34645 ( .A(n28467), .B(n28471), .Z(n28848) );
  XNOR U34646 ( .A(n28462), .B(n28466), .Z(n28849) );
  XNOR U34647 ( .A(n28457), .B(n28461), .Z(n28850) );
  XNOR U34648 ( .A(n28452), .B(n28456), .Z(n28851) );
  XNOR U34649 ( .A(n28447), .B(n28451), .Z(n28852) );
  XNOR U34650 ( .A(n28442), .B(n28446), .Z(n28853) );
  XNOR U34651 ( .A(n28437), .B(n28441), .Z(n28854) );
  XNOR U34652 ( .A(n28432), .B(n28436), .Z(n28855) );
  XNOR U34653 ( .A(n28427), .B(n28431), .Z(n28856) );
  XNOR U34654 ( .A(n28422), .B(n28426), .Z(n28857) );
  XNOR U34655 ( .A(n28417), .B(n28421), .Z(n28858) );
  XNOR U34656 ( .A(n28412), .B(n28416), .Z(n28859) );
  XNOR U34657 ( .A(n28407), .B(n28411), .Z(n28860) );
  XNOR U34658 ( .A(n28402), .B(n28406), .Z(n28861) );
  XNOR U34659 ( .A(n28397), .B(n28401), .Z(n28862) );
  XNOR U34660 ( .A(n28392), .B(n28396), .Z(n28863) );
  XOR U34661 ( .A(n28864), .B(n28391), .Z(n28392) );
  AND U34662 ( .A(a[0]), .B(b[80]), .Z(n28864) );
  XNOR U34663 ( .A(n28865), .B(n28391), .Z(n28393) );
  XNOR U34664 ( .A(n28866), .B(n28867), .Z(n28391) );
  ANDN U34665 ( .B(n28868), .A(n28869), .Z(n28866) );
  AND U34666 ( .A(a[1]), .B(b[79]), .Z(n28865) );
  XOR U34667 ( .A(n28871), .B(n28872), .Z(n28396) );
  ANDN U34668 ( .B(n28873), .A(n28874), .Z(n28871) );
  AND U34669 ( .A(a[2]), .B(b[78]), .Z(n28870) );
  XOR U34670 ( .A(n28876), .B(n28877), .Z(n28401) );
  ANDN U34671 ( .B(n28878), .A(n28879), .Z(n28876) );
  AND U34672 ( .A(a[3]), .B(b[77]), .Z(n28875) );
  XOR U34673 ( .A(n28881), .B(n28882), .Z(n28406) );
  ANDN U34674 ( .B(n28883), .A(n28884), .Z(n28881) );
  AND U34675 ( .A(a[4]), .B(b[76]), .Z(n28880) );
  XOR U34676 ( .A(n28886), .B(n28887), .Z(n28411) );
  ANDN U34677 ( .B(n28888), .A(n28889), .Z(n28886) );
  AND U34678 ( .A(a[5]), .B(b[75]), .Z(n28885) );
  XOR U34679 ( .A(n28891), .B(n28892), .Z(n28416) );
  ANDN U34680 ( .B(n28893), .A(n28894), .Z(n28891) );
  AND U34681 ( .A(a[6]), .B(b[74]), .Z(n28890) );
  XOR U34682 ( .A(n28896), .B(n28897), .Z(n28421) );
  ANDN U34683 ( .B(n28898), .A(n28899), .Z(n28896) );
  AND U34684 ( .A(a[7]), .B(b[73]), .Z(n28895) );
  XOR U34685 ( .A(n28901), .B(n28902), .Z(n28426) );
  ANDN U34686 ( .B(n28903), .A(n28904), .Z(n28901) );
  AND U34687 ( .A(a[8]), .B(b[72]), .Z(n28900) );
  XOR U34688 ( .A(n28906), .B(n28907), .Z(n28431) );
  ANDN U34689 ( .B(n28908), .A(n28909), .Z(n28906) );
  AND U34690 ( .A(a[9]), .B(b[71]), .Z(n28905) );
  XOR U34691 ( .A(n28911), .B(n28912), .Z(n28436) );
  ANDN U34692 ( .B(n28913), .A(n28914), .Z(n28911) );
  AND U34693 ( .A(a[10]), .B(b[70]), .Z(n28910) );
  XOR U34694 ( .A(n28916), .B(n28917), .Z(n28441) );
  ANDN U34695 ( .B(n28918), .A(n28919), .Z(n28916) );
  AND U34696 ( .A(a[11]), .B(b[69]), .Z(n28915) );
  XOR U34697 ( .A(n28921), .B(n28922), .Z(n28446) );
  ANDN U34698 ( .B(n28923), .A(n28924), .Z(n28921) );
  AND U34699 ( .A(a[12]), .B(b[68]), .Z(n28920) );
  XOR U34700 ( .A(n28926), .B(n28927), .Z(n28451) );
  ANDN U34701 ( .B(n28928), .A(n28929), .Z(n28926) );
  AND U34702 ( .A(a[13]), .B(b[67]), .Z(n28925) );
  XOR U34703 ( .A(n28931), .B(n28932), .Z(n28456) );
  ANDN U34704 ( .B(n28933), .A(n28934), .Z(n28931) );
  AND U34705 ( .A(a[14]), .B(b[66]), .Z(n28930) );
  XOR U34706 ( .A(n28936), .B(n28937), .Z(n28461) );
  ANDN U34707 ( .B(n28938), .A(n28939), .Z(n28936) );
  AND U34708 ( .A(a[15]), .B(b[65]), .Z(n28935) );
  XOR U34709 ( .A(n28941), .B(n28942), .Z(n28466) );
  ANDN U34710 ( .B(n28943), .A(n28944), .Z(n28941) );
  AND U34711 ( .A(a[16]), .B(b[64]), .Z(n28940) );
  XOR U34712 ( .A(n28946), .B(n28947), .Z(n28471) );
  ANDN U34713 ( .B(n28948), .A(n28949), .Z(n28946) );
  AND U34714 ( .A(a[17]), .B(b[63]), .Z(n28945) );
  XOR U34715 ( .A(n28951), .B(n28952), .Z(n28476) );
  ANDN U34716 ( .B(n28953), .A(n28954), .Z(n28951) );
  AND U34717 ( .A(a[18]), .B(b[62]), .Z(n28950) );
  XOR U34718 ( .A(n28956), .B(n28957), .Z(n28481) );
  ANDN U34719 ( .B(n28958), .A(n28959), .Z(n28956) );
  AND U34720 ( .A(a[19]), .B(b[61]), .Z(n28955) );
  XOR U34721 ( .A(n28961), .B(n28962), .Z(n28486) );
  ANDN U34722 ( .B(n28963), .A(n28964), .Z(n28961) );
  AND U34723 ( .A(a[20]), .B(b[60]), .Z(n28960) );
  XOR U34724 ( .A(n28966), .B(n28967), .Z(n28491) );
  ANDN U34725 ( .B(n28968), .A(n28969), .Z(n28966) );
  AND U34726 ( .A(a[21]), .B(b[59]), .Z(n28965) );
  XOR U34727 ( .A(n28971), .B(n28972), .Z(n28496) );
  ANDN U34728 ( .B(n28973), .A(n28974), .Z(n28971) );
  AND U34729 ( .A(a[22]), .B(b[58]), .Z(n28970) );
  XOR U34730 ( .A(n28976), .B(n28977), .Z(n28501) );
  ANDN U34731 ( .B(n28978), .A(n28979), .Z(n28976) );
  AND U34732 ( .A(a[23]), .B(b[57]), .Z(n28975) );
  XOR U34733 ( .A(n28981), .B(n28982), .Z(n28506) );
  ANDN U34734 ( .B(n28983), .A(n28984), .Z(n28981) );
  AND U34735 ( .A(a[24]), .B(b[56]), .Z(n28980) );
  XOR U34736 ( .A(n28986), .B(n28987), .Z(n28511) );
  ANDN U34737 ( .B(n28988), .A(n28989), .Z(n28986) );
  AND U34738 ( .A(a[25]), .B(b[55]), .Z(n28985) );
  XOR U34739 ( .A(n28991), .B(n28992), .Z(n28516) );
  ANDN U34740 ( .B(n28993), .A(n28994), .Z(n28991) );
  AND U34741 ( .A(a[26]), .B(b[54]), .Z(n28990) );
  XOR U34742 ( .A(n28996), .B(n28997), .Z(n28521) );
  ANDN U34743 ( .B(n28998), .A(n28999), .Z(n28996) );
  AND U34744 ( .A(a[27]), .B(b[53]), .Z(n28995) );
  XOR U34745 ( .A(n29001), .B(n29002), .Z(n28526) );
  ANDN U34746 ( .B(n29003), .A(n29004), .Z(n29001) );
  AND U34747 ( .A(a[28]), .B(b[52]), .Z(n29000) );
  XOR U34748 ( .A(n29006), .B(n29007), .Z(n28531) );
  ANDN U34749 ( .B(n29008), .A(n29009), .Z(n29006) );
  AND U34750 ( .A(a[29]), .B(b[51]), .Z(n29005) );
  XOR U34751 ( .A(n29011), .B(n29012), .Z(n28536) );
  ANDN U34752 ( .B(n29013), .A(n29014), .Z(n29011) );
  AND U34753 ( .A(a[30]), .B(b[50]), .Z(n29010) );
  XOR U34754 ( .A(n29016), .B(n29017), .Z(n28541) );
  ANDN U34755 ( .B(n29018), .A(n29019), .Z(n29016) );
  AND U34756 ( .A(a[31]), .B(b[49]), .Z(n29015) );
  XOR U34757 ( .A(n29021), .B(n29022), .Z(n28546) );
  ANDN U34758 ( .B(n29023), .A(n29024), .Z(n29021) );
  AND U34759 ( .A(a[32]), .B(b[48]), .Z(n29020) );
  XOR U34760 ( .A(n29026), .B(n29027), .Z(n28551) );
  ANDN U34761 ( .B(n29028), .A(n29029), .Z(n29026) );
  AND U34762 ( .A(a[33]), .B(b[47]), .Z(n29025) );
  XOR U34763 ( .A(n29031), .B(n29032), .Z(n28556) );
  ANDN U34764 ( .B(n29033), .A(n29034), .Z(n29031) );
  AND U34765 ( .A(a[34]), .B(b[46]), .Z(n29030) );
  XOR U34766 ( .A(n29036), .B(n29037), .Z(n28561) );
  ANDN U34767 ( .B(n29038), .A(n29039), .Z(n29036) );
  AND U34768 ( .A(a[35]), .B(b[45]), .Z(n29035) );
  XOR U34769 ( .A(n29041), .B(n29042), .Z(n28566) );
  ANDN U34770 ( .B(n29043), .A(n29044), .Z(n29041) );
  AND U34771 ( .A(a[36]), .B(b[44]), .Z(n29040) );
  XOR U34772 ( .A(n29046), .B(n29047), .Z(n28571) );
  ANDN U34773 ( .B(n29048), .A(n29049), .Z(n29046) );
  AND U34774 ( .A(a[37]), .B(b[43]), .Z(n29045) );
  XOR U34775 ( .A(n29051), .B(n29052), .Z(n28576) );
  ANDN U34776 ( .B(n29053), .A(n29054), .Z(n29051) );
  AND U34777 ( .A(a[38]), .B(b[42]), .Z(n29050) );
  XOR U34778 ( .A(n29056), .B(n29057), .Z(n28581) );
  ANDN U34779 ( .B(n29058), .A(n29059), .Z(n29056) );
  AND U34780 ( .A(a[39]), .B(b[41]), .Z(n29055) );
  XOR U34781 ( .A(n29061), .B(n29062), .Z(n28586) );
  ANDN U34782 ( .B(n29063), .A(n29064), .Z(n29061) );
  AND U34783 ( .A(a[40]), .B(b[40]), .Z(n29060) );
  XOR U34784 ( .A(n29066), .B(n29067), .Z(n28591) );
  ANDN U34785 ( .B(n29068), .A(n29069), .Z(n29066) );
  AND U34786 ( .A(a[41]), .B(b[39]), .Z(n29065) );
  XOR U34787 ( .A(n29071), .B(n29072), .Z(n28596) );
  ANDN U34788 ( .B(n29073), .A(n29074), .Z(n29071) );
  AND U34789 ( .A(a[42]), .B(b[38]), .Z(n29070) );
  XOR U34790 ( .A(n29076), .B(n29077), .Z(n28601) );
  ANDN U34791 ( .B(n29078), .A(n29079), .Z(n29076) );
  AND U34792 ( .A(a[43]), .B(b[37]), .Z(n29075) );
  XOR U34793 ( .A(n29081), .B(n29082), .Z(n28606) );
  ANDN U34794 ( .B(n29083), .A(n29084), .Z(n29081) );
  AND U34795 ( .A(a[44]), .B(b[36]), .Z(n29080) );
  XOR U34796 ( .A(n29086), .B(n29087), .Z(n28611) );
  ANDN U34797 ( .B(n29088), .A(n29089), .Z(n29086) );
  AND U34798 ( .A(a[45]), .B(b[35]), .Z(n29085) );
  XOR U34799 ( .A(n29091), .B(n29092), .Z(n28616) );
  ANDN U34800 ( .B(n29093), .A(n29094), .Z(n29091) );
  AND U34801 ( .A(a[46]), .B(b[34]), .Z(n29090) );
  XOR U34802 ( .A(n29096), .B(n29097), .Z(n28621) );
  ANDN U34803 ( .B(n29098), .A(n29099), .Z(n29096) );
  AND U34804 ( .A(a[47]), .B(b[33]), .Z(n29095) );
  XOR U34805 ( .A(n29101), .B(n29102), .Z(n28626) );
  ANDN U34806 ( .B(n29103), .A(n29104), .Z(n29101) );
  AND U34807 ( .A(a[48]), .B(b[32]), .Z(n29100) );
  XOR U34808 ( .A(n29106), .B(n29107), .Z(n28631) );
  ANDN U34809 ( .B(n29108), .A(n29109), .Z(n29106) );
  AND U34810 ( .A(a[49]), .B(b[31]), .Z(n29105) );
  XOR U34811 ( .A(n29111), .B(n29112), .Z(n28636) );
  ANDN U34812 ( .B(n29113), .A(n29114), .Z(n29111) );
  AND U34813 ( .A(a[50]), .B(b[30]), .Z(n29110) );
  XOR U34814 ( .A(n29116), .B(n29117), .Z(n28641) );
  ANDN U34815 ( .B(n29118), .A(n29119), .Z(n29116) );
  AND U34816 ( .A(a[51]), .B(b[29]), .Z(n29115) );
  XOR U34817 ( .A(n29121), .B(n29122), .Z(n28646) );
  ANDN U34818 ( .B(n29123), .A(n29124), .Z(n29121) );
  AND U34819 ( .A(a[52]), .B(b[28]), .Z(n29120) );
  XOR U34820 ( .A(n29126), .B(n29127), .Z(n28651) );
  ANDN U34821 ( .B(n29128), .A(n29129), .Z(n29126) );
  AND U34822 ( .A(a[53]), .B(b[27]), .Z(n29125) );
  XOR U34823 ( .A(n29131), .B(n29132), .Z(n28656) );
  ANDN U34824 ( .B(n29133), .A(n29134), .Z(n29131) );
  AND U34825 ( .A(a[54]), .B(b[26]), .Z(n29130) );
  XOR U34826 ( .A(n29136), .B(n29137), .Z(n28661) );
  ANDN U34827 ( .B(n29138), .A(n29139), .Z(n29136) );
  AND U34828 ( .A(a[55]), .B(b[25]), .Z(n29135) );
  XOR U34829 ( .A(n29141), .B(n29142), .Z(n28666) );
  ANDN U34830 ( .B(n29143), .A(n29144), .Z(n29141) );
  AND U34831 ( .A(a[56]), .B(b[24]), .Z(n29140) );
  XOR U34832 ( .A(n29146), .B(n29147), .Z(n28671) );
  ANDN U34833 ( .B(n29148), .A(n29149), .Z(n29146) );
  AND U34834 ( .A(a[57]), .B(b[23]), .Z(n29145) );
  XOR U34835 ( .A(n29151), .B(n29152), .Z(n28676) );
  ANDN U34836 ( .B(n29153), .A(n29154), .Z(n29151) );
  AND U34837 ( .A(a[58]), .B(b[22]), .Z(n29150) );
  XOR U34838 ( .A(n29156), .B(n29157), .Z(n28681) );
  ANDN U34839 ( .B(n29158), .A(n29159), .Z(n29156) );
  AND U34840 ( .A(a[59]), .B(b[21]), .Z(n29155) );
  XOR U34841 ( .A(n29161), .B(n29162), .Z(n28686) );
  ANDN U34842 ( .B(n29163), .A(n29164), .Z(n29161) );
  AND U34843 ( .A(a[60]), .B(b[20]), .Z(n29160) );
  XOR U34844 ( .A(n29166), .B(n29167), .Z(n28691) );
  ANDN U34845 ( .B(n29168), .A(n29169), .Z(n29166) );
  AND U34846 ( .A(a[61]), .B(b[19]), .Z(n29165) );
  XOR U34847 ( .A(n29171), .B(n29172), .Z(n28696) );
  ANDN U34848 ( .B(n29173), .A(n29174), .Z(n29171) );
  AND U34849 ( .A(a[62]), .B(b[18]), .Z(n29170) );
  XOR U34850 ( .A(n29176), .B(n29177), .Z(n28701) );
  ANDN U34851 ( .B(n29178), .A(n29179), .Z(n29176) );
  AND U34852 ( .A(a[63]), .B(b[17]), .Z(n29175) );
  XOR U34853 ( .A(n29181), .B(n29182), .Z(n28706) );
  ANDN U34854 ( .B(n29183), .A(n29184), .Z(n29181) );
  AND U34855 ( .A(a[64]), .B(b[16]), .Z(n29180) );
  XOR U34856 ( .A(n29186), .B(n29187), .Z(n28711) );
  ANDN U34857 ( .B(n29188), .A(n29189), .Z(n29186) );
  AND U34858 ( .A(a[65]), .B(b[15]), .Z(n29185) );
  XOR U34859 ( .A(n29191), .B(n29192), .Z(n28716) );
  ANDN U34860 ( .B(n29193), .A(n29194), .Z(n29191) );
  AND U34861 ( .A(a[66]), .B(b[14]), .Z(n29190) );
  XOR U34862 ( .A(n29196), .B(n29197), .Z(n28721) );
  ANDN U34863 ( .B(n29198), .A(n29199), .Z(n29196) );
  AND U34864 ( .A(a[67]), .B(b[13]), .Z(n29195) );
  XOR U34865 ( .A(n29201), .B(n29202), .Z(n28726) );
  ANDN U34866 ( .B(n29203), .A(n29204), .Z(n29201) );
  AND U34867 ( .A(a[68]), .B(b[12]), .Z(n29200) );
  XOR U34868 ( .A(n29206), .B(n29207), .Z(n28731) );
  ANDN U34869 ( .B(n29208), .A(n29209), .Z(n29206) );
  AND U34870 ( .A(a[69]), .B(b[11]), .Z(n29205) );
  XOR U34871 ( .A(n29211), .B(n29212), .Z(n28736) );
  ANDN U34872 ( .B(n29213), .A(n29214), .Z(n29211) );
  AND U34873 ( .A(a[70]), .B(b[10]), .Z(n29210) );
  XOR U34874 ( .A(n29216), .B(n29217), .Z(n28741) );
  ANDN U34875 ( .B(n29218), .A(n29219), .Z(n29216) );
  AND U34876 ( .A(b[9]), .B(a[71]), .Z(n29215) );
  XOR U34877 ( .A(n29221), .B(n29222), .Z(n28746) );
  ANDN U34878 ( .B(n29223), .A(n29224), .Z(n29221) );
  AND U34879 ( .A(b[8]), .B(a[72]), .Z(n29220) );
  XOR U34880 ( .A(n29226), .B(n29227), .Z(n28751) );
  ANDN U34881 ( .B(n29228), .A(n29229), .Z(n29226) );
  AND U34882 ( .A(b[7]), .B(a[73]), .Z(n29225) );
  XOR U34883 ( .A(n29231), .B(n29232), .Z(n28756) );
  ANDN U34884 ( .B(n29233), .A(n29234), .Z(n29231) );
  AND U34885 ( .A(b[6]), .B(a[74]), .Z(n29230) );
  XOR U34886 ( .A(n29236), .B(n29237), .Z(n28761) );
  ANDN U34887 ( .B(n29238), .A(n29239), .Z(n29236) );
  AND U34888 ( .A(b[5]), .B(a[75]), .Z(n29235) );
  XOR U34889 ( .A(n29241), .B(n29242), .Z(n28766) );
  ANDN U34890 ( .B(n29243), .A(n29244), .Z(n29241) );
  AND U34891 ( .A(b[4]), .B(a[76]), .Z(n29240) );
  XOR U34892 ( .A(n29246), .B(n29247), .Z(n28771) );
  ANDN U34893 ( .B(n28783), .A(n28784), .Z(n29246) );
  AND U34894 ( .A(b[2]), .B(a[77]), .Z(n29248) );
  XNOR U34895 ( .A(n29243), .B(n29247), .Z(n29249) );
  XOR U34896 ( .A(n29250), .B(n29251), .Z(n29247) );
  OR U34897 ( .A(n28786), .B(n28787), .Z(n29251) );
  XNOR U34898 ( .A(n29253), .B(n29254), .Z(n29252) );
  XOR U34899 ( .A(n29253), .B(n29256), .Z(n28786) );
  NAND U34900 ( .A(b[1]), .B(a[77]), .Z(n29256) );
  IV U34901 ( .A(n29250), .Z(n29253) );
  NANDN U34902 ( .A(n51), .B(n52), .Z(n29250) );
  XOR U34903 ( .A(n29257), .B(n29258), .Z(n52) );
  NAND U34904 ( .A(a[77]), .B(b[0]), .Z(n51) );
  XNOR U34905 ( .A(n29238), .B(n29242), .Z(n29259) );
  XNOR U34906 ( .A(n29233), .B(n29237), .Z(n29260) );
  XNOR U34907 ( .A(n29228), .B(n29232), .Z(n29261) );
  XNOR U34908 ( .A(n29223), .B(n29227), .Z(n29262) );
  XNOR U34909 ( .A(n29218), .B(n29222), .Z(n29263) );
  XNOR U34910 ( .A(n29213), .B(n29217), .Z(n29264) );
  XNOR U34911 ( .A(n29208), .B(n29212), .Z(n29265) );
  XNOR U34912 ( .A(n29203), .B(n29207), .Z(n29266) );
  XNOR U34913 ( .A(n29198), .B(n29202), .Z(n29267) );
  XNOR U34914 ( .A(n29193), .B(n29197), .Z(n29268) );
  XNOR U34915 ( .A(n29188), .B(n29192), .Z(n29269) );
  XNOR U34916 ( .A(n29183), .B(n29187), .Z(n29270) );
  XNOR U34917 ( .A(n29178), .B(n29182), .Z(n29271) );
  XNOR U34918 ( .A(n29173), .B(n29177), .Z(n29272) );
  XNOR U34919 ( .A(n29168), .B(n29172), .Z(n29273) );
  XNOR U34920 ( .A(n29163), .B(n29167), .Z(n29274) );
  XNOR U34921 ( .A(n29158), .B(n29162), .Z(n29275) );
  XNOR U34922 ( .A(n29153), .B(n29157), .Z(n29276) );
  XNOR U34923 ( .A(n29148), .B(n29152), .Z(n29277) );
  XNOR U34924 ( .A(n29143), .B(n29147), .Z(n29278) );
  XNOR U34925 ( .A(n29138), .B(n29142), .Z(n29279) );
  XNOR U34926 ( .A(n29133), .B(n29137), .Z(n29280) );
  XNOR U34927 ( .A(n29128), .B(n29132), .Z(n29281) );
  XNOR U34928 ( .A(n29123), .B(n29127), .Z(n29282) );
  XNOR U34929 ( .A(n29118), .B(n29122), .Z(n29283) );
  XNOR U34930 ( .A(n29113), .B(n29117), .Z(n29284) );
  XNOR U34931 ( .A(n29108), .B(n29112), .Z(n29285) );
  XNOR U34932 ( .A(n29103), .B(n29107), .Z(n29286) );
  XNOR U34933 ( .A(n29098), .B(n29102), .Z(n29287) );
  XNOR U34934 ( .A(n29093), .B(n29097), .Z(n29288) );
  XNOR U34935 ( .A(n29088), .B(n29092), .Z(n29289) );
  XNOR U34936 ( .A(n29083), .B(n29087), .Z(n29290) );
  XNOR U34937 ( .A(n29078), .B(n29082), .Z(n29291) );
  XNOR U34938 ( .A(n29073), .B(n29077), .Z(n29292) );
  XNOR U34939 ( .A(n29068), .B(n29072), .Z(n29293) );
  XNOR U34940 ( .A(n29063), .B(n29067), .Z(n29294) );
  XNOR U34941 ( .A(n29058), .B(n29062), .Z(n29295) );
  XNOR U34942 ( .A(n29053), .B(n29057), .Z(n29296) );
  XNOR U34943 ( .A(n29048), .B(n29052), .Z(n29297) );
  XNOR U34944 ( .A(n29043), .B(n29047), .Z(n29298) );
  XNOR U34945 ( .A(n29038), .B(n29042), .Z(n29299) );
  XNOR U34946 ( .A(n29033), .B(n29037), .Z(n29300) );
  XNOR U34947 ( .A(n29028), .B(n29032), .Z(n29301) );
  XNOR U34948 ( .A(n29023), .B(n29027), .Z(n29302) );
  XNOR U34949 ( .A(n29018), .B(n29022), .Z(n29303) );
  XNOR U34950 ( .A(n29013), .B(n29017), .Z(n29304) );
  XNOR U34951 ( .A(n29008), .B(n29012), .Z(n29305) );
  XNOR U34952 ( .A(n29003), .B(n29007), .Z(n29306) );
  XNOR U34953 ( .A(n28998), .B(n29002), .Z(n29307) );
  XNOR U34954 ( .A(n28993), .B(n28997), .Z(n29308) );
  XNOR U34955 ( .A(n28988), .B(n28992), .Z(n29309) );
  XNOR U34956 ( .A(n28983), .B(n28987), .Z(n29310) );
  XNOR U34957 ( .A(n28978), .B(n28982), .Z(n29311) );
  XNOR U34958 ( .A(n28973), .B(n28977), .Z(n29312) );
  XNOR U34959 ( .A(n28968), .B(n28972), .Z(n29313) );
  XNOR U34960 ( .A(n28963), .B(n28967), .Z(n29314) );
  XNOR U34961 ( .A(n28958), .B(n28962), .Z(n29315) );
  XNOR U34962 ( .A(n28953), .B(n28957), .Z(n29316) );
  XNOR U34963 ( .A(n28948), .B(n28952), .Z(n29317) );
  XNOR U34964 ( .A(n28943), .B(n28947), .Z(n29318) );
  XNOR U34965 ( .A(n28938), .B(n28942), .Z(n29319) );
  XNOR U34966 ( .A(n28933), .B(n28937), .Z(n29320) );
  XNOR U34967 ( .A(n28928), .B(n28932), .Z(n29321) );
  XNOR U34968 ( .A(n28923), .B(n28927), .Z(n29322) );
  XNOR U34969 ( .A(n28918), .B(n28922), .Z(n29323) );
  XNOR U34970 ( .A(n28913), .B(n28917), .Z(n29324) );
  XNOR U34971 ( .A(n28908), .B(n28912), .Z(n29325) );
  XNOR U34972 ( .A(n28903), .B(n28907), .Z(n29326) );
  XNOR U34973 ( .A(n28898), .B(n28902), .Z(n29327) );
  XNOR U34974 ( .A(n28893), .B(n28897), .Z(n29328) );
  XNOR U34975 ( .A(n28888), .B(n28892), .Z(n29329) );
  XNOR U34976 ( .A(n28883), .B(n28887), .Z(n29330) );
  XNOR U34977 ( .A(n28878), .B(n28882), .Z(n29331) );
  XNOR U34978 ( .A(n28873), .B(n28877), .Z(n29332) );
  XNOR U34979 ( .A(n28868), .B(n28872), .Z(n29333) );
  XNOR U34980 ( .A(n29334), .B(n28867), .Z(n28868) );
  AND U34981 ( .A(a[0]), .B(b[79]), .Z(n29334) );
  XOR U34982 ( .A(n29335), .B(n28867), .Z(n28869) );
  XNOR U34983 ( .A(n29336), .B(n29337), .Z(n28867) );
  ANDN U34984 ( .B(n29338), .A(n29339), .Z(n29336) );
  AND U34985 ( .A(a[1]), .B(b[78]), .Z(n29335) );
  XOR U34986 ( .A(n29341), .B(n29342), .Z(n28872) );
  ANDN U34987 ( .B(n29343), .A(n29344), .Z(n29341) );
  AND U34988 ( .A(a[2]), .B(b[77]), .Z(n29340) );
  XOR U34989 ( .A(n29346), .B(n29347), .Z(n28877) );
  ANDN U34990 ( .B(n29348), .A(n29349), .Z(n29346) );
  AND U34991 ( .A(a[3]), .B(b[76]), .Z(n29345) );
  XOR U34992 ( .A(n29351), .B(n29352), .Z(n28882) );
  ANDN U34993 ( .B(n29353), .A(n29354), .Z(n29351) );
  AND U34994 ( .A(a[4]), .B(b[75]), .Z(n29350) );
  XOR U34995 ( .A(n29356), .B(n29357), .Z(n28887) );
  ANDN U34996 ( .B(n29358), .A(n29359), .Z(n29356) );
  AND U34997 ( .A(a[5]), .B(b[74]), .Z(n29355) );
  XOR U34998 ( .A(n29361), .B(n29362), .Z(n28892) );
  ANDN U34999 ( .B(n29363), .A(n29364), .Z(n29361) );
  AND U35000 ( .A(a[6]), .B(b[73]), .Z(n29360) );
  XOR U35001 ( .A(n29366), .B(n29367), .Z(n28897) );
  ANDN U35002 ( .B(n29368), .A(n29369), .Z(n29366) );
  AND U35003 ( .A(a[7]), .B(b[72]), .Z(n29365) );
  XOR U35004 ( .A(n29371), .B(n29372), .Z(n28902) );
  ANDN U35005 ( .B(n29373), .A(n29374), .Z(n29371) );
  AND U35006 ( .A(a[8]), .B(b[71]), .Z(n29370) );
  XOR U35007 ( .A(n29376), .B(n29377), .Z(n28907) );
  ANDN U35008 ( .B(n29378), .A(n29379), .Z(n29376) );
  AND U35009 ( .A(a[9]), .B(b[70]), .Z(n29375) );
  XOR U35010 ( .A(n29381), .B(n29382), .Z(n28912) );
  ANDN U35011 ( .B(n29383), .A(n29384), .Z(n29381) );
  AND U35012 ( .A(a[10]), .B(b[69]), .Z(n29380) );
  XOR U35013 ( .A(n29386), .B(n29387), .Z(n28917) );
  ANDN U35014 ( .B(n29388), .A(n29389), .Z(n29386) );
  AND U35015 ( .A(a[11]), .B(b[68]), .Z(n29385) );
  XOR U35016 ( .A(n29391), .B(n29392), .Z(n28922) );
  ANDN U35017 ( .B(n29393), .A(n29394), .Z(n29391) );
  AND U35018 ( .A(a[12]), .B(b[67]), .Z(n29390) );
  XOR U35019 ( .A(n29396), .B(n29397), .Z(n28927) );
  ANDN U35020 ( .B(n29398), .A(n29399), .Z(n29396) );
  AND U35021 ( .A(a[13]), .B(b[66]), .Z(n29395) );
  XOR U35022 ( .A(n29401), .B(n29402), .Z(n28932) );
  ANDN U35023 ( .B(n29403), .A(n29404), .Z(n29401) );
  AND U35024 ( .A(a[14]), .B(b[65]), .Z(n29400) );
  XOR U35025 ( .A(n29406), .B(n29407), .Z(n28937) );
  ANDN U35026 ( .B(n29408), .A(n29409), .Z(n29406) );
  AND U35027 ( .A(a[15]), .B(b[64]), .Z(n29405) );
  XOR U35028 ( .A(n29411), .B(n29412), .Z(n28942) );
  ANDN U35029 ( .B(n29413), .A(n29414), .Z(n29411) );
  AND U35030 ( .A(a[16]), .B(b[63]), .Z(n29410) );
  XOR U35031 ( .A(n29416), .B(n29417), .Z(n28947) );
  ANDN U35032 ( .B(n29418), .A(n29419), .Z(n29416) );
  AND U35033 ( .A(a[17]), .B(b[62]), .Z(n29415) );
  XOR U35034 ( .A(n29421), .B(n29422), .Z(n28952) );
  ANDN U35035 ( .B(n29423), .A(n29424), .Z(n29421) );
  AND U35036 ( .A(a[18]), .B(b[61]), .Z(n29420) );
  XOR U35037 ( .A(n29426), .B(n29427), .Z(n28957) );
  ANDN U35038 ( .B(n29428), .A(n29429), .Z(n29426) );
  AND U35039 ( .A(a[19]), .B(b[60]), .Z(n29425) );
  XOR U35040 ( .A(n29431), .B(n29432), .Z(n28962) );
  ANDN U35041 ( .B(n29433), .A(n29434), .Z(n29431) );
  AND U35042 ( .A(a[20]), .B(b[59]), .Z(n29430) );
  XOR U35043 ( .A(n29436), .B(n29437), .Z(n28967) );
  ANDN U35044 ( .B(n29438), .A(n29439), .Z(n29436) );
  AND U35045 ( .A(a[21]), .B(b[58]), .Z(n29435) );
  XOR U35046 ( .A(n29441), .B(n29442), .Z(n28972) );
  ANDN U35047 ( .B(n29443), .A(n29444), .Z(n29441) );
  AND U35048 ( .A(a[22]), .B(b[57]), .Z(n29440) );
  XOR U35049 ( .A(n29446), .B(n29447), .Z(n28977) );
  ANDN U35050 ( .B(n29448), .A(n29449), .Z(n29446) );
  AND U35051 ( .A(a[23]), .B(b[56]), .Z(n29445) );
  XOR U35052 ( .A(n29451), .B(n29452), .Z(n28982) );
  ANDN U35053 ( .B(n29453), .A(n29454), .Z(n29451) );
  AND U35054 ( .A(a[24]), .B(b[55]), .Z(n29450) );
  XOR U35055 ( .A(n29456), .B(n29457), .Z(n28987) );
  ANDN U35056 ( .B(n29458), .A(n29459), .Z(n29456) );
  AND U35057 ( .A(a[25]), .B(b[54]), .Z(n29455) );
  XOR U35058 ( .A(n29461), .B(n29462), .Z(n28992) );
  ANDN U35059 ( .B(n29463), .A(n29464), .Z(n29461) );
  AND U35060 ( .A(a[26]), .B(b[53]), .Z(n29460) );
  XOR U35061 ( .A(n29466), .B(n29467), .Z(n28997) );
  ANDN U35062 ( .B(n29468), .A(n29469), .Z(n29466) );
  AND U35063 ( .A(a[27]), .B(b[52]), .Z(n29465) );
  XOR U35064 ( .A(n29471), .B(n29472), .Z(n29002) );
  ANDN U35065 ( .B(n29473), .A(n29474), .Z(n29471) );
  AND U35066 ( .A(a[28]), .B(b[51]), .Z(n29470) );
  XOR U35067 ( .A(n29476), .B(n29477), .Z(n29007) );
  ANDN U35068 ( .B(n29478), .A(n29479), .Z(n29476) );
  AND U35069 ( .A(a[29]), .B(b[50]), .Z(n29475) );
  XOR U35070 ( .A(n29481), .B(n29482), .Z(n29012) );
  ANDN U35071 ( .B(n29483), .A(n29484), .Z(n29481) );
  AND U35072 ( .A(a[30]), .B(b[49]), .Z(n29480) );
  XOR U35073 ( .A(n29486), .B(n29487), .Z(n29017) );
  ANDN U35074 ( .B(n29488), .A(n29489), .Z(n29486) );
  AND U35075 ( .A(a[31]), .B(b[48]), .Z(n29485) );
  XOR U35076 ( .A(n29491), .B(n29492), .Z(n29022) );
  ANDN U35077 ( .B(n29493), .A(n29494), .Z(n29491) );
  AND U35078 ( .A(a[32]), .B(b[47]), .Z(n29490) );
  XOR U35079 ( .A(n29496), .B(n29497), .Z(n29027) );
  ANDN U35080 ( .B(n29498), .A(n29499), .Z(n29496) );
  AND U35081 ( .A(a[33]), .B(b[46]), .Z(n29495) );
  XOR U35082 ( .A(n29501), .B(n29502), .Z(n29032) );
  ANDN U35083 ( .B(n29503), .A(n29504), .Z(n29501) );
  AND U35084 ( .A(a[34]), .B(b[45]), .Z(n29500) );
  XOR U35085 ( .A(n29506), .B(n29507), .Z(n29037) );
  ANDN U35086 ( .B(n29508), .A(n29509), .Z(n29506) );
  AND U35087 ( .A(a[35]), .B(b[44]), .Z(n29505) );
  XOR U35088 ( .A(n29511), .B(n29512), .Z(n29042) );
  ANDN U35089 ( .B(n29513), .A(n29514), .Z(n29511) );
  AND U35090 ( .A(a[36]), .B(b[43]), .Z(n29510) );
  XOR U35091 ( .A(n29516), .B(n29517), .Z(n29047) );
  ANDN U35092 ( .B(n29518), .A(n29519), .Z(n29516) );
  AND U35093 ( .A(a[37]), .B(b[42]), .Z(n29515) );
  XOR U35094 ( .A(n29521), .B(n29522), .Z(n29052) );
  ANDN U35095 ( .B(n29523), .A(n29524), .Z(n29521) );
  AND U35096 ( .A(a[38]), .B(b[41]), .Z(n29520) );
  XOR U35097 ( .A(n29526), .B(n29527), .Z(n29057) );
  ANDN U35098 ( .B(n29528), .A(n29529), .Z(n29526) );
  AND U35099 ( .A(a[39]), .B(b[40]), .Z(n29525) );
  XOR U35100 ( .A(n29531), .B(n29532), .Z(n29062) );
  ANDN U35101 ( .B(n29533), .A(n29534), .Z(n29531) );
  AND U35102 ( .A(a[40]), .B(b[39]), .Z(n29530) );
  XOR U35103 ( .A(n29536), .B(n29537), .Z(n29067) );
  ANDN U35104 ( .B(n29538), .A(n29539), .Z(n29536) );
  AND U35105 ( .A(a[41]), .B(b[38]), .Z(n29535) );
  XOR U35106 ( .A(n29541), .B(n29542), .Z(n29072) );
  ANDN U35107 ( .B(n29543), .A(n29544), .Z(n29541) );
  AND U35108 ( .A(a[42]), .B(b[37]), .Z(n29540) );
  XOR U35109 ( .A(n29546), .B(n29547), .Z(n29077) );
  ANDN U35110 ( .B(n29548), .A(n29549), .Z(n29546) );
  AND U35111 ( .A(a[43]), .B(b[36]), .Z(n29545) );
  XOR U35112 ( .A(n29551), .B(n29552), .Z(n29082) );
  ANDN U35113 ( .B(n29553), .A(n29554), .Z(n29551) );
  AND U35114 ( .A(a[44]), .B(b[35]), .Z(n29550) );
  XOR U35115 ( .A(n29556), .B(n29557), .Z(n29087) );
  ANDN U35116 ( .B(n29558), .A(n29559), .Z(n29556) );
  AND U35117 ( .A(a[45]), .B(b[34]), .Z(n29555) );
  XOR U35118 ( .A(n29561), .B(n29562), .Z(n29092) );
  ANDN U35119 ( .B(n29563), .A(n29564), .Z(n29561) );
  AND U35120 ( .A(a[46]), .B(b[33]), .Z(n29560) );
  XOR U35121 ( .A(n29566), .B(n29567), .Z(n29097) );
  ANDN U35122 ( .B(n29568), .A(n29569), .Z(n29566) );
  AND U35123 ( .A(a[47]), .B(b[32]), .Z(n29565) );
  XOR U35124 ( .A(n29571), .B(n29572), .Z(n29102) );
  ANDN U35125 ( .B(n29573), .A(n29574), .Z(n29571) );
  AND U35126 ( .A(a[48]), .B(b[31]), .Z(n29570) );
  XOR U35127 ( .A(n29576), .B(n29577), .Z(n29107) );
  ANDN U35128 ( .B(n29578), .A(n29579), .Z(n29576) );
  AND U35129 ( .A(a[49]), .B(b[30]), .Z(n29575) );
  XOR U35130 ( .A(n29581), .B(n29582), .Z(n29112) );
  ANDN U35131 ( .B(n29583), .A(n29584), .Z(n29581) );
  AND U35132 ( .A(a[50]), .B(b[29]), .Z(n29580) );
  XOR U35133 ( .A(n29586), .B(n29587), .Z(n29117) );
  ANDN U35134 ( .B(n29588), .A(n29589), .Z(n29586) );
  AND U35135 ( .A(a[51]), .B(b[28]), .Z(n29585) );
  XOR U35136 ( .A(n29591), .B(n29592), .Z(n29122) );
  ANDN U35137 ( .B(n29593), .A(n29594), .Z(n29591) );
  AND U35138 ( .A(a[52]), .B(b[27]), .Z(n29590) );
  XOR U35139 ( .A(n29596), .B(n29597), .Z(n29127) );
  ANDN U35140 ( .B(n29598), .A(n29599), .Z(n29596) );
  AND U35141 ( .A(a[53]), .B(b[26]), .Z(n29595) );
  XOR U35142 ( .A(n29601), .B(n29602), .Z(n29132) );
  ANDN U35143 ( .B(n29603), .A(n29604), .Z(n29601) );
  AND U35144 ( .A(a[54]), .B(b[25]), .Z(n29600) );
  XOR U35145 ( .A(n29606), .B(n29607), .Z(n29137) );
  ANDN U35146 ( .B(n29608), .A(n29609), .Z(n29606) );
  AND U35147 ( .A(a[55]), .B(b[24]), .Z(n29605) );
  XOR U35148 ( .A(n29611), .B(n29612), .Z(n29142) );
  ANDN U35149 ( .B(n29613), .A(n29614), .Z(n29611) );
  AND U35150 ( .A(a[56]), .B(b[23]), .Z(n29610) );
  XOR U35151 ( .A(n29616), .B(n29617), .Z(n29147) );
  ANDN U35152 ( .B(n29618), .A(n29619), .Z(n29616) );
  AND U35153 ( .A(a[57]), .B(b[22]), .Z(n29615) );
  XOR U35154 ( .A(n29621), .B(n29622), .Z(n29152) );
  ANDN U35155 ( .B(n29623), .A(n29624), .Z(n29621) );
  AND U35156 ( .A(a[58]), .B(b[21]), .Z(n29620) );
  XOR U35157 ( .A(n29626), .B(n29627), .Z(n29157) );
  ANDN U35158 ( .B(n29628), .A(n29629), .Z(n29626) );
  AND U35159 ( .A(a[59]), .B(b[20]), .Z(n29625) );
  XOR U35160 ( .A(n29631), .B(n29632), .Z(n29162) );
  ANDN U35161 ( .B(n29633), .A(n29634), .Z(n29631) );
  AND U35162 ( .A(a[60]), .B(b[19]), .Z(n29630) );
  XOR U35163 ( .A(n29636), .B(n29637), .Z(n29167) );
  ANDN U35164 ( .B(n29638), .A(n29639), .Z(n29636) );
  AND U35165 ( .A(a[61]), .B(b[18]), .Z(n29635) );
  XOR U35166 ( .A(n29641), .B(n29642), .Z(n29172) );
  ANDN U35167 ( .B(n29643), .A(n29644), .Z(n29641) );
  AND U35168 ( .A(a[62]), .B(b[17]), .Z(n29640) );
  XOR U35169 ( .A(n29646), .B(n29647), .Z(n29177) );
  ANDN U35170 ( .B(n29648), .A(n29649), .Z(n29646) );
  AND U35171 ( .A(a[63]), .B(b[16]), .Z(n29645) );
  XOR U35172 ( .A(n29651), .B(n29652), .Z(n29182) );
  ANDN U35173 ( .B(n29653), .A(n29654), .Z(n29651) );
  AND U35174 ( .A(a[64]), .B(b[15]), .Z(n29650) );
  XOR U35175 ( .A(n29656), .B(n29657), .Z(n29187) );
  ANDN U35176 ( .B(n29658), .A(n29659), .Z(n29656) );
  AND U35177 ( .A(a[65]), .B(b[14]), .Z(n29655) );
  XOR U35178 ( .A(n29661), .B(n29662), .Z(n29192) );
  ANDN U35179 ( .B(n29663), .A(n29664), .Z(n29661) );
  AND U35180 ( .A(a[66]), .B(b[13]), .Z(n29660) );
  XOR U35181 ( .A(n29666), .B(n29667), .Z(n29197) );
  ANDN U35182 ( .B(n29668), .A(n29669), .Z(n29666) );
  AND U35183 ( .A(a[67]), .B(b[12]), .Z(n29665) );
  XOR U35184 ( .A(n29671), .B(n29672), .Z(n29202) );
  ANDN U35185 ( .B(n29673), .A(n29674), .Z(n29671) );
  AND U35186 ( .A(a[68]), .B(b[11]), .Z(n29670) );
  XOR U35187 ( .A(n29676), .B(n29677), .Z(n29207) );
  ANDN U35188 ( .B(n29678), .A(n29679), .Z(n29676) );
  AND U35189 ( .A(a[69]), .B(b[10]), .Z(n29675) );
  XOR U35190 ( .A(n29681), .B(n29682), .Z(n29212) );
  ANDN U35191 ( .B(n29683), .A(n29684), .Z(n29681) );
  AND U35192 ( .A(b[9]), .B(a[70]), .Z(n29680) );
  XOR U35193 ( .A(n29686), .B(n29687), .Z(n29217) );
  ANDN U35194 ( .B(n29688), .A(n29689), .Z(n29686) );
  AND U35195 ( .A(b[8]), .B(a[71]), .Z(n29685) );
  XOR U35196 ( .A(n29691), .B(n29692), .Z(n29222) );
  ANDN U35197 ( .B(n29693), .A(n29694), .Z(n29691) );
  AND U35198 ( .A(b[7]), .B(a[72]), .Z(n29690) );
  XOR U35199 ( .A(n29696), .B(n29697), .Z(n29227) );
  ANDN U35200 ( .B(n29698), .A(n29699), .Z(n29696) );
  AND U35201 ( .A(b[6]), .B(a[73]), .Z(n29695) );
  XOR U35202 ( .A(n29701), .B(n29702), .Z(n29232) );
  ANDN U35203 ( .B(n29703), .A(n29704), .Z(n29701) );
  AND U35204 ( .A(b[5]), .B(a[74]), .Z(n29700) );
  XOR U35205 ( .A(n29706), .B(n29707), .Z(n29237) );
  ANDN U35206 ( .B(n29708), .A(n29709), .Z(n29706) );
  AND U35207 ( .A(b[4]), .B(a[75]), .Z(n29705) );
  XOR U35208 ( .A(n29711), .B(n29712), .Z(n29242) );
  ANDN U35209 ( .B(n29254), .A(n29255), .Z(n29711) );
  AND U35210 ( .A(b[2]), .B(a[76]), .Z(n29713) );
  XNOR U35211 ( .A(n29708), .B(n29712), .Z(n29714) );
  XOR U35212 ( .A(n29715), .B(n29716), .Z(n29712) );
  OR U35213 ( .A(n29257), .B(n29258), .Z(n29716) );
  XNOR U35214 ( .A(n29718), .B(n29719), .Z(n29717) );
  XOR U35215 ( .A(n29718), .B(n29721), .Z(n29257) );
  NAND U35216 ( .A(b[1]), .B(a[76]), .Z(n29721) );
  IV U35217 ( .A(n29715), .Z(n29718) );
  NANDN U35218 ( .A(n53), .B(n54), .Z(n29715) );
  XOR U35219 ( .A(n29722), .B(n29723), .Z(n54) );
  NAND U35220 ( .A(a[76]), .B(b[0]), .Z(n53) );
  XNOR U35221 ( .A(n29703), .B(n29707), .Z(n29724) );
  XNOR U35222 ( .A(n29698), .B(n29702), .Z(n29725) );
  XNOR U35223 ( .A(n29693), .B(n29697), .Z(n29726) );
  XNOR U35224 ( .A(n29688), .B(n29692), .Z(n29727) );
  XNOR U35225 ( .A(n29683), .B(n29687), .Z(n29728) );
  XNOR U35226 ( .A(n29678), .B(n29682), .Z(n29729) );
  XNOR U35227 ( .A(n29673), .B(n29677), .Z(n29730) );
  XNOR U35228 ( .A(n29668), .B(n29672), .Z(n29731) );
  XNOR U35229 ( .A(n29663), .B(n29667), .Z(n29732) );
  XNOR U35230 ( .A(n29658), .B(n29662), .Z(n29733) );
  XNOR U35231 ( .A(n29653), .B(n29657), .Z(n29734) );
  XNOR U35232 ( .A(n29648), .B(n29652), .Z(n29735) );
  XNOR U35233 ( .A(n29643), .B(n29647), .Z(n29736) );
  XNOR U35234 ( .A(n29638), .B(n29642), .Z(n29737) );
  XNOR U35235 ( .A(n29633), .B(n29637), .Z(n29738) );
  XNOR U35236 ( .A(n29628), .B(n29632), .Z(n29739) );
  XNOR U35237 ( .A(n29623), .B(n29627), .Z(n29740) );
  XNOR U35238 ( .A(n29618), .B(n29622), .Z(n29741) );
  XNOR U35239 ( .A(n29613), .B(n29617), .Z(n29742) );
  XNOR U35240 ( .A(n29608), .B(n29612), .Z(n29743) );
  XNOR U35241 ( .A(n29603), .B(n29607), .Z(n29744) );
  XNOR U35242 ( .A(n29598), .B(n29602), .Z(n29745) );
  XNOR U35243 ( .A(n29593), .B(n29597), .Z(n29746) );
  XNOR U35244 ( .A(n29588), .B(n29592), .Z(n29747) );
  XNOR U35245 ( .A(n29583), .B(n29587), .Z(n29748) );
  XNOR U35246 ( .A(n29578), .B(n29582), .Z(n29749) );
  XNOR U35247 ( .A(n29573), .B(n29577), .Z(n29750) );
  XNOR U35248 ( .A(n29568), .B(n29572), .Z(n29751) );
  XNOR U35249 ( .A(n29563), .B(n29567), .Z(n29752) );
  XNOR U35250 ( .A(n29558), .B(n29562), .Z(n29753) );
  XNOR U35251 ( .A(n29553), .B(n29557), .Z(n29754) );
  XNOR U35252 ( .A(n29548), .B(n29552), .Z(n29755) );
  XNOR U35253 ( .A(n29543), .B(n29547), .Z(n29756) );
  XNOR U35254 ( .A(n29538), .B(n29542), .Z(n29757) );
  XNOR U35255 ( .A(n29533), .B(n29537), .Z(n29758) );
  XNOR U35256 ( .A(n29528), .B(n29532), .Z(n29759) );
  XNOR U35257 ( .A(n29523), .B(n29527), .Z(n29760) );
  XNOR U35258 ( .A(n29518), .B(n29522), .Z(n29761) );
  XNOR U35259 ( .A(n29513), .B(n29517), .Z(n29762) );
  XNOR U35260 ( .A(n29508), .B(n29512), .Z(n29763) );
  XNOR U35261 ( .A(n29503), .B(n29507), .Z(n29764) );
  XNOR U35262 ( .A(n29498), .B(n29502), .Z(n29765) );
  XNOR U35263 ( .A(n29493), .B(n29497), .Z(n29766) );
  XNOR U35264 ( .A(n29488), .B(n29492), .Z(n29767) );
  XNOR U35265 ( .A(n29483), .B(n29487), .Z(n29768) );
  XNOR U35266 ( .A(n29478), .B(n29482), .Z(n29769) );
  XNOR U35267 ( .A(n29473), .B(n29477), .Z(n29770) );
  XNOR U35268 ( .A(n29468), .B(n29472), .Z(n29771) );
  XNOR U35269 ( .A(n29463), .B(n29467), .Z(n29772) );
  XNOR U35270 ( .A(n29458), .B(n29462), .Z(n29773) );
  XNOR U35271 ( .A(n29453), .B(n29457), .Z(n29774) );
  XNOR U35272 ( .A(n29448), .B(n29452), .Z(n29775) );
  XNOR U35273 ( .A(n29443), .B(n29447), .Z(n29776) );
  XNOR U35274 ( .A(n29438), .B(n29442), .Z(n29777) );
  XNOR U35275 ( .A(n29433), .B(n29437), .Z(n29778) );
  XNOR U35276 ( .A(n29428), .B(n29432), .Z(n29779) );
  XNOR U35277 ( .A(n29423), .B(n29427), .Z(n29780) );
  XNOR U35278 ( .A(n29418), .B(n29422), .Z(n29781) );
  XNOR U35279 ( .A(n29413), .B(n29417), .Z(n29782) );
  XNOR U35280 ( .A(n29408), .B(n29412), .Z(n29783) );
  XNOR U35281 ( .A(n29403), .B(n29407), .Z(n29784) );
  XNOR U35282 ( .A(n29398), .B(n29402), .Z(n29785) );
  XNOR U35283 ( .A(n29393), .B(n29397), .Z(n29786) );
  XNOR U35284 ( .A(n29388), .B(n29392), .Z(n29787) );
  XNOR U35285 ( .A(n29383), .B(n29387), .Z(n29788) );
  XNOR U35286 ( .A(n29378), .B(n29382), .Z(n29789) );
  XNOR U35287 ( .A(n29373), .B(n29377), .Z(n29790) );
  XNOR U35288 ( .A(n29368), .B(n29372), .Z(n29791) );
  XNOR U35289 ( .A(n29363), .B(n29367), .Z(n29792) );
  XNOR U35290 ( .A(n29358), .B(n29362), .Z(n29793) );
  XNOR U35291 ( .A(n29353), .B(n29357), .Z(n29794) );
  XNOR U35292 ( .A(n29348), .B(n29352), .Z(n29795) );
  XNOR U35293 ( .A(n29343), .B(n29347), .Z(n29796) );
  XNOR U35294 ( .A(n29338), .B(n29342), .Z(n29797) );
  XOR U35295 ( .A(n29798), .B(n29337), .Z(n29338) );
  AND U35296 ( .A(a[0]), .B(b[78]), .Z(n29798) );
  XNOR U35297 ( .A(n29799), .B(n29337), .Z(n29339) );
  XNOR U35298 ( .A(n29800), .B(n29801), .Z(n29337) );
  ANDN U35299 ( .B(n29802), .A(n29803), .Z(n29800) );
  AND U35300 ( .A(a[1]), .B(b[77]), .Z(n29799) );
  XOR U35301 ( .A(n29805), .B(n29806), .Z(n29342) );
  ANDN U35302 ( .B(n29807), .A(n29808), .Z(n29805) );
  AND U35303 ( .A(a[2]), .B(b[76]), .Z(n29804) );
  XOR U35304 ( .A(n29810), .B(n29811), .Z(n29347) );
  ANDN U35305 ( .B(n29812), .A(n29813), .Z(n29810) );
  AND U35306 ( .A(a[3]), .B(b[75]), .Z(n29809) );
  XOR U35307 ( .A(n29815), .B(n29816), .Z(n29352) );
  ANDN U35308 ( .B(n29817), .A(n29818), .Z(n29815) );
  AND U35309 ( .A(a[4]), .B(b[74]), .Z(n29814) );
  XOR U35310 ( .A(n29820), .B(n29821), .Z(n29357) );
  ANDN U35311 ( .B(n29822), .A(n29823), .Z(n29820) );
  AND U35312 ( .A(a[5]), .B(b[73]), .Z(n29819) );
  XOR U35313 ( .A(n29825), .B(n29826), .Z(n29362) );
  ANDN U35314 ( .B(n29827), .A(n29828), .Z(n29825) );
  AND U35315 ( .A(a[6]), .B(b[72]), .Z(n29824) );
  XOR U35316 ( .A(n29830), .B(n29831), .Z(n29367) );
  ANDN U35317 ( .B(n29832), .A(n29833), .Z(n29830) );
  AND U35318 ( .A(a[7]), .B(b[71]), .Z(n29829) );
  XOR U35319 ( .A(n29835), .B(n29836), .Z(n29372) );
  ANDN U35320 ( .B(n29837), .A(n29838), .Z(n29835) );
  AND U35321 ( .A(a[8]), .B(b[70]), .Z(n29834) );
  XOR U35322 ( .A(n29840), .B(n29841), .Z(n29377) );
  ANDN U35323 ( .B(n29842), .A(n29843), .Z(n29840) );
  AND U35324 ( .A(a[9]), .B(b[69]), .Z(n29839) );
  XOR U35325 ( .A(n29845), .B(n29846), .Z(n29382) );
  ANDN U35326 ( .B(n29847), .A(n29848), .Z(n29845) );
  AND U35327 ( .A(a[10]), .B(b[68]), .Z(n29844) );
  XOR U35328 ( .A(n29850), .B(n29851), .Z(n29387) );
  ANDN U35329 ( .B(n29852), .A(n29853), .Z(n29850) );
  AND U35330 ( .A(a[11]), .B(b[67]), .Z(n29849) );
  XOR U35331 ( .A(n29855), .B(n29856), .Z(n29392) );
  ANDN U35332 ( .B(n29857), .A(n29858), .Z(n29855) );
  AND U35333 ( .A(a[12]), .B(b[66]), .Z(n29854) );
  XOR U35334 ( .A(n29860), .B(n29861), .Z(n29397) );
  ANDN U35335 ( .B(n29862), .A(n29863), .Z(n29860) );
  AND U35336 ( .A(a[13]), .B(b[65]), .Z(n29859) );
  XOR U35337 ( .A(n29865), .B(n29866), .Z(n29402) );
  ANDN U35338 ( .B(n29867), .A(n29868), .Z(n29865) );
  AND U35339 ( .A(a[14]), .B(b[64]), .Z(n29864) );
  XOR U35340 ( .A(n29870), .B(n29871), .Z(n29407) );
  ANDN U35341 ( .B(n29872), .A(n29873), .Z(n29870) );
  AND U35342 ( .A(a[15]), .B(b[63]), .Z(n29869) );
  XOR U35343 ( .A(n29875), .B(n29876), .Z(n29412) );
  ANDN U35344 ( .B(n29877), .A(n29878), .Z(n29875) );
  AND U35345 ( .A(a[16]), .B(b[62]), .Z(n29874) );
  XOR U35346 ( .A(n29880), .B(n29881), .Z(n29417) );
  ANDN U35347 ( .B(n29882), .A(n29883), .Z(n29880) );
  AND U35348 ( .A(a[17]), .B(b[61]), .Z(n29879) );
  XOR U35349 ( .A(n29885), .B(n29886), .Z(n29422) );
  ANDN U35350 ( .B(n29887), .A(n29888), .Z(n29885) );
  AND U35351 ( .A(a[18]), .B(b[60]), .Z(n29884) );
  XOR U35352 ( .A(n29890), .B(n29891), .Z(n29427) );
  ANDN U35353 ( .B(n29892), .A(n29893), .Z(n29890) );
  AND U35354 ( .A(a[19]), .B(b[59]), .Z(n29889) );
  XOR U35355 ( .A(n29895), .B(n29896), .Z(n29432) );
  ANDN U35356 ( .B(n29897), .A(n29898), .Z(n29895) );
  AND U35357 ( .A(a[20]), .B(b[58]), .Z(n29894) );
  XOR U35358 ( .A(n29900), .B(n29901), .Z(n29437) );
  ANDN U35359 ( .B(n29902), .A(n29903), .Z(n29900) );
  AND U35360 ( .A(a[21]), .B(b[57]), .Z(n29899) );
  XOR U35361 ( .A(n29905), .B(n29906), .Z(n29442) );
  ANDN U35362 ( .B(n29907), .A(n29908), .Z(n29905) );
  AND U35363 ( .A(a[22]), .B(b[56]), .Z(n29904) );
  XOR U35364 ( .A(n29910), .B(n29911), .Z(n29447) );
  ANDN U35365 ( .B(n29912), .A(n29913), .Z(n29910) );
  AND U35366 ( .A(a[23]), .B(b[55]), .Z(n29909) );
  XOR U35367 ( .A(n29915), .B(n29916), .Z(n29452) );
  ANDN U35368 ( .B(n29917), .A(n29918), .Z(n29915) );
  AND U35369 ( .A(a[24]), .B(b[54]), .Z(n29914) );
  XOR U35370 ( .A(n29920), .B(n29921), .Z(n29457) );
  ANDN U35371 ( .B(n29922), .A(n29923), .Z(n29920) );
  AND U35372 ( .A(a[25]), .B(b[53]), .Z(n29919) );
  XOR U35373 ( .A(n29925), .B(n29926), .Z(n29462) );
  ANDN U35374 ( .B(n29927), .A(n29928), .Z(n29925) );
  AND U35375 ( .A(a[26]), .B(b[52]), .Z(n29924) );
  XOR U35376 ( .A(n29930), .B(n29931), .Z(n29467) );
  ANDN U35377 ( .B(n29932), .A(n29933), .Z(n29930) );
  AND U35378 ( .A(a[27]), .B(b[51]), .Z(n29929) );
  XOR U35379 ( .A(n29935), .B(n29936), .Z(n29472) );
  ANDN U35380 ( .B(n29937), .A(n29938), .Z(n29935) );
  AND U35381 ( .A(a[28]), .B(b[50]), .Z(n29934) );
  XOR U35382 ( .A(n29940), .B(n29941), .Z(n29477) );
  ANDN U35383 ( .B(n29942), .A(n29943), .Z(n29940) );
  AND U35384 ( .A(a[29]), .B(b[49]), .Z(n29939) );
  XOR U35385 ( .A(n29945), .B(n29946), .Z(n29482) );
  ANDN U35386 ( .B(n29947), .A(n29948), .Z(n29945) );
  AND U35387 ( .A(a[30]), .B(b[48]), .Z(n29944) );
  XOR U35388 ( .A(n29950), .B(n29951), .Z(n29487) );
  ANDN U35389 ( .B(n29952), .A(n29953), .Z(n29950) );
  AND U35390 ( .A(a[31]), .B(b[47]), .Z(n29949) );
  XOR U35391 ( .A(n29955), .B(n29956), .Z(n29492) );
  ANDN U35392 ( .B(n29957), .A(n29958), .Z(n29955) );
  AND U35393 ( .A(a[32]), .B(b[46]), .Z(n29954) );
  XOR U35394 ( .A(n29960), .B(n29961), .Z(n29497) );
  ANDN U35395 ( .B(n29962), .A(n29963), .Z(n29960) );
  AND U35396 ( .A(a[33]), .B(b[45]), .Z(n29959) );
  XOR U35397 ( .A(n29965), .B(n29966), .Z(n29502) );
  ANDN U35398 ( .B(n29967), .A(n29968), .Z(n29965) );
  AND U35399 ( .A(a[34]), .B(b[44]), .Z(n29964) );
  XOR U35400 ( .A(n29970), .B(n29971), .Z(n29507) );
  ANDN U35401 ( .B(n29972), .A(n29973), .Z(n29970) );
  AND U35402 ( .A(a[35]), .B(b[43]), .Z(n29969) );
  XOR U35403 ( .A(n29975), .B(n29976), .Z(n29512) );
  ANDN U35404 ( .B(n29977), .A(n29978), .Z(n29975) );
  AND U35405 ( .A(a[36]), .B(b[42]), .Z(n29974) );
  XOR U35406 ( .A(n29980), .B(n29981), .Z(n29517) );
  ANDN U35407 ( .B(n29982), .A(n29983), .Z(n29980) );
  AND U35408 ( .A(a[37]), .B(b[41]), .Z(n29979) );
  XOR U35409 ( .A(n29985), .B(n29986), .Z(n29522) );
  ANDN U35410 ( .B(n29987), .A(n29988), .Z(n29985) );
  AND U35411 ( .A(a[38]), .B(b[40]), .Z(n29984) );
  XOR U35412 ( .A(n29990), .B(n29991), .Z(n29527) );
  ANDN U35413 ( .B(n29992), .A(n29993), .Z(n29990) );
  AND U35414 ( .A(a[39]), .B(b[39]), .Z(n29989) );
  XOR U35415 ( .A(n29995), .B(n29996), .Z(n29532) );
  ANDN U35416 ( .B(n29997), .A(n29998), .Z(n29995) );
  AND U35417 ( .A(a[40]), .B(b[38]), .Z(n29994) );
  XOR U35418 ( .A(n30000), .B(n30001), .Z(n29537) );
  ANDN U35419 ( .B(n30002), .A(n30003), .Z(n30000) );
  AND U35420 ( .A(a[41]), .B(b[37]), .Z(n29999) );
  XOR U35421 ( .A(n30005), .B(n30006), .Z(n29542) );
  ANDN U35422 ( .B(n30007), .A(n30008), .Z(n30005) );
  AND U35423 ( .A(a[42]), .B(b[36]), .Z(n30004) );
  XOR U35424 ( .A(n30010), .B(n30011), .Z(n29547) );
  ANDN U35425 ( .B(n30012), .A(n30013), .Z(n30010) );
  AND U35426 ( .A(a[43]), .B(b[35]), .Z(n30009) );
  XOR U35427 ( .A(n30015), .B(n30016), .Z(n29552) );
  ANDN U35428 ( .B(n30017), .A(n30018), .Z(n30015) );
  AND U35429 ( .A(a[44]), .B(b[34]), .Z(n30014) );
  XOR U35430 ( .A(n30020), .B(n30021), .Z(n29557) );
  ANDN U35431 ( .B(n30022), .A(n30023), .Z(n30020) );
  AND U35432 ( .A(a[45]), .B(b[33]), .Z(n30019) );
  XOR U35433 ( .A(n30025), .B(n30026), .Z(n29562) );
  ANDN U35434 ( .B(n30027), .A(n30028), .Z(n30025) );
  AND U35435 ( .A(a[46]), .B(b[32]), .Z(n30024) );
  XOR U35436 ( .A(n30030), .B(n30031), .Z(n29567) );
  ANDN U35437 ( .B(n30032), .A(n30033), .Z(n30030) );
  AND U35438 ( .A(a[47]), .B(b[31]), .Z(n30029) );
  XOR U35439 ( .A(n30035), .B(n30036), .Z(n29572) );
  ANDN U35440 ( .B(n30037), .A(n30038), .Z(n30035) );
  AND U35441 ( .A(a[48]), .B(b[30]), .Z(n30034) );
  XOR U35442 ( .A(n30040), .B(n30041), .Z(n29577) );
  ANDN U35443 ( .B(n30042), .A(n30043), .Z(n30040) );
  AND U35444 ( .A(a[49]), .B(b[29]), .Z(n30039) );
  XOR U35445 ( .A(n30045), .B(n30046), .Z(n29582) );
  ANDN U35446 ( .B(n30047), .A(n30048), .Z(n30045) );
  AND U35447 ( .A(a[50]), .B(b[28]), .Z(n30044) );
  XOR U35448 ( .A(n30050), .B(n30051), .Z(n29587) );
  ANDN U35449 ( .B(n30052), .A(n30053), .Z(n30050) );
  AND U35450 ( .A(a[51]), .B(b[27]), .Z(n30049) );
  XOR U35451 ( .A(n30055), .B(n30056), .Z(n29592) );
  ANDN U35452 ( .B(n30057), .A(n30058), .Z(n30055) );
  AND U35453 ( .A(a[52]), .B(b[26]), .Z(n30054) );
  XOR U35454 ( .A(n30060), .B(n30061), .Z(n29597) );
  ANDN U35455 ( .B(n30062), .A(n30063), .Z(n30060) );
  AND U35456 ( .A(a[53]), .B(b[25]), .Z(n30059) );
  XOR U35457 ( .A(n30065), .B(n30066), .Z(n29602) );
  ANDN U35458 ( .B(n30067), .A(n30068), .Z(n30065) );
  AND U35459 ( .A(a[54]), .B(b[24]), .Z(n30064) );
  XOR U35460 ( .A(n30070), .B(n30071), .Z(n29607) );
  ANDN U35461 ( .B(n30072), .A(n30073), .Z(n30070) );
  AND U35462 ( .A(a[55]), .B(b[23]), .Z(n30069) );
  XOR U35463 ( .A(n30075), .B(n30076), .Z(n29612) );
  ANDN U35464 ( .B(n30077), .A(n30078), .Z(n30075) );
  AND U35465 ( .A(a[56]), .B(b[22]), .Z(n30074) );
  XOR U35466 ( .A(n30080), .B(n30081), .Z(n29617) );
  ANDN U35467 ( .B(n30082), .A(n30083), .Z(n30080) );
  AND U35468 ( .A(a[57]), .B(b[21]), .Z(n30079) );
  XOR U35469 ( .A(n30085), .B(n30086), .Z(n29622) );
  ANDN U35470 ( .B(n30087), .A(n30088), .Z(n30085) );
  AND U35471 ( .A(a[58]), .B(b[20]), .Z(n30084) );
  XOR U35472 ( .A(n30090), .B(n30091), .Z(n29627) );
  ANDN U35473 ( .B(n30092), .A(n30093), .Z(n30090) );
  AND U35474 ( .A(a[59]), .B(b[19]), .Z(n30089) );
  XOR U35475 ( .A(n30095), .B(n30096), .Z(n29632) );
  ANDN U35476 ( .B(n30097), .A(n30098), .Z(n30095) );
  AND U35477 ( .A(a[60]), .B(b[18]), .Z(n30094) );
  XOR U35478 ( .A(n30100), .B(n30101), .Z(n29637) );
  ANDN U35479 ( .B(n30102), .A(n30103), .Z(n30100) );
  AND U35480 ( .A(a[61]), .B(b[17]), .Z(n30099) );
  XOR U35481 ( .A(n30105), .B(n30106), .Z(n29642) );
  ANDN U35482 ( .B(n30107), .A(n30108), .Z(n30105) );
  AND U35483 ( .A(a[62]), .B(b[16]), .Z(n30104) );
  XOR U35484 ( .A(n30110), .B(n30111), .Z(n29647) );
  ANDN U35485 ( .B(n30112), .A(n30113), .Z(n30110) );
  AND U35486 ( .A(a[63]), .B(b[15]), .Z(n30109) );
  XOR U35487 ( .A(n30115), .B(n30116), .Z(n29652) );
  ANDN U35488 ( .B(n30117), .A(n30118), .Z(n30115) );
  AND U35489 ( .A(a[64]), .B(b[14]), .Z(n30114) );
  XOR U35490 ( .A(n30120), .B(n30121), .Z(n29657) );
  ANDN U35491 ( .B(n30122), .A(n30123), .Z(n30120) );
  AND U35492 ( .A(a[65]), .B(b[13]), .Z(n30119) );
  XOR U35493 ( .A(n30125), .B(n30126), .Z(n29662) );
  ANDN U35494 ( .B(n30127), .A(n30128), .Z(n30125) );
  AND U35495 ( .A(a[66]), .B(b[12]), .Z(n30124) );
  XOR U35496 ( .A(n30130), .B(n30131), .Z(n29667) );
  ANDN U35497 ( .B(n30132), .A(n30133), .Z(n30130) );
  AND U35498 ( .A(a[67]), .B(b[11]), .Z(n30129) );
  XOR U35499 ( .A(n30135), .B(n30136), .Z(n29672) );
  ANDN U35500 ( .B(n30137), .A(n30138), .Z(n30135) );
  AND U35501 ( .A(a[68]), .B(b[10]), .Z(n30134) );
  XOR U35502 ( .A(n30140), .B(n30141), .Z(n29677) );
  ANDN U35503 ( .B(n30142), .A(n30143), .Z(n30140) );
  AND U35504 ( .A(b[9]), .B(a[69]), .Z(n30139) );
  XOR U35505 ( .A(n30145), .B(n30146), .Z(n29682) );
  ANDN U35506 ( .B(n30147), .A(n30148), .Z(n30145) );
  AND U35507 ( .A(b[8]), .B(a[70]), .Z(n30144) );
  XOR U35508 ( .A(n30150), .B(n30151), .Z(n29687) );
  ANDN U35509 ( .B(n30152), .A(n30153), .Z(n30150) );
  AND U35510 ( .A(b[7]), .B(a[71]), .Z(n30149) );
  XOR U35511 ( .A(n30155), .B(n30156), .Z(n29692) );
  ANDN U35512 ( .B(n30157), .A(n30158), .Z(n30155) );
  AND U35513 ( .A(b[6]), .B(a[72]), .Z(n30154) );
  XOR U35514 ( .A(n30160), .B(n30161), .Z(n29697) );
  ANDN U35515 ( .B(n30162), .A(n30163), .Z(n30160) );
  AND U35516 ( .A(b[5]), .B(a[73]), .Z(n30159) );
  XOR U35517 ( .A(n30165), .B(n30166), .Z(n29702) );
  ANDN U35518 ( .B(n30167), .A(n30168), .Z(n30165) );
  AND U35519 ( .A(b[4]), .B(a[74]), .Z(n30164) );
  XOR U35520 ( .A(n30170), .B(n30171), .Z(n29707) );
  ANDN U35521 ( .B(n29719), .A(n29720), .Z(n30170) );
  AND U35522 ( .A(b[2]), .B(a[75]), .Z(n30172) );
  XNOR U35523 ( .A(n30167), .B(n30171), .Z(n30173) );
  XOR U35524 ( .A(n30174), .B(n30175), .Z(n30171) );
  OR U35525 ( .A(n29722), .B(n29723), .Z(n30175) );
  XNOR U35526 ( .A(n30177), .B(n30178), .Z(n30176) );
  XOR U35527 ( .A(n30177), .B(n30180), .Z(n29722) );
  NAND U35528 ( .A(b[1]), .B(a[75]), .Z(n30180) );
  IV U35529 ( .A(n30174), .Z(n30177) );
  NANDN U35530 ( .A(n55), .B(n56), .Z(n30174) );
  XOR U35531 ( .A(n30181), .B(n30182), .Z(n56) );
  NAND U35532 ( .A(a[75]), .B(b[0]), .Z(n55) );
  XNOR U35533 ( .A(n30162), .B(n30166), .Z(n30183) );
  XNOR U35534 ( .A(n30157), .B(n30161), .Z(n30184) );
  XNOR U35535 ( .A(n30152), .B(n30156), .Z(n30185) );
  XNOR U35536 ( .A(n30147), .B(n30151), .Z(n30186) );
  XNOR U35537 ( .A(n30142), .B(n30146), .Z(n30187) );
  XNOR U35538 ( .A(n30137), .B(n30141), .Z(n30188) );
  XNOR U35539 ( .A(n30132), .B(n30136), .Z(n30189) );
  XNOR U35540 ( .A(n30127), .B(n30131), .Z(n30190) );
  XNOR U35541 ( .A(n30122), .B(n30126), .Z(n30191) );
  XNOR U35542 ( .A(n30117), .B(n30121), .Z(n30192) );
  XNOR U35543 ( .A(n30112), .B(n30116), .Z(n30193) );
  XNOR U35544 ( .A(n30107), .B(n30111), .Z(n30194) );
  XNOR U35545 ( .A(n30102), .B(n30106), .Z(n30195) );
  XNOR U35546 ( .A(n30097), .B(n30101), .Z(n30196) );
  XNOR U35547 ( .A(n30092), .B(n30096), .Z(n30197) );
  XNOR U35548 ( .A(n30087), .B(n30091), .Z(n30198) );
  XNOR U35549 ( .A(n30082), .B(n30086), .Z(n30199) );
  XNOR U35550 ( .A(n30077), .B(n30081), .Z(n30200) );
  XNOR U35551 ( .A(n30072), .B(n30076), .Z(n30201) );
  XNOR U35552 ( .A(n30067), .B(n30071), .Z(n30202) );
  XNOR U35553 ( .A(n30062), .B(n30066), .Z(n30203) );
  XNOR U35554 ( .A(n30057), .B(n30061), .Z(n30204) );
  XNOR U35555 ( .A(n30052), .B(n30056), .Z(n30205) );
  XNOR U35556 ( .A(n30047), .B(n30051), .Z(n30206) );
  XNOR U35557 ( .A(n30042), .B(n30046), .Z(n30207) );
  XNOR U35558 ( .A(n30037), .B(n30041), .Z(n30208) );
  XNOR U35559 ( .A(n30032), .B(n30036), .Z(n30209) );
  XNOR U35560 ( .A(n30027), .B(n30031), .Z(n30210) );
  XNOR U35561 ( .A(n30022), .B(n30026), .Z(n30211) );
  XNOR U35562 ( .A(n30017), .B(n30021), .Z(n30212) );
  XNOR U35563 ( .A(n30012), .B(n30016), .Z(n30213) );
  XNOR U35564 ( .A(n30007), .B(n30011), .Z(n30214) );
  XNOR U35565 ( .A(n30002), .B(n30006), .Z(n30215) );
  XNOR U35566 ( .A(n29997), .B(n30001), .Z(n30216) );
  XNOR U35567 ( .A(n29992), .B(n29996), .Z(n30217) );
  XNOR U35568 ( .A(n29987), .B(n29991), .Z(n30218) );
  XNOR U35569 ( .A(n29982), .B(n29986), .Z(n30219) );
  XNOR U35570 ( .A(n29977), .B(n29981), .Z(n30220) );
  XNOR U35571 ( .A(n29972), .B(n29976), .Z(n30221) );
  XNOR U35572 ( .A(n29967), .B(n29971), .Z(n30222) );
  XNOR U35573 ( .A(n29962), .B(n29966), .Z(n30223) );
  XNOR U35574 ( .A(n29957), .B(n29961), .Z(n30224) );
  XNOR U35575 ( .A(n29952), .B(n29956), .Z(n30225) );
  XNOR U35576 ( .A(n29947), .B(n29951), .Z(n30226) );
  XNOR U35577 ( .A(n29942), .B(n29946), .Z(n30227) );
  XNOR U35578 ( .A(n29937), .B(n29941), .Z(n30228) );
  XNOR U35579 ( .A(n29932), .B(n29936), .Z(n30229) );
  XNOR U35580 ( .A(n29927), .B(n29931), .Z(n30230) );
  XNOR U35581 ( .A(n29922), .B(n29926), .Z(n30231) );
  XNOR U35582 ( .A(n29917), .B(n29921), .Z(n30232) );
  XNOR U35583 ( .A(n29912), .B(n29916), .Z(n30233) );
  XNOR U35584 ( .A(n29907), .B(n29911), .Z(n30234) );
  XNOR U35585 ( .A(n29902), .B(n29906), .Z(n30235) );
  XNOR U35586 ( .A(n29897), .B(n29901), .Z(n30236) );
  XNOR U35587 ( .A(n29892), .B(n29896), .Z(n30237) );
  XNOR U35588 ( .A(n29887), .B(n29891), .Z(n30238) );
  XNOR U35589 ( .A(n29882), .B(n29886), .Z(n30239) );
  XNOR U35590 ( .A(n29877), .B(n29881), .Z(n30240) );
  XNOR U35591 ( .A(n29872), .B(n29876), .Z(n30241) );
  XNOR U35592 ( .A(n29867), .B(n29871), .Z(n30242) );
  XNOR U35593 ( .A(n29862), .B(n29866), .Z(n30243) );
  XNOR U35594 ( .A(n29857), .B(n29861), .Z(n30244) );
  XNOR U35595 ( .A(n29852), .B(n29856), .Z(n30245) );
  XNOR U35596 ( .A(n29847), .B(n29851), .Z(n30246) );
  XNOR U35597 ( .A(n29842), .B(n29846), .Z(n30247) );
  XNOR U35598 ( .A(n29837), .B(n29841), .Z(n30248) );
  XNOR U35599 ( .A(n29832), .B(n29836), .Z(n30249) );
  XNOR U35600 ( .A(n29827), .B(n29831), .Z(n30250) );
  XNOR U35601 ( .A(n29822), .B(n29826), .Z(n30251) );
  XNOR U35602 ( .A(n29817), .B(n29821), .Z(n30252) );
  XNOR U35603 ( .A(n29812), .B(n29816), .Z(n30253) );
  XNOR U35604 ( .A(n29807), .B(n29811), .Z(n30254) );
  XNOR U35605 ( .A(n29802), .B(n29806), .Z(n30255) );
  XNOR U35606 ( .A(n30256), .B(n29801), .Z(n29802) );
  AND U35607 ( .A(a[0]), .B(b[77]), .Z(n30256) );
  XOR U35608 ( .A(n30257), .B(n29801), .Z(n29803) );
  XNOR U35609 ( .A(n30258), .B(n30259), .Z(n29801) );
  ANDN U35610 ( .B(n30260), .A(n30261), .Z(n30258) );
  AND U35611 ( .A(a[1]), .B(b[76]), .Z(n30257) );
  XOR U35612 ( .A(n30263), .B(n30264), .Z(n29806) );
  ANDN U35613 ( .B(n30265), .A(n30266), .Z(n30263) );
  AND U35614 ( .A(a[2]), .B(b[75]), .Z(n30262) );
  XOR U35615 ( .A(n30268), .B(n30269), .Z(n29811) );
  ANDN U35616 ( .B(n30270), .A(n30271), .Z(n30268) );
  AND U35617 ( .A(a[3]), .B(b[74]), .Z(n30267) );
  XOR U35618 ( .A(n30273), .B(n30274), .Z(n29816) );
  ANDN U35619 ( .B(n30275), .A(n30276), .Z(n30273) );
  AND U35620 ( .A(a[4]), .B(b[73]), .Z(n30272) );
  XOR U35621 ( .A(n30278), .B(n30279), .Z(n29821) );
  ANDN U35622 ( .B(n30280), .A(n30281), .Z(n30278) );
  AND U35623 ( .A(a[5]), .B(b[72]), .Z(n30277) );
  XOR U35624 ( .A(n30283), .B(n30284), .Z(n29826) );
  ANDN U35625 ( .B(n30285), .A(n30286), .Z(n30283) );
  AND U35626 ( .A(a[6]), .B(b[71]), .Z(n30282) );
  XOR U35627 ( .A(n30288), .B(n30289), .Z(n29831) );
  ANDN U35628 ( .B(n30290), .A(n30291), .Z(n30288) );
  AND U35629 ( .A(a[7]), .B(b[70]), .Z(n30287) );
  XOR U35630 ( .A(n30293), .B(n30294), .Z(n29836) );
  ANDN U35631 ( .B(n30295), .A(n30296), .Z(n30293) );
  AND U35632 ( .A(a[8]), .B(b[69]), .Z(n30292) );
  XOR U35633 ( .A(n30298), .B(n30299), .Z(n29841) );
  ANDN U35634 ( .B(n30300), .A(n30301), .Z(n30298) );
  AND U35635 ( .A(a[9]), .B(b[68]), .Z(n30297) );
  XOR U35636 ( .A(n30303), .B(n30304), .Z(n29846) );
  ANDN U35637 ( .B(n30305), .A(n30306), .Z(n30303) );
  AND U35638 ( .A(a[10]), .B(b[67]), .Z(n30302) );
  XOR U35639 ( .A(n30308), .B(n30309), .Z(n29851) );
  ANDN U35640 ( .B(n30310), .A(n30311), .Z(n30308) );
  AND U35641 ( .A(a[11]), .B(b[66]), .Z(n30307) );
  XOR U35642 ( .A(n30313), .B(n30314), .Z(n29856) );
  ANDN U35643 ( .B(n30315), .A(n30316), .Z(n30313) );
  AND U35644 ( .A(a[12]), .B(b[65]), .Z(n30312) );
  XOR U35645 ( .A(n30318), .B(n30319), .Z(n29861) );
  ANDN U35646 ( .B(n30320), .A(n30321), .Z(n30318) );
  AND U35647 ( .A(a[13]), .B(b[64]), .Z(n30317) );
  XOR U35648 ( .A(n30323), .B(n30324), .Z(n29866) );
  ANDN U35649 ( .B(n30325), .A(n30326), .Z(n30323) );
  AND U35650 ( .A(a[14]), .B(b[63]), .Z(n30322) );
  XOR U35651 ( .A(n30328), .B(n30329), .Z(n29871) );
  ANDN U35652 ( .B(n30330), .A(n30331), .Z(n30328) );
  AND U35653 ( .A(a[15]), .B(b[62]), .Z(n30327) );
  XOR U35654 ( .A(n30333), .B(n30334), .Z(n29876) );
  ANDN U35655 ( .B(n30335), .A(n30336), .Z(n30333) );
  AND U35656 ( .A(a[16]), .B(b[61]), .Z(n30332) );
  XOR U35657 ( .A(n30338), .B(n30339), .Z(n29881) );
  ANDN U35658 ( .B(n30340), .A(n30341), .Z(n30338) );
  AND U35659 ( .A(a[17]), .B(b[60]), .Z(n30337) );
  XOR U35660 ( .A(n30343), .B(n30344), .Z(n29886) );
  ANDN U35661 ( .B(n30345), .A(n30346), .Z(n30343) );
  AND U35662 ( .A(a[18]), .B(b[59]), .Z(n30342) );
  XOR U35663 ( .A(n30348), .B(n30349), .Z(n29891) );
  ANDN U35664 ( .B(n30350), .A(n30351), .Z(n30348) );
  AND U35665 ( .A(a[19]), .B(b[58]), .Z(n30347) );
  XOR U35666 ( .A(n30353), .B(n30354), .Z(n29896) );
  ANDN U35667 ( .B(n30355), .A(n30356), .Z(n30353) );
  AND U35668 ( .A(a[20]), .B(b[57]), .Z(n30352) );
  XOR U35669 ( .A(n30358), .B(n30359), .Z(n29901) );
  ANDN U35670 ( .B(n30360), .A(n30361), .Z(n30358) );
  AND U35671 ( .A(a[21]), .B(b[56]), .Z(n30357) );
  XOR U35672 ( .A(n30363), .B(n30364), .Z(n29906) );
  ANDN U35673 ( .B(n30365), .A(n30366), .Z(n30363) );
  AND U35674 ( .A(a[22]), .B(b[55]), .Z(n30362) );
  XOR U35675 ( .A(n30368), .B(n30369), .Z(n29911) );
  ANDN U35676 ( .B(n30370), .A(n30371), .Z(n30368) );
  AND U35677 ( .A(a[23]), .B(b[54]), .Z(n30367) );
  XOR U35678 ( .A(n30373), .B(n30374), .Z(n29916) );
  ANDN U35679 ( .B(n30375), .A(n30376), .Z(n30373) );
  AND U35680 ( .A(a[24]), .B(b[53]), .Z(n30372) );
  XOR U35681 ( .A(n30378), .B(n30379), .Z(n29921) );
  ANDN U35682 ( .B(n30380), .A(n30381), .Z(n30378) );
  AND U35683 ( .A(a[25]), .B(b[52]), .Z(n30377) );
  XOR U35684 ( .A(n30383), .B(n30384), .Z(n29926) );
  ANDN U35685 ( .B(n30385), .A(n30386), .Z(n30383) );
  AND U35686 ( .A(a[26]), .B(b[51]), .Z(n30382) );
  XOR U35687 ( .A(n30388), .B(n30389), .Z(n29931) );
  ANDN U35688 ( .B(n30390), .A(n30391), .Z(n30388) );
  AND U35689 ( .A(a[27]), .B(b[50]), .Z(n30387) );
  XOR U35690 ( .A(n30393), .B(n30394), .Z(n29936) );
  ANDN U35691 ( .B(n30395), .A(n30396), .Z(n30393) );
  AND U35692 ( .A(a[28]), .B(b[49]), .Z(n30392) );
  XOR U35693 ( .A(n30398), .B(n30399), .Z(n29941) );
  ANDN U35694 ( .B(n30400), .A(n30401), .Z(n30398) );
  AND U35695 ( .A(a[29]), .B(b[48]), .Z(n30397) );
  XOR U35696 ( .A(n30403), .B(n30404), .Z(n29946) );
  ANDN U35697 ( .B(n30405), .A(n30406), .Z(n30403) );
  AND U35698 ( .A(a[30]), .B(b[47]), .Z(n30402) );
  XOR U35699 ( .A(n30408), .B(n30409), .Z(n29951) );
  ANDN U35700 ( .B(n30410), .A(n30411), .Z(n30408) );
  AND U35701 ( .A(a[31]), .B(b[46]), .Z(n30407) );
  XOR U35702 ( .A(n30413), .B(n30414), .Z(n29956) );
  ANDN U35703 ( .B(n30415), .A(n30416), .Z(n30413) );
  AND U35704 ( .A(a[32]), .B(b[45]), .Z(n30412) );
  XOR U35705 ( .A(n30418), .B(n30419), .Z(n29961) );
  ANDN U35706 ( .B(n30420), .A(n30421), .Z(n30418) );
  AND U35707 ( .A(a[33]), .B(b[44]), .Z(n30417) );
  XOR U35708 ( .A(n30423), .B(n30424), .Z(n29966) );
  ANDN U35709 ( .B(n30425), .A(n30426), .Z(n30423) );
  AND U35710 ( .A(a[34]), .B(b[43]), .Z(n30422) );
  XOR U35711 ( .A(n30428), .B(n30429), .Z(n29971) );
  ANDN U35712 ( .B(n30430), .A(n30431), .Z(n30428) );
  AND U35713 ( .A(a[35]), .B(b[42]), .Z(n30427) );
  XOR U35714 ( .A(n30433), .B(n30434), .Z(n29976) );
  ANDN U35715 ( .B(n30435), .A(n30436), .Z(n30433) );
  AND U35716 ( .A(a[36]), .B(b[41]), .Z(n30432) );
  XOR U35717 ( .A(n30438), .B(n30439), .Z(n29981) );
  ANDN U35718 ( .B(n30440), .A(n30441), .Z(n30438) );
  AND U35719 ( .A(a[37]), .B(b[40]), .Z(n30437) );
  XOR U35720 ( .A(n30443), .B(n30444), .Z(n29986) );
  ANDN U35721 ( .B(n30445), .A(n30446), .Z(n30443) );
  AND U35722 ( .A(a[38]), .B(b[39]), .Z(n30442) );
  XOR U35723 ( .A(n30448), .B(n30449), .Z(n29991) );
  ANDN U35724 ( .B(n30450), .A(n30451), .Z(n30448) );
  AND U35725 ( .A(a[39]), .B(b[38]), .Z(n30447) );
  XOR U35726 ( .A(n30453), .B(n30454), .Z(n29996) );
  ANDN U35727 ( .B(n30455), .A(n30456), .Z(n30453) );
  AND U35728 ( .A(a[40]), .B(b[37]), .Z(n30452) );
  XOR U35729 ( .A(n30458), .B(n30459), .Z(n30001) );
  ANDN U35730 ( .B(n30460), .A(n30461), .Z(n30458) );
  AND U35731 ( .A(a[41]), .B(b[36]), .Z(n30457) );
  XOR U35732 ( .A(n30463), .B(n30464), .Z(n30006) );
  ANDN U35733 ( .B(n30465), .A(n30466), .Z(n30463) );
  AND U35734 ( .A(a[42]), .B(b[35]), .Z(n30462) );
  XOR U35735 ( .A(n30468), .B(n30469), .Z(n30011) );
  ANDN U35736 ( .B(n30470), .A(n30471), .Z(n30468) );
  AND U35737 ( .A(a[43]), .B(b[34]), .Z(n30467) );
  XOR U35738 ( .A(n30473), .B(n30474), .Z(n30016) );
  ANDN U35739 ( .B(n30475), .A(n30476), .Z(n30473) );
  AND U35740 ( .A(a[44]), .B(b[33]), .Z(n30472) );
  XOR U35741 ( .A(n30478), .B(n30479), .Z(n30021) );
  ANDN U35742 ( .B(n30480), .A(n30481), .Z(n30478) );
  AND U35743 ( .A(a[45]), .B(b[32]), .Z(n30477) );
  XOR U35744 ( .A(n30483), .B(n30484), .Z(n30026) );
  ANDN U35745 ( .B(n30485), .A(n30486), .Z(n30483) );
  AND U35746 ( .A(a[46]), .B(b[31]), .Z(n30482) );
  XOR U35747 ( .A(n30488), .B(n30489), .Z(n30031) );
  ANDN U35748 ( .B(n30490), .A(n30491), .Z(n30488) );
  AND U35749 ( .A(a[47]), .B(b[30]), .Z(n30487) );
  XOR U35750 ( .A(n30493), .B(n30494), .Z(n30036) );
  ANDN U35751 ( .B(n30495), .A(n30496), .Z(n30493) );
  AND U35752 ( .A(a[48]), .B(b[29]), .Z(n30492) );
  XOR U35753 ( .A(n30498), .B(n30499), .Z(n30041) );
  ANDN U35754 ( .B(n30500), .A(n30501), .Z(n30498) );
  AND U35755 ( .A(a[49]), .B(b[28]), .Z(n30497) );
  XOR U35756 ( .A(n30503), .B(n30504), .Z(n30046) );
  ANDN U35757 ( .B(n30505), .A(n30506), .Z(n30503) );
  AND U35758 ( .A(a[50]), .B(b[27]), .Z(n30502) );
  XOR U35759 ( .A(n30508), .B(n30509), .Z(n30051) );
  ANDN U35760 ( .B(n30510), .A(n30511), .Z(n30508) );
  AND U35761 ( .A(a[51]), .B(b[26]), .Z(n30507) );
  XOR U35762 ( .A(n30513), .B(n30514), .Z(n30056) );
  ANDN U35763 ( .B(n30515), .A(n30516), .Z(n30513) );
  AND U35764 ( .A(a[52]), .B(b[25]), .Z(n30512) );
  XOR U35765 ( .A(n30518), .B(n30519), .Z(n30061) );
  ANDN U35766 ( .B(n30520), .A(n30521), .Z(n30518) );
  AND U35767 ( .A(a[53]), .B(b[24]), .Z(n30517) );
  XOR U35768 ( .A(n30523), .B(n30524), .Z(n30066) );
  ANDN U35769 ( .B(n30525), .A(n30526), .Z(n30523) );
  AND U35770 ( .A(a[54]), .B(b[23]), .Z(n30522) );
  XOR U35771 ( .A(n30528), .B(n30529), .Z(n30071) );
  ANDN U35772 ( .B(n30530), .A(n30531), .Z(n30528) );
  AND U35773 ( .A(a[55]), .B(b[22]), .Z(n30527) );
  XOR U35774 ( .A(n30533), .B(n30534), .Z(n30076) );
  ANDN U35775 ( .B(n30535), .A(n30536), .Z(n30533) );
  AND U35776 ( .A(a[56]), .B(b[21]), .Z(n30532) );
  XOR U35777 ( .A(n30538), .B(n30539), .Z(n30081) );
  ANDN U35778 ( .B(n30540), .A(n30541), .Z(n30538) );
  AND U35779 ( .A(a[57]), .B(b[20]), .Z(n30537) );
  XOR U35780 ( .A(n30543), .B(n30544), .Z(n30086) );
  ANDN U35781 ( .B(n30545), .A(n30546), .Z(n30543) );
  AND U35782 ( .A(a[58]), .B(b[19]), .Z(n30542) );
  XOR U35783 ( .A(n30548), .B(n30549), .Z(n30091) );
  ANDN U35784 ( .B(n30550), .A(n30551), .Z(n30548) );
  AND U35785 ( .A(a[59]), .B(b[18]), .Z(n30547) );
  XOR U35786 ( .A(n30553), .B(n30554), .Z(n30096) );
  ANDN U35787 ( .B(n30555), .A(n30556), .Z(n30553) );
  AND U35788 ( .A(a[60]), .B(b[17]), .Z(n30552) );
  XOR U35789 ( .A(n30558), .B(n30559), .Z(n30101) );
  ANDN U35790 ( .B(n30560), .A(n30561), .Z(n30558) );
  AND U35791 ( .A(a[61]), .B(b[16]), .Z(n30557) );
  XOR U35792 ( .A(n30563), .B(n30564), .Z(n30106) );
  ANDN U35793 ( .B(n30565), .A(n30566), .Z(n30563) );
  AND U35794 ( .A(a[62]), .B(b[15]), .Z(n30562) );
  XOR U35795 ( .A(n30568), .B(n30569), .Z(n30111) );
  ANDN U35796 ( .B(n30570), .A(n30571), .Z(n30568) );
  AND U35797 ( .A(a[63]), .B(b[14]), .Z(n30567) );
  XOR U35798 ( .A(n30573), .B(n30574), .Z(n30116) );
  ANDN U35799 ( .B(n30575), .A(n30576), .Z(n30573) );
  AND U35800 ( .A(a[64]), .B(b[13]), .Z(n30572) );
  XOR U35801 ( .A(n30578), .B(n30579), .Z(n30121) );
  ANDN U35802 ( .B(n30580), .A(n30581), .Z(n30578) );
  AND U35803 ( .A(a[65]), .B(b[12]), .Z(n30577) );
  XOR U35804 ( .A(n30583), .B(n30584), .Z(n30126) );
  ANDN U35805 ( .B(n30585), .A(n30586), .Z(n30583) );
  AND U35806 ( .A(a[66]), .B(b[11]), .Z(n30582) );
  XOR U35807 ( .A(n30588), .B(n30589), .Z(n30131) );
  ANDN U35808 ( .B(n30590), .A(n30591), .Z(n30588) );
  AND U35809 ( .A(a[67]), .B(b[10]), .Z(n30587) );
  XOR U35810 ( .A(n30593), .B(n30594), .Z(n30136) );
  ANDN U35811 ( .B(n30595), .A(n30596), .Z(n30593) );
  AND U35812 ( .A(b[9]), .B(a[68]), .Z(n30592) );
  XOR U35813 ( .A(n30598), .B(n30599), .Z(n30141) );
  ANDN U35814 ( .B(n30600), .A(n30601), .Z(n30598) );
  AND U35815 ( .A(b[8]), .B(a[69]), .Z(n30597) );
  XOR U35816 ( .A(n30603), .B(n30604), .Z(n30146) );
  ANDN U35817 ( .B(n30605), .A(n30606), .Z(n30603) );
  AND U35818 ( .A(b[7]), .B(a[70]), .Z(n30602) );
  XOR U35819 ( .A(n30608), .B(n30609), .Z(n30151) );
  ANDN U35820 ( .B(n30610), .A(n30611), .Z(n30608) );
  AND U35821 ( .A(b[6]), .B(a[71]), .Z(n30607) );
  XOR U35822 ( .A(n30613), .B(n30614), .Z(n30156) );
  ANDN U35823 ( .B(n30615), .A(n30616), .Z(n30613) );
  AND U35824 ( .A(b[5]), .B(a[72]), .Z(n30612) );
  XOR U35825 ( .A(n30618), .B(n30619), .Z(n30161) );
  ANDN U35826 ( .B(n30620), .A(n30621), .Z(n30618) );
  AND U35827 ( .A(b[4]), .B(a[73]), .Z(n30617) );
  XOR U35828 ( .A(n30623), .B(n30624), .Z(n30166) );
  ANDN U35829 ( .B(n30178), .A(n30179), .Z(n30623) );
  AND U35830 ( .A(b[2]), .B(a[74]), .Z(n30625) );
  XNOR U35831 ( .A(n30620), .B(n30624), .Z(n30626) );
  XOR U35832 ( .A(n30627), .B(n30628), .Z(n30624) );
  OR U35833 ( .A(n30181), .B(n30182), .Z(n30628) );
  XNOR U35834 ( .A(n30630), .B(n30631), .Z(n30629) );
  XOR U35835 ( .A(n30630), .B(n30633), .Z(n30181) );
  NAND U35836 ( .A(b[1]), .B(a[74]), .Z(n30633) );
  IV U35837 ( .A(n30627), .Z(n30630) );
  NANDN U35838 ( .A(n57), .B(n58), .Z(n30627) );
  XOR U35839 ( .A(n30634), .B(n30635), .Z(n58) );
  NAND U35840 ( .A(a[74]), .B(b[0]), .Z(n57) );
  XNOR U35841 ( .A(n30615), .B(n30619), .Z(n30636) );
  XNOR U35842 ( .A(n30610), .B(n30614), .Z(n30637) );
  XNOR U35843 ( .A(n30605), .B(n30609), .Z(n30638) );
  XNOR U35844 ( .A(n30600), .B(n30604), .Z(n30639) );
  XNOR U35845 ( .A(n30595), .B(n30599), .Z(n30640) );
  XNOR U35846 ( .A(n30590), .B(n30594), .Z(n30641) );
  XNOR U35847 ( .A(n30585), .B(n30589), .Z(n30642) );
  XNOR U35848 ( .A(n30580), .B(n30584), .Z(n30643) );
  XNOR U35849 ( .A(n30575), .B(n30579), .Z(n30644) );
  XNOR U35850 ( .A(n30570), .B(n30574), .Z(n30645) );
  XNOR U35851 ( .A(n30565), .B(n30569), .Z(n30646) );
  XNOR U35852 ( .A(n30560), .B(n30564), .Z(n30647) );
  XNOR U35853 ( .A(n30555), .B(n30559), .Z(n30648) );
  XNOR U35854 ( .A(n30550), .B(n30554), .Z(n30649) );
  XNOR U35855 ( .A(n30545), .B(n30549), .Z(n30650) );
  XNOR U35856 ( .A(n30540), .B(n30544), .Z(n30651) );
  XNOR U35857 ( .A(n30535), .B(n30539), .Z(n30652) );
  XNOR U35858 ( .A(n30530), .B(n30534), .Z(n30653) );
  XNOR U35859 ( .A(n30525), .B(n30529), .Z(n30654) );
  XNOR U35860 ( .A(n30520), .B(n30524), .Z(n30655) );
  XNOR U35861 ( .A(n30515), .B(n30519), .Z(n30656) );
  XNOR U35862 ( .A(n30510), .B(n30514), .Z(n30657) );
  XNOR U35863 ( .A(n30505), .B(n30509), .Z(n30658) );
  XNOR U35864 ( .A(n30500), .B(n30504), .Z(n30659) );
  XNOR U35865 ( .A(n30495), .B(n30499), .Z(n30660) );
  XNOR U35866 ( .A(n30490), .B(n30494), .Z(n30661) );
  XNOR U35867 ( .A(n30485), .B(n30489), .Z(n30662) );
  XNOR U35868 ( .A(n30480), .B(n30484), .Z(n30663) );
  XNOR U35869 ( .A(n30475), .B(n30479), .Z(n30664) );
  XNOR U35870 ( .A(n30470), .B(n30474), .Z(n30665) );
  XNOR U35871 ( .A(n30465), .B(n30469), .Z(n30666) );
  XNOR U35872 ( .A(n30460), .B(n30464), .Z(n30667) );
  XNOR U35873 ( .A(n30455), .B(n30459), .Z(n30668) );
  XNOR U35874 ( .A(n30450), .B(n30454), .Z(n30669) );
  XNOR U35875 ( .A(n30445), .B(n30449), .Z(n30670) );
  XNOR U35876 ( .A(n30440), .B(n30444), .Z(n30671) );
  XNOR U35877 ( .A(n30435), .B(n30439), .Z(n30672) );
  XNOR U35878 ( .A(n30430), .B(n30434), .Z(n30673) );
  XNOR U35879 ( .A(n30425), .B(n30429), .Z(n30674) );
  XNOR U35880 ( .A(n30420), .B(n30424), .Z(n30675) );
  XNOR U35881 ( .A(n30415), .B(n30419), .Z(n30676) );
  XNOR U35882 ( .A(n30410), .B(n30414), .Z(n30677) );
  XNOR U35883 ( .A(n30405), .B(n30409), .Z(n30678) );
  XNOR U35884 ( .A(n30400), .B(n30404), .Z(n30679) );
  XNOR U35885 ( .A(n30395), .B(n30399), .Z(n30680) );
  XNOR U35886 ( .A(n30390), .B(n30394), .Z(n30681) );
  XNOR U35887 ( .A(n30385), .B(n30389), .Z(n30682) );
  XNOR U35888 ( .A(n30380), .B(n30384), .Z(n30683) );
  XNOR U35889 ( .A(n30375), .B(n30379), .Z(n30684) );
  XNOR U35890 ( .A(n30370), .B(n30374), .Z(n30685) );
  XNOR U35891 ( .A(n30365), .B(n30369), .Z(n30686) );
  XNOR U35892 ( .A(n30360), .B(n30364), .Z(n30687) );
  XNOR U35893 ( .A(n30355), .B(n30359), .Z(n30688) );
  XNOR U35894 ( .A(n30350), .B(n30354), .Z(n30689) );
  XNOR U35895 ( .A(n30345), .B(n30349), .Z(n30690) );
  XNOR U35896 ( .A(n30340), .B(n30344), .Z(n30691) );
  XNOR U35897 ( .A(n30335), .B(n30339), .Z(n30692) );
  XNOR U35898 ( .A(n30330), .B(n30334), .Z(n30693) );
  XNOR U35899 ( .A(n30325), .B(n30329), .Z(n30694) );
  XNOR U35900 ( .A(n30320), .B(n30324), .Z(n30695) );
  XNOR U35901 ( .A(n30315), .B(n30319), .Z(n30696) );
  XNOR U35902 ( .A(n30310), .B(n30314), .Z(n30697) );
  XNOR U35903 ( .A(n30305), .B(n30309), .Z(n30698) );
  XNOR U35904 ( .A(n30300), .B(n30304), .Z(n30699) );
  XNOR U35905 ( .A(n30295), .B(n30299), .Z(n30700) );
  XNOR U35906 ( .A(n30290), .B(n30294), .Z(n30701) );
  XNOR U35907 ( .A(n30285), .B(n30289), .Z(n30702) );
  XNOR U35908 ( .A(n30280), .B(n30284), .Z(n30703) );
  XNOR U35909 ( .A(n30275), .B(n30279), .Z(n30704) );
  XNOR U35910 ( .A(n30270), .B(n30274), .Z(n30705) );
  XNOR U35911 ( .A(n30265), .B(n30269), .Z(n30706) );
  XNOR U35912 ( .A(n30260), .B(n30264), .Z(n30707) );
  XOR U35913 ( .A(n30708), .B(n30259), .Z(n30260) );
  AND U35914 ( .A(a[0]), .B(b[76]), .Z(n30708) );
  XNOR U35915 ( .A(n30709), .B(n30259), .Z(n30261) );
  XNOR U35916 ( .A(n30710), .B(n30711), .Z(n30259) );
  ANDN U35917 ( .B(n30712), .A(n30713), .Z(n30710) );
  AND U35918 ( .A(a[1]), .B(b[75]), .Z(n30709) );
  XOR U35919 ( .A(n30715), .B(n30716), .Z(n30264) );
  ANDN U35920 ( .B(n30717), .A(n30718), .Z(n30715) );
  AND U35921 ( .A(a[2]), .B(b[74]), .Z(n30714) );
  XOR U35922 ( .A(n30720), .B(n30721), .Z(n30269) );
  ANDN U35923 ( .B(n30722), .A(n30723), .Z(n30720) );
  AND U35924 ( .A(a[3]), .B(b[73]), .Z(n30719) );
  XOR U35925 ( .A(n30725), .B(n30726), .Z(n30274) );
  ANDN U35926 ( .B(n30727), .A(n30728), .Z(n30725) );
  AND U35927 ( .A(a[4]), .B(b[72]), .Z(n30724) );
  XOR U35928 ( .A(n30730), .B(n30731), .Z(n30279) );
  ANDN U35929 ( .B(n30732), .A(n30733), .Z(n30730) );
  AND U35930 ( .A(a[5]), .B(b[71]), .Z(n30729) );
  XOR U35931 ( .A(n30735), .B(n30736), .Z(n30284) );
  ANDN U35932 ( .B(n30737), .A(n30738), .Z(n30735) );
  AND U35933 ( .A(a[6]), .B(b[70]), .Z(n30734) );
  XOR U35934 ( .A(n30740), .B(n30741), .Z(n30289) );
  ANDN U35935 ( .B(n30742), .A(n30743), .Z(n30740) );
  AND U35936 ( .A(a[7]), .B(b[69]), .Z(n30739) );
  XOR U35937 ( .A(n30745), .B(n30746), .Z(n30294) );
  ANDN U35938 ( .B(n30747), .A(n30748), .Z(n30745) );
  AND U35939 ( .A(a[8]), .B(b[68]), .Z(n30744) );
  XOR U35940 ( .A(n30750), .B(n30751), .Z(n30299) );
  ANDN U35941 ( .B(n30752), .A(n30753), .Z(n30750) );
  AND U35942 ( .A(a[9]), .B(b[67]), .Z(n30749) );
  XOR U35943 ( .A(n30755), .B(n30756), .Z(n30304) );
  ANDN U35944 ( .B(n30757), .A(n30758), .Z(n30755) );
  AND U35945 ( .A(a[10]), .B(b[66]), .Z(n30754) );
  XOR U35946 ( .A(n30760), .B(n30761), .Z(n30309) );
  ANDN U35947 ( .B(n30762), .A(n30763), .Z(n30760) );
  AND U35948 ( .A(a[11]), .B(b[65]), .Z(n30759) );
  XOR U35949 ( .A(n30765), .B(n30766), .Z(n30314) );
  ANDN U35950 ( .B(n30767), .A(n30768), .Z(n30765) );
  AND U35951 ( .A(a[12]), .B(b[64]), .Z(n30764) );
  XOR U35952 ( .A(n30770), .B(n30771), .Z(n30319) );
  ANDN U35953 ( .B(n30772), .A(n30773), .Z(n30770) );
  AND U35954 ( .A(a[13]), .B(b[63]), .Z(n30769) );
  XOR U35955 ( .A(n30775), .B(n30776), .Z(n30324) );
  ANDN U35956 ( .B(n30777), .A(n30778), .Z(n30775) );
  AND U35957 ( .A(a[14]), .B(b[62]), .Z(n30774) );
  XOR U35958 ( .A(n30780), .B(n30781), .Z(n30329) );
  ANDN U35959 ( .B(n30782), .A(n30783), .Z(n30780) );
  AND U35960 ( .A(a[15]), .B(b[61]), .Z(n30779) );
  XOR U35961 ( .A(n30785), .B(n30786), .Z(n30334) );
  ANDN U35962 ( .B(n30787), .A(n30788), .Z(n30785) );
  AND U35963 ( .A(a[16]), .B(b[60]), .Z(n30784) );
  XOR U35964 ( .A(n30790), .B(n30791), .Z(n30339) );
  ANDN U35965 ( .B(n30792), .A(n30793), .Z(n30790) );
  AND U35966 ( .A(a[17]), .B(b[59]), .Z(n30789) );
  XOR U35967 ( .A(n30795), .B(n30796), .Z(n30344) );
  ANDN U35968 ( .B(n30797), .A(n30798), .Z(n30795) );
  AND U35969 ( .A(a[18]), .B(b[58]), .Z(n30794) );
  XOR U35970 ( .A(n30800), .B(n30801), .Z(n30349) );
  ANDN U35971 ( .B(n30802), .A(n30803), .Z(n30800) );
  AND U35972 ( .A(a[19]), .B(b[57]), .Z(n30799) );
  XOR U35973 ( .A(n30805), .B(n30806), .Z(n30354) );
  ANDN U35974 ( .B(n30807), .A(n30808), .Z(n30805) );
  AND U35975 ( .A(a[20]), .B(b[56]), .Z(n30804) );
  XOR U35976 ( .A(n30810), .B(n30811), .Z(n30359) );
  ANDN U35977 ( .B(n30812), .A(n30813), .Z(n30810) );
  AND U35978 ( .A(a[21]), .B(b[55]), .Z(n30809) );
  XOR U35979 ( .A(n30815), .B(n30816), .Z(n30364) );
  ANDN U35980 ( .B(n30817), .A(n30818), .Z(n30815) );
  AND U35981 ( .A(a[22]), .B(b[54]), .Z(n30814) );
  XOR U35982 ( .A(n30820), .B(n30821), .Z(n30369) );
  ANDN U35983 ( .B(n30822), .A(n30823), .Z(n30820) );
  AND U35984 ( .A(a[23]), .B(b[53]), .Z(n30819) );
  XOR U35985 ( .A(n30825), .B(n30826), .Z(n30374) );
  ANDN U35986 ( .B(n30827), .A(n30828), .Z(n30825) );
  AND U35987 ( .A(a[24]), .B(b[52]), .Z(n30824) );
  XOR U35988 ( .A(n30830), .B(n30831), .Z(n30379) );
  ANDN U35989 ( .B(n30832), .A(n30833), .Z(n30830) );
  AND U35990 ( .A(a[25]), .B(b[51]), .Z(n30829) );
  XOR U35991 ( .A(n30835), .B(n30836), .Z(n30384) );
  ANDN U35992 ( .B(n30837), .A(n30838), .Z(n30835) );
  AND U35993 ( .A(a[26]), .B(b[50]), .Z(n30834) );
  XOR U35994 ( .A(n30840), .B(n30841), .Z(n30389) );
  ANDN U35995 ( .B(n30842), .A(n30843), .Z(n30840) );
  AND U35996 ( .A(a[27]), .B(b[49]), .Z(n30839) );
  XOR U35997 ( .A(n30845), .B(n30846), .Z(n30394) );
  ANDN U35998 ( .B(n30847), .A(n30848), .Z(n30845) );
  AND U35999 ( .A(a[28]), .B(b[48]), .Z(n30844) );
  XOR U36000 ( .A(n30850), .B(n30851), .Z(n30399) );
  ANDN U36001 ( .B(n30852), .A(n30853), .Z(n30850) );
  AND U36002 ( .A(a[29]), .B(b[47]), .Z(n30849) );
  XOR U36003 ( .A(n30855), .B(n30856), .Z(n30404) );
  ANDN U36004 ( .B(n30857), .A(n30858), .Z(n30855) );
  AND U36005 ( .A(a[30]), .B(b[46]), .Z(n30854) );
  XOR U36006 ( .A(n30860), .B(n30861), .Z(n30409) );
  ANDN U36007 ( .B(n30862), .A(n30863), .Z(n30860) );
  AND U36008 ( .A(a[31]), .B(b[45]), .Z(n30859) );
  XOR U36009 ( .A(n30865), .B(n30866), .Z(n30414) );
  ANDN U36010 ( .B(n30867), .A(n30868), .Z(n30865) );
  AND U36011 ( .A(a[32]), .B(b[44]), .Z(n30864) );
  XOR U36012 ( .A(n30870), .B(n30871), .Z(n30419) );
  ANDN U36013 ( .B(n30872), .A(n30873), .Z(n30870) );
  AND U36014 ( .A(a[33]), .B(b[43]), .Z(n30869) );
  XOR U36015 ( .A(n30875), .B(n30876), .Z(n30424) );
  ANDN U36016 ( .B(n30877), .A(n30878), .Z(n30875) );
  AND U36017 ( .A(a[34]), .B(b[42]), .Z(n30874) );
  XOR U36018 ( .A(n30880), .B(n30881), .Z(n30429) );
  ANDN U36019 ( .B(n30882), .A(n30883), .Z(n30880) );
  AND U36020 ( .A(a[35]), .B(b[41]), .Z(n30879) );
  XOR U36021 ( .A(n30885), .B(n30886), .Z(n30434) );
  ANDN U36022 ( .B(n30887), .A(n30888), .Z(n30885) );
  AND U36023 ( .A(a[36]), .B(b[40]), .Z(n30884) );
  XOR U36024 ( .A(n30890), .B(n30891), .Z(n30439) );
  ANDN U36025 ( .B(n30892), .A(n30893), .Z(n30890) );
  AND U36026 ( .A(a[37]), .B(b[39]), .Z(n30889) );
  XOR U36027 ( .A(n30895), .B(n30896), .Z(n30444) );
  ANDN U36028 ( .B(n30897), .A(n30898), .Z(n30895) );
  AND U36029 ( .A(a[38]), .B(b[38]), .Z(n30894) );
  XOR U36030 ( .A(n30900), .B(n30901), .Z(n30449) );
  ANDN U36031 ( .B(n30902), .A(n30903), .Z(n30900) );
  AND U36032 ( .A(a[39]), .B(b[37]), .Z(n30899) );
  XOR U36033 ( .A(n30905), .B(n30906), .Z(n30454) );
  ANDN U36034 ( .B(n30907), .A(n30908), .Z(n30905) );
  AND U36035 ( .A(a[40]), .B(b[36]), .Z(n30904) );
  XOR U36036 ( .A(n30910), .B(n30911), .Z(n30459) );
  ANDN U36037 ( .B(n30912), .A(n30913), .Z(n30910) );
  AND U36038 ( .A(a[41]), .B(b[35]), .Z(n30909) );
  XOR U36039 ( .A(n30915), .B(n30916), .Z(n30464) );
  ANDN U36040 ( .B(n30917), .A(n30918), .Z(n30915) );
  AND U36041 ( .A(a[42]), .B(b[34]), .Z(n30914) );
  XOR U36042 ( .A(n30920), .B(n30921), .Z(n30469) );
  ANDN U36043 ( .B(n30922), .A(n30923), .Z(n30920) );
  AND U36044 ( .A(a[43]), .B(b[33]), .Z(n30919) );
  XOR U36045 ( .A(n30925), .B(n30926), .Z(n30474) );
  ANDN U36046 ( .B(n30927), .A(n30928), .Z(n30925) );
  AND U36047 ( .A(a[44]), .B(b[32]), .Z(n30924) );
  XOR U36048 ( .A(n30930), .B(n30931), .Z(n30479) );
  ANDN U36049 ( .B(n30932), .A(n30933), .Z(n30930) );
  AND U36050 ( .A(a[45]), .B(b[31]), .Z(n30929) );
  XOR U36051 ( .A(n30935), .B(n30936), .Z(n30484) );
  ANDN U36052 ( .B(n30937), .A(n30938), .Z(n30935) );
  AND U36053 ( .A(a[46]), .B(b[30]), .Z(n30934) );
  XOR U36054 ( .A(n30940), .B(n30941), .Z(n30489) );
  ANDN U36055 ( .B(n30942), .A(n30943), .Z(n30940) );
  AND U36056 ( .A(a[47]), .B(b[29]), .Z(n30939) );
  XOR U36057 ( .A(n30945), .B(n30946), .Z(n30494) );
  ANDN U36058 ( .B(n30947), .A(n30948), .Z(n30945) );
  AND U36059 ( .A(a[48]), .B(b[28]), .Z(n30944) );
  XOR U36060 ( .A(n30950), .B(n30951), .Z(n30499) );
  ANDN U36061 ( .B(n30952), .A(n30953), .Z(n30950) );
  AND U36062 ( .A(a[49]), .B(b[27]), .Z(n30949) );
  XOR U36063 ( .A(n30955), .B(n30956), .Z(n30504) );
  ANDN U36064 ( .B(n30957), .A(n30958), .Z(n30955) );
  AND U36065 ( .A(a[50]), .B(b[26]), .Z(n30954) );
  XOR U36066 ( .A(n30960), .B(n30961), .Z(n30509) );
  ANDN U36067 ( .B(n30962), .A(n30963), .Z(n30960) );
  AND U36068 ( .A(a[51]), .B(b[25]), .Z(n30959) );
  XOR U36069 ( .A(n30965), .B(n30966), .Z(n30514) );
  ANDN U36070 ( .B(n30967), .A(n30968), .Z(n30965) );
  AND U36071 ( .A(a[52]), .B(b[24]), .Z(n30964) );
  XOR U36072 ( .A(n30970), .B(n30971), .Z(n30519) );
  ANDN U36073 ( .B(n30972), .A(n30973), .Z(n30970) );
  AND U36074 ( .A(a[53]), .B(b[23]), .Z(n30969) );
  XOR U36075 ( .A(n30975), .B(n30976), .Z(n30524) );
  ANDN U36076 ( .B(n30977), .A(n30978), .Z(n30975) );
  AND U36077 ( .A(a[54]), .B(b[22]), .Z(n30974) );
  XOR U36078 ( .A(n30980), .B(n30981), .Z(n30529) );
  ANDN U36079 ( .B(n30982), .A(n30983), .Z(n30980) );
  AND U36080 ( .A(a[55]), .B(b[21]), .Z(n30979) );
  XOR U36081 ( .A(n30985), .B(n30986), .Z(n30534) );
  ANDN U36082 ( .B(n30987), .A(n30988), .Z(n30985) );
  AND U36083 ( .A(a[56]), .B(b[20]), .Z(n30984) );
  XOR U36084 ( .A(n30990), .B(n30991), .Z(n30539) );
  ANDN U36085 ( .B(n30992), .A(n30993), .Z(n30990) );
  AND U36086 ( .A(a[57]), .B(b[19]), .Z(n30989) );
  XOR U36087 ( .A(n30995), .B(n30996), .Z(n30544) );
  ANDN U36088 ( .B(n30997), .A(n30998), .Z(n30995) );
  AND U36089 ( .A(a[58]), .B(b[18]), .Z(n30994) );
  XOR U36090 ( .A(n31000), .B(n31001), .Z(n30549) );
  ANDN U36091 ( .B(n31002), .A(n31003), .Z(n31000) );
  AND U36092 ( .A(a[59]), .B(b[17]), .Z(n30999) );
  XOR U36093 ( .A(n31005), .B(n31006), .Z(n30554) );
  ANDN U36094 ( .B(n31007), .A(n31008), .Z(n31005) );
  AND U36095 ( .A(a[60]), .B(b[16]), .Z(n31004) );
  XOR U36096 ( .A(n31010), .B(n31011), .Z(n30559) );
  ANDN U36097 ( .B(n31012), .A(n31013), .Z(n31010) );
  AND U36098 ( .A(a[61]), .B(b[15]), .Z(n31009) );
  XOR U36099 ( .A(n31015), .B(n31016), .Z(n30564) );
  ANDN U36100 ( .B(n31017), .A(n31018), .Z(n31015) );
  AND U36101 ( .A(a[62]), .B(b[14]), .Z(n31014) );
  XOR U36102 ( .A(n31020), .B(n31021), .Z(n30569) );
  ANDN U36103 ( .B(n31022), .A(n31023), .Z(n31020) );
  AND U36104 ( .A(a[63]), .B(b[13]), .Z(n31019) );
  XOR U36105 ( .A(n31025), .B(n31026), .Z(n30574) );
  ANDN U36106 ( .B(n31027), .A(n31028), .Z(n31025) );
  AND U36107 ( .A(a[64]), .B(b[12]), .Z(n31024) );
  XOR U36108 ( .A(n31030), .B(n31031), .Z(n30579) );
  ANDN U36109 ( .B(n31032), .A(n31033), .Z(n31030) );
  AND U36110 ( .A(a[65]), .B(b[11]), .Z(n31029) );
  XOR U36111 ( .A(n31035), .B(n31036), .Z(n30584) );
  ANDN U36112 ( .B(n31037), .A(n31038), .Z(n31035) );
  AND U36113 ( .A(a[66]), .B(b[10]), .Z(n31034) );
  XOR U36114 ( .A(n31040), .B(n31041), .Z(n30589) );
  ANDN U36115 ( .B(n31042), .A(n31043), .Z(n31040) );
  AND U36116 ( .A(b[9]), .B(a[67]), .Z(n31039) );
  XOR U36117 ( .A(n31045), .B(n31046), .Z(n30594) );
  ANDN U36118 ( .B(n31047), .A(n31048), .Z(n31045) );
  AND U36119 ( .A(b[8]), .B(a[68]), .Z(n31044) );
  XOR U36120 ( .A(n31050), .B(n31051), .Z(n30599) );
  ANDN U36121 ( .B(n31052), .A(n31053), .Z(n31050) );
  AND U36122 ( .A(b[7]), .B(a[69]), .Z(n31049) );
  XOR U36123 ( .A(n31055), .B(n31056), .Z(n30604) );
  ANDN U36124 ( .B(n31057), .A(n31058), .Z(n31055) );
  AND U36125 ( .A(b[6]), .B(a[70]), .Z(n31054) );
  XOR U36126 ( .A(n31060), .B(n31061), .Z(n30609) );
  ANDN U36127 ( .B(n31062), .A(n31063), .Z(n31060) );
  AND U36128 ( .A(b[5]), .B(a[71]), .Z(n31059) );
  XOR U36129 ( .A(n31065), .B(n31066), .Z(n30614) );
  ANDN U36130 ( .B(n31067), .A(n31068), .Z(n31065) );
  AND U36131 ( .A(b[4]), .B(a[72]), .Z(n31064) );
  XOR U36132 ( .A(n31070), .B(n31071), .Z(n30619) );
  ANDN U36133 ( .B(n30631), .A(n30632), .Z(n31070) );
  AND U36134 ( .A(b[2]), .B(a[73]), .Z(n31072) );
  XNOR U36135 ( .A(n31067), .B(n31071), .Z(n31073) );
  XOR U36136 ( .A(n31074), .B(n31075), .Z(n31071) );
  OR U36137 ( .A(n30634), .B(n30635), .Z(n31075) );
  XNOR U36138 ( .A(n31077), .B(n31078), .Z(n31076) );
  XOR U36139 ( .A(n31077), .B(n31080), .Z(n30634) );
  NAND U36140 ( .A(b[1]), .B(a[73]), .Z(n31080) );
  IV U36141 ( .A(n31074), .Z(n31077) );
  NANDN U36142 ( .A(n59), .B(n60), .Z(n31074) );
  XOR U36143 ( .A(n31081), .B(n31082), .Z(n60) );
  NAND U36144 ( .A(a[73]), .B(b[0]), .Z(n59) );
  XNOR U36145 ( .A(n31062), .B(n31066), .Z(n31083) );
  XNOR U36146 ( .A(n31057), .B(n31061), .Z(n31084) );
  XNOR U36147 ( .A(n31052), .B(n31056), .Z(n31085) );
  XNOR U36148 ( .A(n31047), .B(n31051), .Z(n31086) );
  XNOR U36149 ( .A(n31042), .B(n31046), .Z(n31087) );
  XNOR U36150 ( .A(n31037), .B(n31041), .Z(n31088) );
  XNOR U36151 ( .A(n31032), .B(n31036), .Z(n31089) );
  XNOR U36152 ( .A(n31027), .B(n31031), .Z(n31090) );
  XNOR U36153 ( .A(n31022), .B(n31026), .Z(n31091) );
  XNOR U36154 ( .A(n31017), .B(n31021), .Z(n31092) );
  XNOR U36155 ( .A(n31012), .B(n31016), .Z(n31093) );
  XNOR U36156 ( .A(n31007), .B(n31011), .Z(n31094) );
  XNOR U36157 ( .A(n31002), .B(n31006), .Z(n31095) );
  XNOR U36158 ( .A(n30997), .B(n31001), .Z(n31096) );
  XNOR U36159 ( .A(n30992), .B(n30996), .Z(n31097) );
  XNOR U36160 ( .A(n30987), .B(n30991), .Z(n31098) );
  XNOR U36161 ( .A(n30982), .B(n30986), .Z(n31099) );
  XNOR U36162 ( .A(n30977), .B(n30981), .Z(n31100) );
  XNOR U36163 ( .A(n30972), .B(n30976), .Z(n31101) );
  XNOR U36164 ( .A(n30967), .B(n30971), .Z(n31102) );
  XNOR U36165 ( .A(n30962), .B(n30966), .Z(n31103) );
  XNOR U36166 ( .A(n30957), .B(n30961), .Z(n31104) );
  XNOR U36167 ( .A(n30952), .B(n30956), .Z(n31105) );
  XNOR U36168 ( .A(n30947), .B(n30951), .Z(n31106) );
  XNOR U36169 ( .A(n30942), .B(n30946), .Z(n31107) );
  XNOR U36170 ( .A(n30937), .B(n30941), .Z(n31108) );
  XNOR U36171 ( .A(n30932), .B(n30936), .Z(n31109) );
  XNOR U36172 ( .A(n30927), .B(n30931), .Z(n31110) );
  XNOR U36173 ( .A(n30922), .B(n30926), .Z(n31111) );
  XNOR U36174 ( .A(n30917), .B(n30921), .Z(n31112) );
  XNOR U36175 ( .A(n30912), .B(n30916), .Z(n31113) );
  XNOR U36176 ( .A(n30907), .B(n30911), .Z(n31114) );
  XNOR U36177 ( .A(n30902), .B(n30906), .Z(n31115) );
  XNOR U36178 ( .A(n30897), .B(n30901), .Z(n31116) );
  XNOR U36179 ( .A(n30892), .B(n30896), .Z(n31117) );
  XNOR U36180 ( .A(n30887), .B(n30891), .Z(n31118) );
  XNOR U36181 ( .A(n30882), .B(n30886), .Z(n31119) );
  XNOR U36182 ( .A(n30877), .B(n30881), .Z(n31120) );
  XNOR U36183 ( .A(n30872), .B(n30876), .Z(n31121) );
  XNOR U36184 ( .A(n30867), .B(n30871), .Z(n31122) );
  XNOR U36185 ( .A(n30862), .B(n30866), .Z(n31123) );
  XNOR U36186 ( .A(n30857), .B(n30861), .Z(n31124) );
  XNOR U36187 ( .A(n30852), .B(n30856), .Z(n31125) );
  XNOR U36188 ( .A(n30847), .B(n30851), .Z(n31126) );
  XNOR U36189 ( .A(n30842), .B(n30846), .Z(n31127) );
  XNOR U36190 ( .A(n30837), .B(n30841), .Z(n31128) );
  XNOR U36191 ( .A(n30832), .B(n30836), .Z(n31129) );
  XNOR U36192 ( .A(n30827), .B(n30831), .Z(n31130) );
  XNOR U36193 ( .A(n30822), .B(n30826), .Z(n31131) );
  XNOR U36194 ( .A(n30817), .B(n30821), .Z(n31132) );
  XNOR U36195 ( .A(n30812), .B(n30816), .Z(n31133) );
  XNOR U36196 ( .A(n30807), .B(n30811), .Z(n31134) );
  XNOR U36197 ( .A(n30802), .B(n30806), .Z(n31135) );
  XNOR U36198 ( .A(n30797), .B(n30801), .Z(n31136) );
  XNOR U36199 ( .A(n30792), .B(n30796), .Z(n31137) );
  XNOR U36200 ( .A(n30787), .B(n30791), .Z(n31138) );
  XNOR U36201 ( .A(n30782), .B(n30786), .Z(n31139) );
  XNOR U36202 ( .A(n30777), .B(n30781), .Z(n31140) );
  XNOR U36203 ( .A(n30772), .B(n30776), .Z(n31141) );
  XNOR U36204 ( .A(n30767), .B(n30771), .Z(n31142) );
  XNOR U36205 ( .A(n30762), .B(n30766), .Z(n31143) );
  XNOR U36206 ( .A(n30757), .B(n30761), .Z(n31144) );
  XNOR U36207 ( .A(n30752), .B(n30756), .Z(n31145) );
  XNOR U36208 ( .A(n30747), .B(n30751), .Z(n31146) );
  XNOR U36209 ( .A(n30742), .B(n30746), .Z(n31147) );
  XNOR U36210 ( .A(n30737), .B(n30741), .Z(n31148) );
  XNOR U36211 ( .A(n30732), .B(n30736), .Z(n31149) );
  XNOR U36212 ( .A(n30727), .B(n30731), .Z(n31150) );
  XNOR U36213 ( .A(n30722), .B(n30726), .Z(n31151) );
  XNOR U36214 ( .A(n30717), .B(n30721), .Z(n31152) );
  XNOR U36215 ( .A(n30712), .B(n30716), .Z(n31153) );
  XNOR U36216 ( .A(n31154), .B(n30711), .Z(n30712) );
  AND U36217 ( .A(a[0]), .B(b[75]), .Z(n31154) );
  XOR U36218 ( .A(n31155), .B(n30711), .Z(n30713) );
  XNOR U36219 ( .A(n31156), .B(n31157), .Z(n30711) );
  ANDN U36220 ( .B(n31158), .A(n31159), .Z(n31156) );
  AND U36221 ( .A(a[1]), .B(b[74]), .Z(n31155) );
  XOR U36222 ( .A(n31161), .B(n31162), .Z(n30716) );
  ANDN U36223 ( .B(n31163), .A(n31164), .Z(n31161) );
  AND U36224 ( .A(a[2]), .B(b[73]), .Z(n31160) );
  XOR U36225 ( .A(n31166), .B(n31167), .Z(n30721) );
  ANDN U36226 ( .B(n31168), .A(n31169), .Z(n31166) );
  AND U36227 ( .A(a[3]), .B(b[72]), .Z(n31165) );
  XOR U36228 ( .A(n31171), .B(n31172), .Z(n30726) );
  ANDN U36229 ( .B(n31173), .A(n31174), .Z(n31171) );
  AND U36230 ( .A(a[4]), .B(b[71]), .Z(n31170) );
  XOR U36231 ( .A(n31176), .B(n31177), .Z(n30731) );
  ANDN U36232 ( .B(n31178), .A(n31179), .Z(n31176) );
  AND U36233 ( .A(a[5]), .B(b[70]), .Z(n31175) );
  XOR U36234 ( .A(n31181), .B(n31182), .Z(n30736) );
  ANDN U36235 ( .B(n31183), .A(n31184), .Z(n31181) );
  AND U36236 ( .A(a[6]), .B(b[69]), .Z(n31180) );
  XOR U36237 ( .A(n31186), .B(n31187), .Z(n30741) );
  ANDN U36238 ( .B(n31188), .A(n31189), .Z(n31186) );
  AND U36239 ( .A(a[7]), .B(b[68]), .Z(n31185) );
  XOR U36240 ( .A(n31191), .B(n31192), .Z(n30746) );
  ANDN U36241 ( .B(n31193), .A(n31194), .Z(n31191) );
  AND U36242 ( .A(a[8]), .B(b[67]), .Z(n31190) );
  XOR U36243 ( .A(n31196), .B(n31197), .Z(n30751) );
  ANDN U36244 ( .B(n31198), .A(n31199), .Z(n31196) );
  AND U36245 ( .A(a[9]), .B(b[66]), .Z(n31195) );
  XOR U36246 ( .A(n31201), .B(n31202), .Z(n30756) );
  ANDN U36247 ( .B(n31203), .A(n31204), .Z(n31201) );
  AND U36248 ( .A(a[10]), .B(b[65]), .Z(n31200) );
  XOR U36249 ( .A(n31206), .B(n31207), .Z(n30761) );
  ANDN U36250 ( .B(n31208), .A(n31209), .Z(n31206) );
  AND U36251 ( .A(a[11]), .B(b[64]), .Z(n31205) );
  XOR U36252 ( .A(n31211), .B(n31212), .Z(n30766) );
  ANDN U36253 ( .B(n31213), .A(n31214), .Z(n31211) );
  AND U36254 ( .A(a[12]), .B(b[63]), .Z(n31210) );
  XOR U36255 ( .A(n31216), .B(n31217), .Z(n30771) );
  ANDN U36256 ( .B(n31218), .A(n31219), .Z(n31216) );
  AND U36257 ( .A(a[13]), .B(b[62]), .Z(n31215) );
  XOR U36258 ( .A(n31221), .B(n31222), .Z(n30776) );
  ANDN U36259 ( .B(n31223), .A(n31224), .Z(n31221) );
  AND U36260 ( .A(a[14]), .B(b[61]), .Z(n31220) );
  XOR U36261 ( .A(n31226), .B(n31227), .Z(n30781) );
  ANDN U36262 ( .B(n31228), .A(n31229), .Z(n31226) );
  AND U36263 ( .A(a[15]), .B(b[60]), .Z(n31225) );
  XOR U36264 ( .A(n31231), .B(n31232), .Z(n30786) );
  ANDN U36265 ( .B(n31233), .A(n31234), .Z(n31231) );
  AND U36266 ( .A(a[16]), .B(b[59]), .Z(n31230) );
  XOR U36267 ( .A(n31236), .B(n31237), .Z(n30791) );
  ANDN U36268 ( .B(n31238), .A(n31239), .Z(n31236) );
  AND U36269 ( .A(a[17]), .B(b[58]), .Z(n31235) );
  XOR U36270 ( .A(n31241), .B(n31242), .Z(n30796) );
  ANDN U36271 ( .B(n31243), .A(n31244), .Z(n31241) );
  AND U36272 ( .A(a[18]), .B(b[57]), .Z(n31240) );
  XOR U36273 ( .A(n31246), .B(n31247), .Z(n30801) );
  ANDN U36274 ( .B(n31248), .A(n31249), .Z(n31246) );
  AND U36275 ( .A(a[19]), .B(b[56]), .Z(n31245) );
  XOR U36276 ( .A(n31251), .B(n31252), .Z(n30806) );
  ANDN U36277 ( .B(n31253), .A(n31254), .Z(n31251) );
  AND U36278 ( .A(a[20]), .B(b[55]), .Z(n31250) );
  XOR U36279 ( .A(n31256), .B(n31257), .Z(n30811) );
  ANDN U36280 ( .B(n31258), .A(n31259), .Z(n31256) );
  AND U36281 ( .A(a[21]), .B(b[54]), .Z(n31255) );
  XOR U36282 ( .A(n31261), .B(n31262), .Z(n30816) );
  ANDN U36283 ( .B(n31263), .A(n31264), .Z(n31261) );
  AND U36284 ( .A(a[22]), .B(b[53]), .Z(n31260) );
  XOR U36285 ( .A(n31266), .B(n31267), .Z(n30821) );
  ANDN U36286 ( .B(n31268), .A(n31269), .Z(n31266) );
  AND U36287 ( .A(a[23]), .B(b[52]), .Z(n31265) );
  XOR U36288 ( .A(n31271), .B(n31272), .Z(n30826) );
  ANDN U36289 ( .B(n31273), .A(n31274), .Z(n31271) );
  AND U36290 ( .A(a[24]), .B(b[51]), .Z(n31270) );
  XOR U36291 ( .A(n31276), .B(n31277), .Z(n30831) );
  ANDN U36292 ( .B(n31278), .A(n31279), .Z(n31276) );
  AND U36293 ( .A(a[25]), .B(b[50]), .Z(n31275) );
  XOR U36294 ( .A(n31281), .B(n31282), .Z(n30836) );
  ANDN U36295 ( .B(n31283), .A(n31284), .Z(n31281) );
  AND U36296 ( .A(a[26]), .B(b[49]), .Z(n31280) );
  XOR U36297 ( .A(n31286), .B(n31287), .Z(n30841) );
  ANDN U36298 ( .B(n31288), .A(n31289), .Z(n31286) );
  AND U36299 ( .A(a[27]), .B(b[48]), .Z(n31285) );
  XOR U36300 ( .A(n31291), .B(n31292), .Z(n30846) );
  ANDN U36301 ( .B(n31293), .A(n31294), .Z(n31291) );
  AND U36302 ( .A(a[28]), .B(b[47]), .Z(n31290) );
  XOR U36303 ( .A(n31296), .B(n31297), .Z(n30851) );
  ANDN U36304 ( .B(n31298), .A(n31299), .Z(n31296) );
  AND U36305 ( .A(a[29]), .B(b[46]), .Z(n31295) );
  XOR U36306 ( .A(n31301), .B(n31302), .Z(n30856) );
  ANDN U36307 ( .B(n31303), .A(n31304), .Z(n31301) );
  AND U36308 ( .A(a[30]), .B(b[45]), .Z(n31300) );
  XOR U36309 ( .A(n31306), .B(n31307), .Z(n30861) );
  ANDN U36310 ( .B(n31308), .A(n31309), .Z(n31306) );
  AND U36311 ( .A(a[31]), .B(b[44]), .Z(n31305) );
  XOR U36312 ( .A(n31311), .B(n31312), .Z(n30866) );
  ANDN U36313 ( .B(n31313), .A(n31314), .Z(n31311) );
  AND U36314 ( .A(a[32]), .B(b[43]), .Z(n31310) );
  XOR U36315 ( .A(n31316), .B(n31317), .Z(n30871) );
  ANDN U36316 ( .B(n31318), .A(n31319), .Z(n31316) );
  AND U36317 ( .A(a[33]), .B(b[42]), .Z(n31315) );
  XOR U36318 ( .A(n31321), .B(n31322), .Z(n30876) );
  ANDN U36319 ( .B(n31323), .A(n31324), .Z(n31321) );
  AND U36320 ( .A(a[34]), .B(b[41]), .Z(n31320) );
  XOR U36321 ( .A(n31326), .B(n31327), .Z(n30881) );
  ANDN U36322 ( .B(n31328), .A(n31329), .Z(n31326) );
  AND U36323 ( .A(a[35]), .B(b[40]), .Z(n31325) );
  XOR U36324 ( .A(n31331), .B(n31332), .Z(n30886) );
  ANDN U36325 ( .B(n31333), .A(n31334), .Z(n31331) );
  AND U36326 ( .A(a[36]), .B(b[39]), .Z(n31330) );
  XOR U36327 ( .A(n31336), .B(n31337), .Z(n30891) );
  ANDN U36328 ( .B(n31338), .A(n31339), .Z(n31336) );
  AND U36329 ( .A(a[37]), .B(b[38]), .Z(n31335) );
  XOR U36330 ( .A(n31341), .B(n31342), .Z(n30896) );
  ANDN U36331 ( .B(n31343), .A(n31344), .Z(n31341) );
  AND U36332 ( .A(a[38]), .B(b[37]), .Z(n31340) );
  XOR U36333 ( .A(n31346), .B(n31347), .Z(n30901) );
  ANDN U36334 ( .B(n31348), .A(n31349), .Z(n31346) );
  AND U36335 ( .A(a[39]), .B(b[36]), .Z(n31345) );
  XOR U36336 ( .A(n31351), .B(n31352), .Z(n30906) );
  ANDN U36337 ( .B(n31353), .A(n31354), .Z(n31351) );
  AND U36338 ( .A(a[40]), .B(b[35]), .Z(n31350) );
  XOR U36339 ( .A(n31356), .B(n31357), .Z(n30911) );
  ANDN U36340 ( .B(n31358), .A(n31359), .Z(n31356) );
  AND U36341 ( .A(a[41]), .B(b[34]), .Z(n31355) );
  XOR U36342 ( .A(n31361), .B(n31362), .Z(n30916) );
  ANDN U36343 ( .B(n31363), .A(n31364), .Z(n31361) );
  AND U36344 ( .A(a[42]), .B(b[33]), .Z(n31360) );
  XOR U36345 ( .A(n31366), .B(n31367), .Z(n30921) );
  ANDN U36346 ( .B(n31368), .A(n31369), .Z(n31366) );
  AND U36347 ( .A(a[43]), .B(b[32]), .Z(n31365) );
  XOR U36348 ( .A(n31371), .B(n31372), .Z(n30926) );
  ANDN U36349 ( .B(n31373), .A(n31374), .Z(n31371) );
  AND U36350 ( .A(a[44]), .B(b[31]), .Z(n31370) );
  XOR U36351 ( .A(n31376), .B(n31377), .Z(n30931) );
  ANDN U36352 ( .B(n31378), .A(n31379), .Z(n31376) );
  AND U36353 ( .A(a[45]), .B(b[30]), .Z(n31375) );
  XOR U36354 ( .A(n31381), .B(n31382), .Z(n30936) );
  ANDN U36355 ( .B(n31383), .A(n31384), .Z(n31381) );
  AND U36356 ( .A(a[46]), .B(b[29]), .Z(n31380) );
  XOR U36357 ( .A(n31386), .B(n31387), .Z(n30941) );
  ANDN U36358 ( .B(n31388), .A(n31389), .Z(n31386) );
  AND U36359 ( .A(a[47]), .B(b[28]), .Z(n31385) );
  XOR U36360 ( .A(n31391), .B(n31392), .Z(n30946) );
  ANDN U36361 ( .B(n31393), .A(n31394), .Z(n31391) );
  AND U36362 ( .A(a[48]), .B(b[27]), .Z(n31390) );
  XOR U36363 ( .A(n31396), .B(n31397), .Z(n30951) );
  ANDN U36364 ( .B(n31398), .A(n31399), .Z(n31396) );
  AND U36365 ( .A(a[49]), .B(b[26]), .Z(n31395) );
  XOR U36366 ( .A(n31401), .B(n31402), .Z(n30956) );
  ANDN U36367 ( .B(n31403), .A(n31404), .Z(n31401) );
  AND U36368 ( .A(a[50]), .B(b[25]), .Z(n31400) );
  XOR U36369 ( .A(n31406), .B(n31407), .Z(n30961) );
  ANDN U36370 ( .B(n31408), .A(n31409), .Z(n31406) );
  AND U36371 ( .A(a[51]), .B(b[24]), .Z(n31405) );
  XOR U36372 ( .A(n31411), .B(n31412), .Z(n30966) );
  ANDN U36373 ( .B(n31413), .A(n31414), .Z(n31411) );
  AND U36374 ( .A(a[52]), .B(b[23]), .Z(n31410) );
  XOR U36375 ( .A(n31416), .B(n31417), .Z(n30971) );
  ANDN U36376 ( .B(n31418), .A(n31419), .Z(n31416) );
  AND U36377 ( .A(a[53]), .B(b[22]), .Z(n31415) );
  XOR U36378 ( .A(n31421), .B(n31422), .Z(n30976) );
  ANDN U36379 ( .B(n31423), .A(n31424), .Z(n31421) );
  AND U36380 ( .A(a[54]), .B(b[21]), .Z(n31420) );
  XOR U36381 ( .A(n31426), .B(n31427), .Z(n30981) );
  ANDN U36382 ( .B(n31428), .A(n31429), .Z(n31426) );
  AND U36383 ( .A(a[55]), .B(b[20]), .Z(n31425) );
  XOR U36384 ( .A(n31431), .B(n31432), .Z(n30986) );
  ANDN U36385 ( .B(n31433), .A(n31434), .Z(n31431) );
  AND U36386 ( .A(a[56]), .B(b[19]), .Z(n31430) );
  XOR U36387 ( .A(n31436), .B(n31437), .Z(n30991) );
  ANDN U36388 ( .B(n31438), .A(n31439), .Z(n31436) );
  AND U36389 ( .A(a[57]), .B(b[18]), .Z(n31435) );
  XOR U36390 ( .A(n31441), .B(n31442), .Z(n30996) );
  ANDN U36391 ( .B(n31443), .A(n31444), .Z(n31441) );
  AND U36392 ( .A(a[58]), .B(b[17]), .Z(n31440) );
  XOR U36393 ( .A(n31446), .B(n31447), .Z(n31001) );
  ANDN U36394 ( .B(n31448), .A(n31449), .Z(n31446) );
  AND U36395 ( .A(a[59]), .B(b[16]), .Z(n31445) );
  XOR U36396 ( .A(n31451), .B(n31452), .Z(n31006) );
  ANDN U36397 ( .B(n31453), .A(n31454), .Z(n31451) );
  AND U36398 ( .A(a[60]), .B(b[15]), .Z(n31450) );
  XOR U36399 ( .A(n31456), .B(n31457), .Z(n31011) );
  ANDN U36400 ( .B(n31458), .A(n31459), .Z(n31456) );
  AND U36401 ( .A(a[61]), .B(b[14]), .Z(n31455) );
  XOR U36402 ( .A(n31461), .B(n31462), .Z(n31016) );
  ANDN U36403 ( .B(n31463), .A(n31464), .Z(n31461) );
  AND U36404 ( .A(a[62]), .B(b[13]), .Z(n31460) );
  XOR U36405 ( .A(n31466), .B(n31467), .Z(n31021) );
  ANDN U36406 ( .B(n31468), .A(n31469), .Z(n31466) );
  AND U36407 ( .A(a[63]), .B(b[12]), .Z(n31465) );
  XOR U36408 ( .A(n31471), .B(n31472), .Z(n31026) );
  ANDN U36409 ( .B(n31473), .A(n31474), .Z(n31471) );
  AND U36410 ( .A(a[64]), .B(b[11]), .Z(n31470) );
  XOR U36411 ( .A(n31476), .B(n31477), .Z(n31031) );
  ANDN U36412 ( .B(n31478), .A(n31479), .Z(n31476) );
  AND U36413 ( .A(a[65]), .B(b[10]), .Z(n31475) );
  XOR U36414 ( .A(n31481), .B(n31482), .Z(n31036) );
  ANDN U36415 ( .B(n31483), .A(n31484), .Z(n31481) );
  AND U36416 ( .A(b[9]), .B(a[66]), .Z(n31480) );
  XOR U36417 ( .A(n31486), .B(n31487), .Z(n31041) );
  ANDN U36418 ( .B(n31488), .A(n31489), .Z(n31486) );
  AND U36419 ( .A(b[8]), .B(a[67]), .Z(n31485) );
  XOR U36420 ( .A(n31491), .B(n31492), .Z(n31046) );
  ANDN U36421 ( .B(n31493), .A(n31494), .Z(n31491) );
  AND U36422 ( .A(b[7]), .B(a[68]), .Z(n31490) );
  XOR U36423 ( .A(n31496), .B(n31497), .Z(n31051) );
  ANDN U36424 ( .B(n31498), .A(n31499), .Z(n31496) );
  AND U36425 ( .A(b[6]), .B(a[69]), .Z(n31495) );
  XOR U36426 ( .A(n31501), .B(n31502), .Z(n31056) );
  ANDN U36427 ( .B(n31503), .A(n31504), .Z(n31501) );
  AND U36428 ( .A(b[5]), .B(a[70]), .Z(n31500) );
  XOR U36429 ( .A(n31506), .B(n31507), .Z(n31061) );
  ANDN U36430 ( .B(n31508), .A(n31509), .Z(n31506) );
  AND U36431 ( .A(b[4]), .B(a[71]), .Z(n31505) );
  XOR U36432 ( .A(n31511), .B(n31512), .Z(n31066) );
  ANDN U36433 ( .B(n31078), .A(n31079), .Z(n31511) );
  AND U36434 ( .A(b[2]), .B(a[72]), .Z(n31513) );
  XNOR U36435 ( .A(n31508), .B(n31512), .Z(n31514) );
  XOR U36436 ( .A(n31515), .B(n31516), .Z(n31512) );
  OR U36437 ( .A(n31081), .B(n31082), .Z(n31516) );
  XNOR U36438 ( .A(n31518), .B(n31519), .Z(n31517) );
  XOR U36439 ( .A(n31518), .B(n31521), .Z(n31081) );
  NAND U36440 ( .A(b[1]), .B(a[72]), .Z(n31521) );
  IV U36441 ( .A(n31515), .Z(n31518) );
  NANDN U36442 ( .A(n61), .B(n62), .Z(n31515) );
  XOR U36443 ( .A(n31522), .B(n31523), .Z(n62) );
  NAND U36444 ( .A(a[72]), .B(b[0]), .Z(n61) );
  XNOR U36445 ( .A(n31503), .B(n31507), .Z(n31524) );
  XNOR U36446 ( .A(n31498), .B(n31502), .Z(n31525) );
  XNOR U36447 ( .A(n31493), .B(n31497), .Z(n31526) );
  XNOR U36448 ( .A(n31488), .B(n31492), .Z(n31527) );
  XNOR U36449 ( .A(n31483), .B(n31487), .Z(n31528) );
  XNOR U36450 ( .A(n31478), .B(n31482), .Z(n31529) );
  XNOR U36451 ( .A(n31473), .B(n31477), .Z(n31530) );
  XNOR U36452 ( .A(n31468), .B(n31472), .Z(n31531) );
  XNOR U36453 ( .A(n31463), .B(n31467), .Z(n31532) );
  XNOR U36454 ( .A(n31458), .B(n31462), .Z(n31533) );
  XNOR U36455 ( .A(n31453), .B(n31457), .Z(n31534) );
  XNOR U36456 ( .A(n31448), .B(n31452), .Z(n31535) );
  XNOR U36457 ( .A(n31443), .B(n31447), .Z(n31536) );
  XNOR U36458 ( .A(n31438), .B(n31442), .Z(n31537) );
  XNOR U36459 ( .A(n31433), .B(n31437), .Z(n31538) );
  XNOR U36460 ( .A(n31428), .B(n31432), .Z(n31539) );
  XNOR U36461 ( .A(n31423), .B(n31427), .Z(n31540) );
  XNOR U36462 ( .A(n31418), .B(n31422), .Z(n31541) );
  XNOR U36463 ( .A(n31413), .B(n31417), .Z(n31542) );
  XNOR U36464 ( .A(n31408), .B(n31412), .Z(n31543) );
  XNOR U36465 ( .A(n31403), .B(n31407), .Z(n31544) );
  XNOR U36466 ( .A(n31398), .B(n31402), .Z(n31545) );
  XNOR U36467 ( .A(n31393), .B(n31397), .Z(n31546) );
  XNOR U36468 ( .A(n31388), .B(n31392), .Z(n31547) );
  XNOR U36469 ( .A(n31383), .B(n31387), .Z(n31548) );
  XNOR U36470 ( .A(n31378), .B(n31382), .Z(n31549) );
  XNOR U36471 ( .A(n31373), .B(n31377), .Z(n31550) );
  XNOR U36472 ( .A(n31368), .B(n31372), .Z(n31551) );
  XNOR U36473 ( .A(n31363), .B(n31367), .Z(n31552) );
  XNOR U36474 ( .A(n31358), .B(n31362), .Z(n31553) );
  XNOR U36475 ( .A(n31353), .B(n31357), .Z(n31554) );
  XNOR U36476 ( .A(n31348), .B(n31352), .Z(n31555) );
  XNOR U36477 ( .A(n31343), .B(n31347), .Z(n31556) );
  XNOR U36478 ( .A(n31338), .B(n31342), .Z(n31557) );
  XNOR U36479 ( .A(n31333), .B(n31337), .Z(n31558) );
  XNOR U36480 ( .A(n31328), .B(n31332), .Z(n31559) );
  XNOR U36481 ( .A(n31323), .B(n31327), .Z(n31560) );
  XNOR U36482 ( .A(n31318), .B(n31322), .Z(n31561) );
  XNOR U36483 ( .A(n31313), .B(n31317), .Z(n31562) );
  XNOR U36484 ( .A(n31308), .B(n31312), .Z(n31563) );
  XNOR U36485 ( .A(n31303), .B(n31307), .Z(n31564) );
  XNOR U36486 ( .A(n31298), .B(n31302), .Z(n31565) );
  XNOR U36487 ( .A(n31293), .B(n31297), .Z(n31566) );
  XNOR U36488 ( .A(n31288), .B(n31292), .Z(n31567) );
  XNOR U36489 ( .A(n31283), .B(n31287), .Z(n31568) );
  XNOR U36490 ( .A(n31278), .B(n31282), .Z(n31569) );
  XNOR U36491 ( .A(n31273), .B(n31277), .Z(n31570) );
  XNOR U36492 ( .A(n31268), .B(n31272), .Z(n31571) );
  XNOR U36493 ( .A(n31263), .B(n31267), .Z(n31572) );
  XNOR U36494 ( .A(n31258), .B(n31262), .Z(n31573) );
  XNOR U36495 ( .A(n31253), .B(n31257), .Z(n31574) );
  XNOR U36496 ( .A(n31248), .B(n31252), .Z(n31575) );
  XNOR U36497 ( .A(n31243), .B(n31247), .Z(n31576) );
  XNOR U36498 ( .A(n31238), .B(n31242), .Z(n31577) );
  XNOR U36499 ( .A(n31233), .B(n31237), .Z(n31578) );
  XNOR U36500 ( .A(n31228), .B(n31232), .Z(n31579) );
  XNOR U36501 ( .A(n31223), .B(n31227), .Z(n31580) );
  XNOR U36502 ( .A(n31218), .B(n31222), .Z(n31581) );
  XNOR U36503 ( .A(n31213), .B(n31217), .Z(n31582) );
  XNOR U36504 ( .A(n31208), .B(n31212), .Z(n31583) );
  XNOR U36505 ( .A(n31203), .B(n31207), .Z(n31584) );
  XNOR U36506 ( .A(n31198), .B(n31202), .Z(n31585) );
  XNOR U36507 ( .A(n31193), .B(n31197), .Z(n31586) );
  XNOR U36508 ( .A(n31188), .B(n31192), .Z(n31587) );
  XNOR U36509 ( .A(n31183), .B(n31187), .Z(n31588) );
  XNOR U36510 ( .A(n31178), .B(n31182), .Z(n31589) );
  XNOR U36511 ( .A(n31173), .B(n31177), .Z(n31590) );
  XNOR U36512 ( .A(n31168), .B(n31172), .Z(n31591) );
  XNOR U36513 ( .A(n31163), .B(n31167), .Z(n31592) );
  XNOR U36514 ( .A(n31158), .B(n31162), .Z(n31593) );
  XOR U36515 ( .A(n31594), .B(n31157), .Z(n31158) );
  AND U36516 ( .A(a[0]), .B(b[74]), .Z(n31594) );
  XNOR U36517 ( .A(n31595), .B(n31157), .Z(n31159) );
  XNOR U36518 ( .A(n31596), .B(n31597), .Z(n31157) );
  ANDN U36519 ( .B(n31598), .A(n31599), .Z(n31596) );
  AND U36520 ( .A(a[1]), .B(b[73]), .Z(n31595) );
  XOR U36521 ( .A(n31601), .B(n31602), .Z(n31162) );
  ANDN U36522 ( .B(n31603), .A(n31604), .Z(n31601) );
  AND U36523 ( .A(a[2]), .B(b[72]), .Z(n31600) );
  XOR U36524 ( .A(n31606), .B(n31607), .Z(n31167) );
  ANDN U36525 ( .B(n31608), .A(n31609), .Z(n31606) );
  AND U36526 ( .A(a[3]), .B(b[71]), .Z(n31605) );
  XOR U36527 ( .A(n31611), .B(n31612), .Z(n31172) );
  ANDN U36528 ( .B(n31613), .A(n31614), .Z(n31611) );
  AND U36529 ( .A(a[4]), .B(b[70]), .Z(n31610) );
  XOR U36530 ( .A(n31616), .B(n31617), .Z(n31177) );
  ANDN U36531 ( .B(n31618), .A(n31619), .Z(n31616) );
  AND U36532 ( .A(a[5]), .B(b[69]), .Z(n31615) );
  XOR U36533 ( .A(n31621), .B(n31622), .Z(n31182) );
  ANDN U36534 ( .B(n31623), .A(n31624), .Z(n31621) );
  AND U36535 ( .A(a[6]), .B(b[68]), .Z(n31620) );
  XOR U36536 ( .A(n31626), .B(n31627), .Z(n31187) );
  ANDN U36537 ( .B(n31628), .A(n31629), .Z(n31626) );
  AND U36538 ( .A(a[7]), .B(b[67]), .Z(n31625) );
  XOR U36539 ( .A(n31631), .B(n31632), .Z(n31192) );
  ANDN U36540 ( .B(n31633), .A(n31634), .Z(n31631) );
  AND U36541 ( .A(a[8]), .B(b[66]), .Z(n31630) );
  XOR U36542 ( .A(n31636), .B(n31637), .Z(n31197) );
  ANDN U36543 ( .B(n31638), .A(n31639), .Z(n31636) );
  AND U36544 ( .A(a[9]), .B(b[65]), .Z(n31635) );
  XOR U36545 ( .A(n31641), .B(n31642), .Z(n31202) );
  ANDN U36546 ( .B(n31643), .A(n31644), .Z(n31641) );
  AND U36547 ( .A(a[10]), .B(b[64]), .Z(n31640) );
  XOR U36548 ( .A(n31646), .B(n31647), .Z(n31207) );
  ANDN U36549 ( .B(n31648), .A(n31649), .Z(n31646) );
  AND U36550 ( .A(a[11]), .B(b[63]), .Z(n31645) );
  XOR U36551 ( .A(n31651), .B(n31652), .Z(n31212) );
  ANDN U36552 ( .B(n31653), .A(n31654), .Z(n31651) );
  AND U36553 ( .A(a[12]), .B(b[62]), .Z(n31650) );
  XOR U36554 ( .A(n31656), .B(n31657), .Z(n31217) );
  ANDN U36555 ( .B(n31658), .A(n31659), .Z(n31656) );
  AND U36556 ( .A(a[13]), .B(b[61]), .Z(n31655) );
  XOR U36557 ( .A(n31661), .B(n31662), .Z(n31222) );
  ANDN U36558 ( .B(n31663), .A(n31664), .Z(n31661) );
  AND U36559 ( .A(a[14]), .B(b[60]), .Z(n31660) );
  XOR U36560 ( .A(n31666), .B(n31667), .Z(n31227) );
  ANDN U36561 ( .B(n31668), .A(n31669), .Z(n31666) );
  AND U36562 ( .A(a[15]), .B(b[59]), .Z(n31665) );
  XOR U36563 ( .A(n31671), .B(n31672), .Z(n31232) );
  ANDN U36564 ( .B(n31673), .A(n31674), .Z(n31671) );
  AND U36565 ( .A(a[16]), .B(b[58]), .Z(n31670) );
  XOR U36566 ( .A(n31676), .B(n31677), .Z(n31237) );
  ANDN U36567 ( .B(n31678), .A(n31679), .Z(n31676) );
  AND U36568 ( .A(a[17]), .B(b[57]), .Z(n31675) );
  XOR U36569 ( .A(n31681), .B(n31682), .Z(n31242) );
  ANDN U36570 ( .B(n31683), .A(n31684), .Z(n31681) );
  AND U36571 ( .A(a[18]), .B(b[56]), .Z(n31680) );
  XOR U36572 ( .A(n31686), .B(n31687), .Z(n31247) );
  ANDN U36573 ( .B(n31688), .A(n31689), .Z(n31686) );
  AND U36574 ( .A(a[19]), .B(b[55]), .Z(n31685) );
  XOR U36575 ( .A(n31691), .B(n31692), .Z(n31252) );
  ANDN U36576 ( .B(n31693), .A(n31694), .Z(n31691) );
  AND U36577 ( .A(a[20]), .B(b[54]), .Z(n31690) );
  XOR U36578 ( .A(n31696), .B(n31697), .Z(n31257) );
  ANDN U36579 ( .B(n31698), .A(n31699), .Z(n31696) );
  AND U36580 ( .A(a[21]), .B(b[53]), .Z(n31695) );
  XOR U36581 ( .A(n31701), .B(n31702), .Z(n31262) );
  ANDN U36582 ( .B(n31703), .A(n31704), .Z(n31701) );
  AND U36583 ( .A(a[22]), .B(b[52]), .Z(n31700) );
  XOR U36584 ( .A(n31706), .B(n31707), .Z(n31267) );
  ANDN U36585 ( .B(n31708), .A(n31709), .Z(n31706) );
  AND U36586 ( .A(a[23]), .B(b[51]), .Z(n31705) );
  XOR U36587 ( .A(n31711), .B(n31712), .Z(n31272) );
  ANDN U36588 ( .B(n31713), .A(n31714), .Z(n31711) );
  AND U36589 ( .A(a[24]), .B(b[50]), .Z(n31710) );
  XOR U36590 ( .A(n31716), .B(n31717), .Z(n31277) );
  ANDN U36591 ( .B(n31718), .A(n31719), .Z(n31716) );
  AND U36592 ( .A(a[25]), .B(b[49]), .Z(n31715) );
  XOR U36593 ( .A(n31721), .B(n31722), .Z(n31282) );
  ANDN U36594 ( .B(n31723), .A(n31724), .Z(n31721) );
  AND U36595 ( .A(a[26]), .B(b[48]), .Z(n31720) );
  XOR U36596 ( .A(n31726), .B(n31727), .Z(n31287) );
  ANDN U36597 ( .B(n31728), .A(n31729), .Z(n31726) );
  AND U36598 ( .A(a[27]), .B(b[47]), .Z(n31725) );
  XOR U36599 ( .A(n31731), .B(n31732), .Z(n31292) );
  ANDN U36600 ( .B(n31733), .A(n31734), .Z(n31731) );
  AND U36601 ( .A(a[28]), .B(b[46]), .Z(n31730) );
  XOR U36602 ( .A(n31736), .B(n31737), .Z(n31297) );
  ANDN U36603 ( .B(n31738), .A(n31739), .Z(n31736) );
  AND U36604 ( .A(a[29]), .B(b[45]), .Z(n31735) );
  XOR U36605 ( .A(n31741), .B(n31742), .Z(n31302) );
  ANDN U36606 ( .B(n31743), .A(n31744), .Z(n31741) );
  AND U36607 ( .A(a[30]), .B(b[44]), .Z(n31740) );
  XOR U36608 ( .A(n31746), .B(n31747), .Z(n31307) );
  ANDN U36609 ( .B(n31748), .A(n31749), .Z(n31746) );
  AND U36610 ( .A(a[31]), .B(b[43]), .Z(n31745) );
  XOR U36611 ( .A(n31751), .B(n31752), .Z(n31312) );
  ANDN U36612 ( .B(n31753), .A(n31754), .Z(n31751) );
  AND U36613 ( .A(a[32]), .B(b[42]), .Z(n31750) );
  XOR U36614 ( .A(n31756), .B(n31757), .Z(n31317) );
  ANDN U36615 ( .B(n31758), .A(n31759), .Z(n31756) );
  AND U36616 ( .A(a[33]), .B(b[41]), .Z(n31755) );
  XOR U36617 ( .A(n31761), .B(n31762), .Z(n31322) );
  ANDN U36618 ( .B(n31763), .A(n31764), .Z(n31761) );
  AND U36619 ( .A(a[34]), .B(b[40]), .Z(n31760) );
  XOR U36620 ( .A(n31766), .B(n31767), .Z(n31327) );
  ANDN U36621 ( .B(n31768), .A(n31769), .Z(n31766) );
  AND U36622 ( .A(a[35]), .B(b[39]), .Z(n31765) );
  XOR U36623 ( .A(n31771), .B(n31772), .Z(n31332) );
  ANDN U36624 ( .B(n31773), .A(n31774), .Z(n31771) );
  AND U36625 ( .A(a[36]), .B(b[38]), .Z(n31770) );
  XOR U36626 ( .A(n31776), .B(n31777), .Z(n31337) );
  ANDN U36627 ( .B(n31778), .A(n31779), .Z(n31776) );
  AND U36628 ( .A(a[37]), .B(b[37]), .Z(n31775) );
  XOR U36629 ( .A(n31781), .B(n31782), .Z(n31342) );
  ANDN U36630 ( .B(n31783), .A(n31784), .Z(n31781) );
  AND U36631 ( .A(a[38]), .B(b[36]), .Z(n31780) );
  XOR U36632 ( .A(n31786), .B(n31787), .Z(n31347) );
  ANDN U36633 ( .B(n31788), .A(n31789), .Z(n31786) );
  AND U36634 ( .A(a[39]), .B(b[35]), .Z(n31785) );
  XOR U36635 ( .A(n31791), .B(n31792), .Z(n31352) );
  ANDN U36636 ( .B(n31793), .A(n31794), .Z(n31791) );
  AND U36637 ( .A(a[40]), .B(b[34]), .Z(n31790) );
  XOR U36638 ( .A(n31796), .B(n31797), .Z(n31357) );
  ANDN U36639 ( .B(n31798), .A(n31799), .Z(n31796) );
  AND U36640 ( .A(a[41]), .B(b[33]), .Z(n31795) );
  XOR U36641 ( .A(n31801), .B(n31802), .Z(n31362) );
  ANDN U36642 ( .B(n31803), .A(n31804), .Z(n31801) );
  AND U36643 ( .A(a[42]), .B(b[32]), .Z(n31800) );
  XOR U36644 ( .A(n31806), .B(n31807), .Z(n31367) );
  ANDN U36645 ( .B(n31808), .A(n31809), .Z(n31806) );
  AND U36646 ( .A(a[43]), .B(b[31]), .Z(n31805) );
  XOR U36647 ( .A(n31811), .B(n31812), .Z(n31372) );
  ANDN U36648 ( .B(n31813), .A(n31814), .Z(n31811) );
  AND U36649 ( .A(a[44]), .B(b[30]), .Z(n31810) );
  XOR U36650 ( .A(n31816), .B(n31817), .Z(n31377) );
  ANDN U36651 ( .B(n31818), .A(n31819), .Z(n31816) );
  AND U36652 ( .A(a[45]), .B(b[29]), .Z(n31815) );
  XOR U36653 ( .A(n31821), .B(n31822), .Z(n31382) );
  ANDN U36654 ( .B(n31823), .A(n31824), .Z(n31821) );
  AND U36655 ( .A(a[46]), .B(b[28]), .Z(n31820) );
  XOR U36656 ( .A(n31826), .B(n31827), .Z(n31387) );
  ANDN U36657 ( .B(n31828), .A(n31829), .Z(n31826) );
  AND U36658 ( .A(a[47]), .B(b[27]), .Z(n31825) );
  XOR U36659 ( .A(n31831), .B(n31832), .Z(n31392) );
  ANDN U36660 ( .B(n31833), .A(n31834), .Z(n31831) );
  AND U36661 ( .A(a[48]), .B(b[26]), .Z(n31830) );
  XOR U36662 ( .A(n31836), .B(n31837), .Z(n31397) );
  ANDN U36663 ( .B(n31838), .A(n31839), .Z(n31836) );
  AND U36664 ( .A(a[49]), .B(b[25]), .Z(n31835) );
  XOR U36665 ( .A(n31841), .B(n31842), .Z(n31402) );
  ANDN U36666 ( .B(n31843), .A(n31844), .Z(n31841) );
  AND U36667 ( .A(a[50]), .B(b[24]), .Z(n31840) );
  XOR U36668 ( .A(n31846), .B(n31847), .Z(n31407) );
  ANDN U36669 ( .B(n31848), .A(n31849), .Z(n31846) );
  AND U36670 ( .A(a[51]), .B(b[23]), .Z(n31845) );
  XOR U36671 ( .A(n31851), .B(n31852), .Z(n31412) );
  ANDN U36672 ( .B(n31853), .A(n31854), .Z(n31851) );
  AND U36673 ( .A(a[52]), .B(b[22]), .Z(n31850) );
  XOR U36674 ( .A(n31856), .B(n31857), .Z(n31417) );
  ANDN U36675 ( .B(n31858), .A(n31859), .Z(n31856) );
  AND U36676 ( .A(a[53]), .B(b[21]), .Z(n31855) );
  XOR U36677 ( .A(n31861), .B(n31862), .Z(n31422) );
  ANDN U36678 ( .B(n31863), .A(n31864), .Z(n31861) );
  AND U36679 ( .A(a[54]), .B(b[20]), .Z(n31860) );
  XOR U36680 ( .A(n31866), .B(n31867), .Z(n31427) );
  ANDN U36681 ( .B(n31868), .A(n31869), .Z(n31866) );
  AND U36682 ( .A(a[55]), .B(b[19]), .Z(n31865) );
  XOR U36683 ( .A(n31871), .B(n31872), .Z(n31432) );
  ANDN U36684 ( .B(n31873), .A(n31874), .Z(n31871) );
  AND U36685 ( .A(a[56]), .B(b[18]), .Z(n31870) );
  XOR U36686 ( .A(n31876), .B(n31877), .Z(n31437) );
  ANDN U36687 ( .B(n31878), .A(n31879), .Z(n31876) );
  AND U36688 ( .A(a[57]), .B(b[17]), .Z(n31875) );
  XOR U36689 ( .A(n31881), .B(n31882), .Z(n31442) );
  ANDN U36690 ( .B(n31883), .A(n31884), .Z(n31881) );
  AND U36691 ( .A(a[58]), .B(b[16]), .Z(n31880) );
  XOR U36692 ( .A(n31886), .B(n31887), .Z(n31447) );
  ANDN U36693 ( .B(n31888), .A(n31889), .Z(n31886) );
  AND U36694 ( .A(a[59]), .B(b[15]), .Z(n31885) );
  XOR U36695 ( .A(n31891), .B(n31892), .Z(n31452) );
  ANDN U36696 ( .B(n31893), .A(n31894), .Z(n31891) );
  AND U36697 ( .A(a[60]), .B(b[14]), .Z(n31890) );
  XOR U36698 ( .A(n31896), .B(n31897), .Z(n31457) );
  ANDN U36699 ( .B(n31898), .A(n31899), .Z(n31896) );
  AND U36700 ( .A(a[61]), .B(b[13]), .Z(n31895) );
  XOR U36701 ( .A(n31901), .B(n31902), .Z(n31462) );
  ANDN U36702 ( .B(n31903), .A(n31904), .Z(n31901) );
  AND U36703 ( .A(a[62]), .B(b[12]), .Z(n31900) );
  XOR U36704 ( .A(n31906), .B(n31907), .Z(n31467) );
  ANDN U36705 ( .B(n31908), .A(n31909), .Z(n31906) );
  AND U36706 ( .A(a[63]), .B(b[11]), .Z(n31905) );
  XOR U36707 ( .A(n31911), .B(n31912), .Z(n31472) );
  ANDN U36708 ( .B(n31913), .A(n31914), .Z(n31911) );
  AND U36709 ( .A(a[64]), .B(b[10]), .Z(n31910) );
  XOR U36710 ( .A(n31916), .B(n31917), .Z(n31477) );
  ANDN U36711 ( .B(n31918), .A(n31919), .Z(n31916) );
  AND U36712 ( .A(b[9]), .B(a[65]), .Z(n31915) );
  XOR U36713 ( .A(n31921), .B(n31922), .Z(n31482) );
  ANDN U36714 ( .B(n31923), .A(n31924), .Z(n31921) );
  AND U36715 ( .A(b[8]), .B(a[66]), .Z(n31920) );
  XOR U36716 ( .A(n31926), .B(n31927), .Z(n31487) );
  ANDN U36717 ( .B(n31928), .A(n31929), .Z(n31926) );
  AND U36718 ( .A(b[7]), .B(a[67]), .Z(n31925) );
  XOR U36719 ( .A(n31931), .B(n31932), .Z(n31492) );
  ANDN U36720 ( .B(n31933), .A(n31934), .Z(n31931) );
  AND U36721 ( .A(b[6]), .B(a[68]), .Z(n31930) );
  XOR U36722 ( .A(n31936), .B(n31937), .Z(n31497) );
  ANDN U36723 ( .B(n31938), .A(n31939), .Z(n31936) );
  AND U36724 ( .A(b[5]), .B(a[69]), .Z(n31935) );
  XOR U36725 ( .A(n31941), .B(n31942), .Z(n31502) );
  ANDN U36726 ( .B(n31943), .A(n31944), .Z(n31941) );
  AND U36727 ( .A(b[4]), .B(a[70]), .Z(n31940) );
  XOR U36728 ( .A(n31946), .B(n31947), .Z(n31507) );
  ANDN U36729 ( .B(n31519), .A(n31520), .Z(n31946) );
  AND U36730 ( .A(b[2]), .B(a[71]), .Z(n31948) );
  XNOR U36731 ( .A(n31943), .B(n31947), .Z(n31949) );
  XOR U36732 ( .A(n31950), .B(n31951), .Z(n31947) );
  OR U36733 ( .A(n31522), .B(n31523), .Z(n31951) );
  XNOR U36734 ( .A(n31953), .B(n31954), .Z(n31952) );
  XOR U36735 ( .A(n31953), .B(n31956), .Z(n31522) );
  NAND U36736 ( .A(b[1]), .B(a[71]), .Z(n31956) );
  IV U36737 ( .A(n31950), .Z(n31953) );
  NANDN U36738 ( .A(n63), .B(n64), .Z(n31950) );
  XOR U36739 ( .A(n31957), .B(n31958), .Z(n64) );
  NAND U36740 ( .A(a[71]), .B(b[0]), .Z(n63) );
  XNOR U36741 ( .A(n31938), .B(n31942), .Z(n31959) );
  XNOR U36742 ( .A(n31933), .B(n31937), .Z(n31960) );
  XNOR U36743 ( .A(n31928), .B(n31932), .Z(n31961) );
  XNOR U36744 ( .A(n31923), .B(n31927), .Z(n31962) );
  XNOR U36745 ( .A(n31918), .B(n31922), .Z(n31963) );
  XNOR U36746 ( .A(n31913), .B(n31917), .Z(n31964) );
  XNOR U36747 ( .A(n31908), .B(n31912), .Z(n31965) );
  XNOR U36748 ( .A(n31903), .B(n31907), .Z(n31966) );
  XNOR U36749 ( .A(n31898), .B(n31902), .Z(n31967) );
  XNOR U36750 ( .A(n31893), .B(n31897), .Z(n31968) );
  XNOR U36751 ( .A(n31888), .B(n31892), .Z(n31969) );
  XNOR U36752 ( .A(n31883), .B(n31887), .Z(n31970) );
  XNOR U36753 ( .A(n31878), .B(n31882), .Z(n31971) );
  XNOR U36754 ( .A(n31873), .B(n31877), .Z(n31972) );
  XNOR U36755 ( .A(n31868), .B(n31872), .Z(n31973) );
  XNOR U36756 ( .A(n31863), .B(n31867), .Z(n31974) );
  XNOR U36757 ( .A(n31858), .B(n31862), .Z(n31975) );
  XNOR U36758 ( .A(n31853), .B(n31857), .Z(n31976) );
  XNOR U36759 ( .A(n31848), .B(n31852), .Z(n31977) );
  XNOR U36760 ( .A(n31843), .B(n31847), .Z(n31978) );
  XNOR U36761 ( .A(n31838), .B(n31842), .Z(n31979) );
  XNOR U36762 ( .A(n31833), .B(n31837), .Z(n31980) );
  XNOR U36763 ( .A(n31828), .B(n31832), .Z(n31981) );
  XNOR U36764 ( .A(n31823), .B(n31827), .Z(n31982) );
  XNOR U36765 ( .A(n31818), .B(n31822), .Z(n31983) );
  XNOR U36766 ( .A(n31813), .B(n31817), .Z(n31984) );
  XNOR U36767 ( .A(n31808), .B(n31812), .Z(n31985) );
  XNOR U36768 ( .A(n31803), .B(n31807), .Z(n31986) );
  XNOR U36769 ( .A(n31798), .B(n31802), .Z(n31987) );
  XNOR U36770 ( .A(n31793), .B(n31797), .Z(n31988) );
  XNOR U36771 ( .A(n31788), .B(n31792), .Z(n31989) );
  XNOR U36772 ( .A(n31783), .B(n31787), .Z(n31990) );
  XNOR U36773 ( .A(n31778), .B(n31782), .Z(n31991) );
  XNOR U36774 ( .A(n31773), .B(n31777), .Z(n31992) );
  XNOR U36775 ( .A(n31768), .B(n31772), .Z(n31993) );
  XNOR U36776 ( .A(n31763), .B(n31767), .Z(n31994) );
  XNOR U36777 ( .A(n31758), .B(n31762), .Z(n31995) );
  XNOR U36778 ( .A(n31753), .B(n31757), .Z(n31996) );
  XNOR U36779 ( .A(n31748), .B(n31752), .Z(n31997) );
  XNOR U36780 ( .A(n31743), .B(n31747), .Z(n31998) );
  XNOR U36781 ( .A(n31738), .B(n31742), .Z(n31999) );
  XNOR U36782 ( .A(n31733), .B(n31737), .Z(n32000) );
  XNOR U36783 ( .A(n31728), .B(n31732), .Z(n32001) );
  XNOR U36784 ( .A(n31723), .B(n31727), .Z(n32002) );
  XNOR U36785 ( .A(n31718), .B(n31722), .Z(n32003) );
  XNOR U36786 ( .A(n31713), .B(n31717), .Z(n32004) );
  XNOR U36787 ( .A(n31708), .B(n31712), .Z(n32005) );
  XNOR U36788 ( .A(n31703), .B(n31707), .Z(n32006) );
  XNOR U36789 ( .A(n31698), .B(n31702), .Z(n32007) );
  XNOR U36790 ( .A(n31693), .B(n31697), .Z(n32008) );
  XNOR U36791 ( .A(n31688), .B(n31692), .Z(n32009) );
  XNOR U36792 ( .A(n31683), .B(n31687), .Z(n32010) );
  XNOR U36793 ( .A(n31678), .B(n31682), .Z(n32011) );
  XNOR U36794 ( .A(n31673), .B(n31677), .Z(n32012) );
  XNOR U36795 ( .A(n31668), .B(n31672), .Z(n32013) );
  XNOR U36796 ( .A(n31663), .B(n31667), .Z(n32014) );
  XNOR U36797 ( .A(n31658), .B(n31662), .Z(n32015) );
  XNOR U36798 ( .A(n31653), .B(n31657), .Z(n32016) );
  XNOR U36799 ( .A(n31648), .B(n31652), .Z(n32017) );
  XNOR U36800 ( .A(n31643), .B(n31647), .Z(n32018) );
  XNOR U36801 ( .A(n31638), .B(n31642), .Z(n32019) );
  XNOR U36802 ( .A(n31633), .B(n31637), .Z(n32020) );
  XNOR U36803 ( .A(n31628), .B(n31632), .Z(n32021) );
  XNOR U36804 ( .A(n31623), .B(n31627), .Z(n32022) );
  XNOR U36805 ( .A(n31618), .B(n31622), .Z(n32023) );
  XNOR U36806 ( .A(n31613), .B(n31617), .Z(n32024) );
  XNOR U36807 ( .A(n31608), .B(n31612), .Z(n32025) );
  XNOR U36808 ( .A(n31603), .B(n31607), .Z(n32026) );
  XNOR U36809 ( .A(n31598), .B(n31602), .Z(n32027) );
  XNOR U36810 ( .A(n32028), .B(n31597), .Z(n31598) );
  AND U36811 ( .A(a[0]), .B(b[73]), .Z(n32028) );
  XOR U36812 ( .A(n32029), .B(n31597), .Z(n31599) );
  XNOR U36813 ( .A(n32030), .B(n32031), .Z(n31597) );
  ANDN U36814 ( .B(n32032), .A(n32033), .Z(n32030) );
  AND U36815 ( .A(a[1]), .B(b[72]), .Z(n32029) );
  XOR U36816 ( .A(n32035), .B(n32036), .Z(n31602) );
  ANDN U36817 ( .B(n32037), .A(n32038), .Z(n32035) );
  AND U36818 ( .A(a[2]), .B(b[71]), .Z(n32034) );
  XOR U36819 ( .A(n32040), .B(n32041), .Z(n31607) );
  ANDN U36820 ( .B(n32042), .A(n32043), .Z(n32040) );
  AND U36821 ( .A(a[3]), .B(b[70]), .Z(n32039) );
  XOR U36822 ( .A(n32045), .B(n32046), .Z(n31612) );
  ANDN U36823 ( .B(n32047), .A(n32048), .Z(n32045) );
  AND U36824 ( .A(a[4]), .B(b[69]), .Z(n32044) );
  XOR U36825 ( .A(n32050), .B(n32051), .Z(n31617) );
  ANDN U36826 ( .B(n32052), .A(n32053), .Z(n32050) );
  AND U36827 ( .A(a[5]), .B(b[68]), .Z(n32049) );
  XOR U36828 ( .A(n32055), .B(n32056), .Z(n31622) );
  ANDN U36829 ( .B(n32057), .A(n32058), .Z(n32055) );
  AND U36830 ( .A(a[6]), .B(b[67]), .Z(n32054) );
  XOR U36831 ( .A(n32060), .B(n32061), .Z(n31627) );
  ANDN U36832 ( .B(n32062), .A(n32063), .Z(n32060) );
  AND U36833 ( .A(a[7]), .B(b[66]), .Z(n32059) );
  XOR U36834 ( .A(n32065), .B(n32066), .Z(n31632) );
  ANDN U36835 ( .B(n32067), .A(n32068), .Z(n32065) );
  AND U36836 ( .A(a[8]), .B(b[65]), .Z(n32064) );
  XOR U36837 ( .A(n32070), .B(n32071), .Z(n31637) );
  ANDN U36838 ( .B(n32072), .A(n32073), .Z(n32070) );
  AND U36839 ( .A(a[9]), .B(b[64]), .Z(n32069) );
  XOR U36840 ( .A(n32075), .B(n32076), .Z(n31642) );
  ANDN U36841 ( .B(n32077), .A(n32078), .Z(n32075) );
  AND U36842 ( .A(a[10]), .B(b[63]), .Z(n32074) );
  XOR U36843 ( .A(n32080), .B(n32081), .Z(n31647) );
  ANDN U36844 ( .B(n32082), .A(n32083), .Z(n32080) );
  AND U36845 ( .A(a[11]), .B(b[62]), .Z(n32079) );
  XOR U36846 ( .A(n32085), .B(n32086), .Z(n31652) );
  ANDN U36847 ( .B(n32087), .A(n32088), .Z(n32085) );
  AND U36848 ( .A(a[12]), .B(b[61]), .Z(n32084) );
  XOR U36849 ( .A(n32090), .B(n32091), .Z(n31657) );
  ANDN U36850 ( .B(n32092), .A(n32093), .Z(n32090) );
  AND U36851 ( .A(a[13]), .B(b[60]), .Z(n32089) );
  XOR U36852 ( .A(n32095), .B(n32096), .Z(n31662) );
  ANDN U36853 ( .B(n32097), .A(n32098), .Z(n32095) );
  AND U36854 ( .A(a[14]), .B(b[59]), .Z(n32094) );
  XOR U36855 ( .A(n32100), .B(n32101), .Z(n31667) );
  ANDN U36856 ( .B(n32102), .A(n32103), .Z(n32100) );
  AND U36857 ( .A(a[15]), .B(b[58]), .Z(n32099) );
  XOR U36858 ( .A(n32105), .B(n32106), .Z(n31672) );
  ANDN U36859 ( .B(n32107), .A(n32108), .Z(n32105) );
  AND U36860 ( .A(a[16]), .B(b[57]), .Z(n32104) );
  XOR U36861 ( .A(n32110), .B(n32111), .Z(n31677) );
  ANDN U36862 ( .B(n32112), .A(n32113), .Z(n32110) );
  AND U36863 ( .A(a[17]), .B(b[56]), .Z(n32109) );
  XOR U36864 ( .A(n32115), .B(n32116), .Z(n31682) );
  ANDN U36865 ( .B(n32117), .A(n32118), .Z(n32115) );
  AND U36866 ( .A(a[18]), .B(b[55]), .Z(n32114) );
  XOR U36867 ( .A(n32120), .B(n32121), .Z(n31687) );
  ANDN U36868 ( .B(n32122), .A(n32123), .Z(n32120) );
  AND U36869 ( .A(a[19]), .B(b[54]), .Z(n32119) );
  XOR U36870 ( .A(n32125), .B(n32126), .Z(n31692) );
  ANDN U36871 ( .B(n32127), .A(n32128), .Z(n32125) );
  AND U36872 ( .A(a[20]), .B(b[53]), .Z(n32124) );
  XOR U36873 ( .A(n32130), .B(n32131), .Z(n31697) );
  ANDN U36874 ( .B(n32132), .A(n32133), .Z(n32130) );
  AND U36875 ( .A(a[21]), .B(b[52]), .Z(n32129) );
  XOR U36876 ( .A(n32135), .B(n32136), .Z(n31702) );
  ANDN U36877 ( .B(n32137), .A(n32138), .Z(n32135) );
  AND U36878 ( .A(a[22]), .B(b[51]), .Z(n32134) );
  XOR U36879 ( .A(n32140), .B(n32141), .Z(n31707) );
  ANDN U36880 ( .B(n32142), .A(n32143), .Z(n32140) );
  AND U36881 ( .A(a[23]), .B(b[50]), .Z(n32139) );
  XOR U36882 ( .A(n32145), .B(n32146), .Z(n31712) );
  ANDN U36883 ( .B(n32147), .A(n32148), .Z(n32145) );
  AND U36884 ( .A(a[24]), .B(b[49]), .Z(n32144) );
  XOR U36885 ( .A(n32150), .B(n32151), .Z(n31717) );
  ANDN U36886 ( .B(n32152), .A(n32153), .Z(n32150) );
  AND U36887 ( .A(a[25]), .B(b[48]), .Z(n32149) );
  XOR U36888 ( .A(n32155), .B(n32156), .Z(n31722) );
  ANDN U36889 ( .B(n32157), .A(n32158), .Z(n32155) );
  AND U36890 ( .A(a[26]), .B(b[47]), .Z(n32154) );
  XOR U36891 ( .A(n32160), .B(n32161), .Z(n31727) );
  ANDN U36892 ( .B(n32162), .A(n32163), .Z(n32160) );
  AND U36893 ( .A(a[27]), .B(b[46]), .Z(n32159) );
  XOR U36894 ( .A(n32165), .B(n32166), .Z(n31732) );
  ANDN U36895 ( .B(n32167), .A(n32168), .Z(n32165) );
  AND U36896 ( .A(a[28]), .B(b[45]), .Z(n32164) );
  XOR U36897 ( .A(n32170), .B(n32171), .Z(n31737) );
  ANDN U36898 ( .B(n32172), .A(n32173), .Z(n32170) );
  AND U36899 ( .A(a[29]), .B(b[44]), .Z(n32169) );
  XOR U36900 ( .A(n32175), .B(n32176), .Z(n31742) );
  ANDN U36901 ( .B(n32177), .A(n32178), .Z(n32175) );
  AND U36902 ( .A(a[30]), .B(b[43]), .Z(n32174) );
  XOR U36903 ( .A(n32180), .B(n32181), .Z(n31747) );
  ANDN U36904 ( .B(n32182), .A(n32183), .Z(n32180) );
  AND U36905 ( .A(a[31]), .B(b[42]), .Z(n32179) );
  XOR U36906 ( .A(n32185), .B(n32186), .Z(n31752) );
  ANDN U36907 ( .B(n32187), .A(n32188), .Z(n32185) );
  AND U36908 ( .A(a[32]), .B(b[41]), .Z(n32184) );
  XOR U36909 ( .A(n32190), .B(n32191), .Z(n31757) );
  ANDN U36910 ( .B(n32192), .A(n32193), .Z(n32190) );
  AND U36911 ( .A(a[33]), .B(b[40]), .Z(n32189) );
  XOR U36912 ( .A(n32195), .B(n32196), .Z(n31762) );
  ANDN U36913 ( .B(n32197), .A(n32198), .Z(n32195) );
  AND U36914 ( .A(a[34]), .B(b[39]), .Z(n32194) );
  XOR U36915 ( .A(n32200), .B(n32201), .Z(n31767) );
  ANDN U36916 ( .B(n32202), .A(n32203), .Z(n32200) );
  AND U36917 ( .A(a[35]), .B(b[38]), .Z(n32199) );
  XOR U36918 ( .A(n32205), .B(n32206), .Z(n31772) );
  ANDN U36919 ( .B(n32207), .A(n32208), .Z(n32205) );
  AND U36920 ( .A(a[36]), .B(b[37]), .Z(n32204) );
  XOR U36921 ( .A(n32210), .B(n32211), .Z(n31777) );
  ANDN U36922 ( .B(n32212), .A(n32213), .Z(n32210) );
  AND U36923 ( .A(a[37]), .B(b[36]), .Z(n32209) );
  XOR U36924 ( .A(n32215), .B(n32216), .Z(n31782) );
  ANDN U36925 ( .B(n32217), .A(n32218), .Z(n32215) );
  AND U36926 ( .A(a[38]), .B(b[35]), .Z(n32214) );
  XOR U36927 ( .A(n32220), .B(n32221), .Z(n31787) );
  ANDN U36928 ( .B(n32222), .A(n32223), .Z(n32220) );
  AND U36929 ( .A(a[39]), .B(b[34]), .Z(n32219) );
  XOR U36930 ( .A(n32225), .B(n32226), .Z(n31792) );
  ANDN U36931 ( .B(n32227), .A(n32228), .Z(n32225) );
  AND U36932 ( .A(a[40]), .B(b[33]), .Z(n32224) );
  XOR U36933 ( .A(n32230), .B(n32231), .Z(n31797) );
  ANDN U36934 ( .B(n32232), .A(n32233), .Z(n32230) );
  AND U36935 ( .A(a[41]), .B(b[32]), .Z(n32229) );
  XOR U36936 ( .A(n32235), .B(n32236), .Z(n31802) );
  ANDN U36937 ( .B(n32237), .A(n32238), .Z(n32235) );
  AND U36938 ( .A(a[42]), .B(b[31]), .Z(n32234) );
  XOR U36939 ( .A(n32240), .B(n32241), .Z(n31807) );
  ANDN U36940 ( .B(n32242), .A(n32243), .Z(n32240) );
  AND U36941 ( .A(a[43]), .B(b[30]), .Z(n32239) );
  XOR U36942 ( .A(n32245), .B(n32246), .Z(n31812) );
  ANDN U36943 ( .B(n32247), .A(n32248), .Z(n32245) );
  AND U36944 ( .A(a[44]), .B(b[29]), .Z(n32244) );
  XOR U36945 ( .A(n32250), .B(n32251), .Z(n31817) );
  ANDN U36946 ( .B(n32252), .A(n32253), .Z(n32250) );
  AND U36947 ( .A(a[45]), .B(b[28]), .Z(n32249) );
  XOR U36948 ( .A(n32255), .B(n32256), .Z(n31822) );
  ANDN U36949 ( .B(n32257), .A(n32258), .Z(n32255) );
  AND U36950 ( .A(a[46]), .B(b[27]), .Z(n32254) );
  XOR U36951 ( .A(n32260), .B(n32261), .Z(n31827) );
  ANDN U36952 ( .B(n32262), .A(n32263), .Z(n32260) );
  AND U36953 ( .A(a[47]), .B(b[26]), .Z(n32259) );
  XOR U36954 ( .A(n32265), .B(n32266), .Z(n31832) );
  ANDN U36955 ( .B(n32267), .A(n32268), .Z(n32265) );
  AND U36956 ( .A(a[48]), .B(b[25]), .Z(n32264) );
  XOR U36957 ( .A(n32270), .B(n32271), .Z(n31837) );
  ANDN U36958 ( .B(n32272), .A(n32273), .Z(n32270) );
  AND U36959 ( .A(a[49]), .B(b[24]), .Z(n32269) );
  XOR U36960 ( .A(n32275), .B(n32276), .Z(n31842) );
  ANDN U36961 ( .B(n32277), .A(n32278), .Z(n32275) );
  AND U36962 ( .A(a[50]), .B(b[23]), .Z(n32274) );
  XOR U36963 ( .A(n32280), .B(n32281), .Z(n31847) );
  ANDN U36964 ( .B(n32282), .A(n32283), .Z(n32280) );
  AND U36965 ( .A(a[51]), .B(b[22]), .Z(n32279) );
  XOR U36966 ( .A(n32285), .B(n32286), .Z(n31852) );
  ANDN U36967 ( .B(n32287), .A(n32288), .Z(n32285) );
  AND U36968 ( .A(a[52]), .B(b[21]), .Z(n32284) );
  XOR U36969 ( .A(n32290), .B(n32291), .Z(n31857) );
  ANDN U36970 ( .B(n32292), .A(n32293), .Z(n32290) );
  AND U36971 ( .A(a[53]), .B(b[20]), .Z(n32289) );
  XOR U36972 ( .A(n32295), .B(n32296), .Z(n31862) );
  ANDN U36973 ( .B(n32297), .A(n32298), .Z(n32295) );
  AND U36974 ( .A(a[54]), .B(b[19]), .Z(n32294) );
  XOR U36975 ( .A(n32300), .B(n32301), .Z(n31867) );
  ANDN U36976 ( .B(n32302), .A(n32303), .Z(n32300) );
  AND U36977 ( .A(a[55]), .B(b[18]), .Z(n32299) );
  XOR U36978 ( .A(n32305), .B(n32306), .Z(n31872) );
  ANDN U36979 ( .B(n32307), .A(n32308), .Z(n32305) );
  AND U36980 ( .A(a[56]), .B(b[17]), .Z(n32304) );
  XOR U36981 ( .A(n32310), .B(n32311), .Z(n31877) );
  ANDN U36982 ( .B(n32312), .A(n32313), .Z(n32310) );
  AND U36983 ( .A(a[57]), .B(b[16]), .Z(n32309) );
  XOR U36984 ( .A(n32315), .B(n32316), .Z(n31882) );
  ANDN U36985 ( .B(n32317), .A(n32318), .Z(n32315) );
  AND U36986 ( .A(a[58]), .B(b[15]), .Z(n32314) );
  XOR U36987 ( .A(n32320), .B(n32321), .Z(n31887) );
  ANDN U36988 ( .B(n32322), .A(n32323), .Z(n32320) );
  AND U36989 ( .A(a[59]), .B(b[14]), .Z(n32319) );
  XOR U36990 ( .A(n32325), .B(n32326), .Z(n31892) );
  ANDN U36991 ( .B(n32327), .A(n32328), .Z(n32325) );
  AND U36992 ( .A(a[60]), .B(b[13]), .Z(n32324) );
  XOR U36993 ( .A(n32330), .B(n32331), .Z(n31897) );
  ANDN U36994 ( .B(n32332), .A(n32333), .Z(n32330) );
  AND U36995 ( .A(a[61]), .B(b[12]), .Z(n32329) );
  XOR U36996 ( .A(n32335), .B(n32336), .Z(n31902) );
  ANDN U36997 ( .B(n32337), .A(n32338), .Z(n32335) );
  AND U36998 ( .A(a[62]), .B(b[11]), .Z(n32334) );
  XOR U36999 ( .A(n32340), .B(n32341), .Z(n31907) );
  ANDN U37000 ( .B(n32342), .A(n32343), .Z(n32340) );
  AND U37001 ( .A(a[63]), .B(b[10]), .Z(n32339) );
  XOR U37002 ( .A(n32345), .B(n32346), .Z(n31912) );
  ANDN U37003 ( .B(n32347), .A(n32348), .Z(n32345) );
  AND U37004 ( .A(b[9]), .B(a[64]), .Z(n32344) );
  XOR U37005 ( .A(n32350), .B(n32351), .Z(n31917) );
  ANDN U37006 ( .B(n32352), .A(n32353), .Z(n32350) );
  AND U37007 ( .A(b[8]), .B(a[65]), .Z(n32349) );
  XOR U37008 ( .A(n32355), .B(n32356), .Z(n31922) );
  ANDN U37009 ( .B(n32357), .A(n32358), .Z(n32355) );
  AND U37010 ( .A(b[7]), .B(a[66]), .Z(n32354) );
  XOR U37011 ( .A(n32360), .B(n32361), .Z(n31927) );
  ANDN U37012 ( .B(n32362), .A(n32363), .Z(n32360) );
  AND U37013 ( .A(b[6]), .B(a[67]), .Z(n32359) );
  XOR U37014 ( .A(n32365), .B(n32366), .Z(n31932) );
  ANDN U37015 ( .B(n32367), .A(n32368), .Z(n32365) );
  AND U37016 ( .A(b[5]), .B(a[68]), .Z(n32364) );
  XOR U37017 ( .A(n32370), .B(n32371), .Z(n31937) );
  ANDN U37018 ( .B(n32372), .A(n32373), .Z(n32370) );
  AND U37019 ( .A(b[4]), .B(a[69]), .Z(n32369) );
  XOR U37020 ( .A(n32375), .B(n32376), .Z(n31942) );
  ANDN U37021 ( .B(n31954), .A(n31955), .Z(n32375) );
  AND U37022 ( .A(b[2]), .B(a[70]), .Z(n32377) );
  XNOR U37023 ( .A(n32372), .B(n32376), .Z(n32378) );
  XOR U37024 ( .A(n32379), .B(n32380), .Z(n32376) );
  OR U37025 ( .A(n31957), .B(n31958), .Z(n32380) );
  XNOR U37026 ( .A(n32382), .B(n32383), .Z(n32381) );
  XOR U37027 ( .A(n32382), .B(n32385), .Z(n31957) );
  NAND U37028 ( .A(b[1]), .B(a[70]), .Z(n32385) );
  IV U37029 ( .A(n32379), .Z(n32382) );
  NANDN U37030 ( .A(n65), .B(n66), .Z(n32379) );
  XOR U37031 ( .A(n32386), .B(n32387), .Z(n66) );
  NAND U37032 ( .A(a[70]), .B(b[0]), .Z(n65) );
  XNOR U37033 ( .A(n32367), .B(n32371), .Z(n32388) );
  XNOR U37034 ( .A(n32362), .B(n32366), .Z(n32389) );
  XNOR U37035 ( .A(n32357), .B(n32361), .Z(n32390) );
  XNOR U37036 ( .A(n32352), .B(n32356), .Z(n32391) );
  XNOR U37037 ( .A(n32347), .B(n32351), .Z(n32392) );
  XNOR U37038 ( .A(n32342), .B(n32346), .Z(n32393) );
  XNOR U37039 ( .A(n32337), .B(n32341), .Z(n32394) );
  XNOR U37040 ( .A(n32332), .B(n32336), .Z(n32395) );
  XNOR U37041 ( .A(n32327), .B(n32331), .Z(n32396) );
  XNOR U37042 ( .A(n32322), .B(n32326), .Z(n32397) );
  XNOR U37043 ( .A(n32317), .B(n32321), .Z(n32398) );
  XNOR U37044 ( .A(n32312), .B(n32316), .Z(n32399) );
  XNOR U37045 ( .A(n32307), .B(n32311), .Z(n32400) );
  XNOR U37046 ( .A(n32302), .B(n32306), .Z(n32401) );
  XNOR U37047 ( .A(n32297), .B(n32301), .Z(n32402) );
  XNOR U37048 ( .A(n32292), .B(n32296), .Z(n32403) );
  XNOR U37049 ( .A(n32287), .B(n32291), .Z(n32404) );
  XNOR U37050 ( .A(n32282), .B(n32286), .Z(n32405) );
  XNOR U37051 ( .A(n32277), .B(n32281), .Z(n32406) );
  XNOR U37052 ( .A(n32272), .B(n32276), .Z(n32407) );
  XNOR U37053 ( .A(n32267), .B(n32271), .Z(n32408) );
  XNOR U37054 ( .A(n32262), .B(n32266), .Z(n32409) );
  XNOR U37055 ( .A(n32257), .B(n32261), .Z(n32410) );
  XNOR U37056 ( .A(n32252), .B(n32256), .Z(n32411) );
  XNOR U37057 ( .A(n32247), .B(n32251), .Z(n32412) );
  XNOR U37058 ( .A(n32242), .B(n32246), .Z(n32413) );
  XNOR U37059 ( .A(n32237), .B(n32241), .Z(n32414) );
  XNOR U37060 ( .A(n32232), .B(n32236), .Z(n32415) );
  XNOR U37061 ( .A(n32227), .B(n32231), .Z(n32416) );
  XNOR U37062 ( .A(n32222), .B(n32226), .Z(n32417) );
  XNOR U37063 ( .A(n32217), .B(n32221), .Z(n32418) );
  XNOR U37064 ( .A(n32212), .B(n32216), .Z(n32419) );
  XNOR U37065 ( .A(n32207), .B(n32211), .Z(n32420) );
  XNOR U37066 ( .A(n32202), .B(n32206), .Z(n32421) );
  XNOR U37067 ( .A(n32197), .B(n32201), .Z(n32422) );
  XNOR U37068 ( .A(n32192), .B(n32196), .Z(n32423) );
  XNOR U37069 ( .A(n32187), .B(n32191), .Z(n32424) );
  XNOR U37070 ( .A(n32182), .B(n32186), .Z(n32425) );
  XNOR U37071 ( .A(n32177), .B(n32181), .Z(n32426) );
  XNOR U37072 ( .A(n32172), .B(n32176), .Z(n32427) );
  XNOR U37073 ( .A(n32167), .B(n32171), .Z(n32428) );
  XNOR U37074 ( .A(n32162), .B(n32166), .Z(n32429) );
  XNOR U37075 ( .A(n32157), .B(n32161), .Z(n32430) );
  XNOR U37076 ( .A(n32152), .B(n32156), .Z(n32431) );
  XNOR U37077 ( .A(n32147), .B(n32151), .Z(n32432) );
  XNOR U37078 ( .A(n32142), .B(n32146), .Z(n32433) );
  XNOR U37079 ( .A(n32137), .B(n32141), .Z(n32434) );
  XNOR U37080 ( .A(n32132), .B(n32136), .Z(n32435) );
  XNOR U37081 ( .A(n32127), .B(n32131), .Z(n32436) );
  XNOR U37082 ( .A(n32122), .B(n32126), .Z(n32437) );
  XNOR U37083 ( .A(n32117), .B(n32121), .Z(n32438) );
  XNOR U37084 ( .A(n32112), .B(n32116), .Z(n32439) );
  XNOR U37085 ( .A(n32107), .B(n32111), .Z(n32440) );
  XNOR U37086 ( .A(n32102), .B(n32106), .Z(n32441) );
  XNOR U37087 ( .A(n32097), .B(n32101), .Z(n32442) );
  XNOR U37088 ( .A(n32092), .B(n32096), .Z(n32443) );
  XNOR U37089 ( .A(n32087), .B(n32091), .Z(n32444) );
  XNOR U37090 ( .A(n32082), .B(n32086), .Z(n32445) );
  XNOR U37091 ( .A(n32077), .B(n32081), .Z(n32446) );
  XNOR U37092 ( .A(n32072), .B(n32076), .Z(n32447) );
  XNOR U37093 ( .A(n32067), .B(n32071), .Z(n32448) );
  XNOR U37094 ( .A(n32062), .B(n32066), .Z(n32449) );
  XNOR U37095 ( .A(n32057), .B(n32061), .Z(n32450) );
  XNOR U37096 ( .A(n32052), .B(n32056), .Z(n32451) );
  XNOR U37097 ( .A(n32047), .B(n32051), .Z(n32452) );
  XNOR U37098 ( .A(n32042), .B(n32046), .Z(n32453) );
  XNOR U37099 ( .A(n32037), .B(n32041), .Z(n32454) );
  XNOR U37100 ( .A(n32032), .B(n32036), .Z(n32455) );
  XOR U37101 ( .A(n32456), .B(n32031), .Z(n32032) );
  AND U37102 ( .A(a[0]), .B(b[72]), .Z(n32456) );
  XNOR U37103 ( .A(n32457), .B(n32031), .Z(n32033) );
  XNOR U37104 ( .A(n32458), .B(n32459), .Z(n32031) );
  ANDN U37105 ( .B(n32460), .A(n32461), .Z(n32458) );
  AND U37106 ( .A(a[1]), .B(b[71]), .Z(n32457) );
  XOR U37107 ( .A(n32463), .B(n32464), .Z(n32036) );
  ANDN U37108 ( .B(n32465), .A(n32466), .Z(n32463) );
  AND U37109 ( .A(a[2]), .B(b[70]), .Z(n32462) );
  XOR U37110 ( .A(n32468), .B(n32469), .Z(n32041) );
  ANDN U37111 ( .B(n32470), .A(n32471), .Z(n32468) );
  AND U37112 ( .A(a[3]), .B(b[69]), .Z(n32467) );
  XOR U37113 ( .A(n32473), .B(n32474), .Z(n32046) );
  ANDN U37114 ( .B(n32475), .A(n32476), .Z(n32473) );
  AND U37115 ( .A(a[4]), .B(b[68]), .Z(n32472) );
  XOR U37116 ( .A(n32478), .B(n32479), .Z(n32051) );
  ANDN U37117 ( .B(n32480), .A(n32481), .Z(n32478) );
  AND U37118 ( .A(a[5]), .B(b[67]), .Z(n32477) );
  XOR U37119 ( .A(n32483), .B(n32484), .Z(n32056) );
  ANDN U37120 ( .B(n32485), .A(n32486), .Z(n32483) );
  AND U37121 ( .A(a[6]), .B(b[66]), .Z(n32482) );
  XOR U37122 ( .A(n32488), .B(n32489), .Z(n32061) );
  ANDN U37123 ( .B(n32490), .A(n32491), .Z(n32488) );
  AND U37124 ( .A(a[7]), .B(b[65]), .Z(n32487) );
  XOR U37125 ( .A(n32493), .B(n32494), .Z(n32066) );
  ANDN U37126 ( .B(n32495), .A(n32496), .Z(n32493) );
  AND U37127 ( .A(a[8]), .B(b[64]), .Z(n32492) );
  XOR U37128 ( .A(n32498), .B(n32499), .Z(n32071) );
  ANDN U37129 ( .B(n32500), .A(n32501), .Z(n32498) );
  AND U37130 ( .A(a[9]), .B(b[63]), .Z(n32497) );
  XOR U37131 ( .A(n32503), .B(n32504), .Z(n32076) );
  ANDN U37132 ( .B(n32505), .A(n32506), .Z(n32503) );
  AND U37133 ( .A(a[10]), .B(b[62]), .Z(n32502) );
  XOR U37134 ( .A(n32508), .B(n32509), .Z(n32081) );
  ANDN U37135 ( .B(n32510), .A(n32511), .Z(n32508) );
  AND U37136 ( .A(a[11]), .B(b[61]), .Z(n32507) );
  XOR U37137 ( .A(n32513), .B(n32514), .Z(n32086) );
  ANDN U37138 ( .B(n32515), .A(n32516), .Z(n32513) );
  AND U37139 ( .A(a[12]), .B(b[60]), .Z(n32512) );
  XOR U37140 ( .A(n32518), .B(n32519), .Z(n32091) );
  ANDN U37141 ( .B(n32520), .A(n32521), .Z(n32518) );
  AND U37142 ( .A(a[13]), .B(b[59]), .Z(n32517) );
  XOR U37143 ( .A(n32523), .B(n32524), .Z(n32096) );
  ANDN U37144 ( .B(n32525), .A(n32526), .Z(n32523) );
  AND U37145 ( .A(a[14]), .B(b[58]), .Z(n32522) );
  XOR U37146 ( .A(n32528), .B(n32529), .Z(n32101) );
  ANDN U37147 ( .B(n32530), .A(n32531), .Z(n32528) );
  AND U37148 ( .A(a[15]), .B(b[57]), .Z(n32527) );
  XOR U37149 ( .A(n32533), .B(n32534), .Z(n32106) );
  ANDN U37150 ( .B(n32535), .A(n32536), .Z(n32533) );
  AND U37151 ( .A(a[16]), .B(b[56]), .Z(n32532) );
  XOR U37152 ( .A(n32538), .B(n32539), .Z(n32111) );
  ANDN U37153 ( .B(n32540), .A(n32541), .Z(n32538) );
  AND U37154 ( .A(a[17]), .B(b[55]), .Z(n32537) );
  XOR U37155 ( .A(n32543), .B(n32544), .Z(n32116) );
  ANDN U37156 ( .B(n32545), .A(n32546), .Z(n32543) );
  AND U37157 ( .A(a[18]), .B(b[54]), .Z(n32542) );
  XOR U37158 ( .A(n32548), .B(n32549), .Z(n32121) );
  ANDN U37159 ( .B(n32550), .A(n32551), .Z(n32548) );
  AND U37160 ( .A(a[19]), .B(b[53]), .Z(n32547) );
  XOR U37161 ( .A(n32553), .B(n32554), .Z(n32126) );
  ANDN U37162 ( .B(n32555), .A(n32556), .Z(n32553) );
  AND U37163 ( .A(a[20]), .B(b[52]), .Z(n32552) );
  XOR U37164 ( .A(n32558), .B(n32559), .Z(n32131) );
  ANDN U37165 ( .B(n32560), .A(n32561), .Z(n32558) );
  AND U37166 ( .A(a[21]), .B(b[51]), .Z(n32557) );
  XOR U37167 ( .A(n32563), .B(n32564), .Z(n32136) );
  ANDN U37168 ( .B(n32565), .A(n32566), .Z(n32563) );
  AND U37169 ( .A(a[22]), .B(b[50]), .Z(n32562) );
  XOR U37170 ( .A(n32568), .B(n32569), .Z(n32141) );
  ANDN U37171 ( .B(n32570), .A(n32571), .Z(n32568) );
  AND U37172 ( .A(a[23]), .B(b[49]), .Z(n32567) );
  XOR U37173 ( .A(n32573), .B(n32574), .Z(n32146) );
  ANDN U37174 ( .B(n32575), .A(n32576), .Z(n32573) );
  AND U37175 ( .A(a[24]), .B(b[48]), .Z(n32572) );
  XOR U37176 ( .A(n32578), .B(n32579), .Z(n32151) );
  ANDN U37177 ( .B(n32580), .A(n32581), .Z(n32578) );
  AND U37178 ( .A(a[25]), .B(b[47]), .Z(n32577) );
  XOR U37179 ( .A(n32583), .B(n32584), .Z(n32156) );
  ANDN U37180 ( .B(n32585), .A(n32586), .Z(n32583) );
  AND U37181 ( .A(a[26]), .B(b[46]), .Z(n32582) );
  XOR U37182 ( .A(n32588), .B(n32589), .Z(n32161) );
  ANDN U37183 ( .B(n32590), .A(n32591), .Z(n32588) );
  AND U37184 ( .A(a[27]), .B(b[45]), .Z(n32587) );
  XOR U37185 ( .A(n32593), .B(n32594), .Z(n32166) );
  ANDN U37186 ( .B(n32595), .A(n32596), .Z(n32593) );
  AND U37187 ( .A(a[28]), .B(b[44]), .Z(n32592) );
  XOR U37188 ( .A(n32598), .B(n32599), .Z(n32171) );
  ANDN U37189 ( .B(n32600), .A(n32601), .Z(n32598) );
  AND U37190 ( .A(a[29]), .B(b[43]), .Z(n32597) );
  XOR U37191 ( .A(n32603), .B(n32604), .Z(n32176) );
  ANDN U37192 ( .B(n32605), .A(n32606), .Z(n32603) );
  AND U37193 ( .A(a[30]), .B(b[42]), .Z(n32602) );
  XOR U37194 ( .A(n32608), .B(n32609), .Z(n32181) );
  ANDN U37195 ( .B(n32610), .A(n32611), .Z(n32608) );
  AND U37196 ( .A(a[31]), .B(b[41]), .Z(n32607) );
  XOR U37197 ( .A(n32613), .B(n32614), .Z(n32186) );
  ANDN U37198 ( .B(n32615), .A(n32616), .Z(n32613) );
  AND U37199 ( .A(a[32]), .B(b[40]), .Z(n32612) );
  XOR U37200 ( .A(n32618), .B(n32619), .Z(n32191) );
  ANDN U37201 ( .B(n32620), .A(n32621), .Z(n32618) );
  AND U37202 ( .A(a[33]), .B(b[39]), .Z(n32617) );
  XOR U37203 ( .A(n32623), .B(n32624), .Z(n32196) );
  ANDN U37204 ( .B(n32625), .A(n32626), .Z(n32623) );
  AND U37205 ( .A(a[34]), .B(b[38]), .Z(n32622) );
  XOR U37206 ( .A(n32628), .B(n32629), .Z(n32201) );
  ANDN U37207 ( .B(n32630), .A(n32631), .Z(n32628) );
  AND U37208 ( .A(a[35]), .B(b[37]), .Z(n32627) );
  XOR U37209 ( .A(n32633), .B(n32634), .Z(n32206) );
  ANDN U37210 ( .B(n32635), .A(n32636), .Z(n32633) );
  AND U37211 ( .A(a[36]), .B(b[36]), .Z(n32632) );
  XOR U37212 ( .A(n32638), .B(n32639), .Z(n32211) );
  ANDN U37213 ( .B(n32640), .A(n32641), .Z(n32638) );
  AND U37214 ( .A(a[37]), .B(b[35]), .Z(n32637) );
  XOR U37215 ( .A(n32643), .B(n32644), .Z(n32216) );
  ANDN U37216 ( .B(n32645), .A(n32646), .Z(n32643) );
  AND U37217 ( .A(a[38]), .B(b[34]), .Z(n32642) );
  XOR U37218 ( .A(n32648), .B(n32649), .Z(n32221) );
  ANDN U37219 ( .B(n32650), .A(n32651), .Z(n32648) );
  AND U37220 ( .A(a[39]), .B(b[33]), .Z(n32647) );
  XOR U37221 ( .A(n32653), .B(n32654), .Z(n32226) );
  ANDN U37222 ( .B(n32655), .A(n32656), .Z(n32653) );
  AND U37223 ( .A(a[40]), .B(b[32]), .Z(n32652) );
  XOR U37224 ( .A(n32658), .B(n32659), .Z(n32231) );
  ANDN U37225 ( .B(n32660), .A(n32661), .Z(n32658) );
  AND U37226 ( .A(a[41]), .B(b[31]), .Z(n32657) );
  XOR U37227 ( .A(n32663), .B(n32664), .Z(n32236) );
  ANDN U37228 ( .B(n32665), .A(n32666), .Z(n32663) );
  AND U37229 ( .A(a[42]), .B(b[30]), .Z(n32662) );
  XOR U37230 ( .A(n32668), .B(n32669), .Z(n32241) );
  ANDN U37231 ( .B(n32670), .A(n32671), .Z(n32668) );
  AND U37232 ( .A(a[43]), .B(b[29]), .Z(n32667) );
  XOR U37233 ( .A(n32673), .B(n32674), .Z(n32246) );
  ANDN U37234 ( .B(n32675), .A(n32676), .Z(n32673) );
  AND U37235 ( .A(a[44]), .B(b[28]), .Z(n32672) );
  XOR U37236 ( .A(n32678), .B(n32679), .Z(n32251) );
  ANDN U37237 ( .B(n32680), .A(n32681), .Z(n32678) );
  AND U37238 ( .A(a[45]), .B(b[27]), .Z(n32677) );
  XOR U37239 ( .A(n32683), .B(n32684), .Z(n32256) );
  ANDN U37240 ( .B(n32685), .A(n32686), .Z(n32683) );
  AND U37241 ( .A(a[46]), .B(b[26]), .Z(n32682) );
  XOR U37242 ( .A(n32688), .B(n32689), .Z(n32261) );
  ANDN U37243 ( .B(n32690), .A(n32691), .Z(n32688) );
  AND U37244 ( .A(a[47]), .B(b[25]), .Z(n32687) );
  XOR U37245 ( .A(n32693), .B(n32694), .Z(n32266) );
  ANDN U37246 ( .B(n32695), .A(n32696), .Z(n32693) );
  AND U37247 ( .A(a[48]), .B(b[24]), .Z(n32692) );
  XOR U37248 ( .A(n32698), .B(n32699), .Z(n32271) );
  ANDN U37249 ( .B(n32700), .A(n32701), .Z(n32698) );
  AND U37250 ( .A(a[49]), .B(b[23]), .Z(n32697) );
  XOR U37251 ( .A(n32703), .B(n32704), .Z(n32276) );
  ANDN U37252 ( .B(n32705), .A(n32706), .Z(n32703) );
  AND U37253 ( .A(a[50]), .B(b[22]), .Z(n32702) );
  XOR U37254 ( .A(n32708), .B(n32709), .Z(n32281) );
  ANDN U37255 ( .B(n32710), .A(n32711), .Z(n32708) );
  AND U37256 ( .A(a[51]), .B(b[21]), .Z(n32707) );
  XOR U37257 ( .A(n32713), .B(n32714), .Z(n32286) );
  ANDN U37258 ( .B(n32715), .A(n32716), .Z(n32713) );
  AND U37259 ( .A(a[52]), .B(b[20]), .Z(n32712) );
  XOR U37260 ( .A(n32718), .B(n32719), .Z(n32291) );
  ANDN U37261 ( .B(n32720), .A(n32721), .Z(n32718) );
  AND U37262 ( .A(a[53]), .B(b[19]), .Z(n32717) );
  XOR U37263 ( .A(n32723), .B(n32724), .Z(n32296) );
  ANDN U37264 ( .B(n32725), .A(n32726), .Z(n32723) );
  AND U37265 ( .A(a[54]), .B(b[18]), .Z(n32722) );
  XOR U37266 ( .A(n32728), .B(n32729), .Z(n32301) );
  ANDN U37267 ( .B(n32730), .A(n32731), .Z(n32728) );
  AND U37268 ( .A(a[55]), .B(b[17]), .Z(n32727) );
  XOR U37269 ( .A(n32733), .B(n32734), .Z(n32306) );
  ANDN U37270 ( .B(n32735), .A(n32736), .Z(n32733) );
  AND U37271 ( .A(a[56]), .B(b[16]), .Z(n32732) );
  XOR U37272 ( .A(n32738), .B(n32739), .Z(n32311) );
  ANDN U37273 ( .B(n32740), .A(n32741), .Z(n32738) );
  AND U37274 ( .A(a[57]), .B(b[15]), .Z(n32737) );
  XOR U37275 ( .A(n32743), .B(n32744), .Z(n32316) );
  ANDN U37276 ( .B(n32745), .A(n32746), .Z(n32743) );
  AND U37277 ( .A(a[58]), .B(b[14]), .Z(n32742) );
  XOR U37278 ( .A(n32748), .B(n32749), .Z(n32321) );
  ANDN U37279 ( .B(n32750), .A(n32751), .Z(n32748) );
  AND U37280 ( .A(a[59]), .B(b[13]), .Z(n32747) );
  XOR U37281 ( .A(n32753), .B(n32754), .Z(n32326) );
  ANDN U37282 ( .B(n32755), .A(n32756), .Z(n32753) );
  AND U37283 ( .A(a[60]), .B(b[12]), .Z(n32752) );
  XOR U37284 ( .A(n32758), .B(n32759), .Z(n32331) );
  ANDN U37285 ( .B(n32760), .A(n32761), .Z(n32758) );
  AND U37286 ( .A(a[61]), .B(b[11]), .Z(n32757) );
  XOR U37287 ( .A(n32763), .B(n32764), .Z(n32336) );
  ANDN U37288 ( .B(n32765), .A(n32766), .Z(n32763) );
  AND U37289 ( .A(a[62]), .B(b[10]), .Z(n32762) );
  XOR U37290 ( .A(n32768), .B(n32769), .Z(n32341) );
  ANDN U37291 ( .B(n32770), .A(n32771), .Z(n32768) );
  AND U37292 ( .A(b[9]), .B(a[63]), .Z(n32767) );
  XOR U37293 ( .A(n32773), .B(n32774), .Z(n32346) );
  ANDN U37294 ( .B(n32775), .A(n32776), .Z(n32773) );
  AND U37295 ( .A(b[8]), .B(a[64]), .Z(n32772) );
  XOR U37296 ( .A(n32778), .B(n32779), .Z(n32351) );
  ANDN U37297 ( .B(n32780), .A(n32781), .Z(n32778) );
  AND U37298 ( .A(b[7]), .B(a[65]), .Z(n32777) );
  XOR U37299 ( .A(n32783), .B(n32784), .Z(n32356) );
  ANDN U37300 ( .B(n32785), .A(n32786), .Z(n32783) );
  AND U37301 ( .A(b[6]), .B(a[66]), .Z(n32782) );
  XOR U37302 ( .A(n32788), .B(n32789), .Z(n32361) );
  ANDN U37303 ( .B(n32790), .A(n32791), .Z(n32788) );
  AND U37304 ( .A(b[5]), .B(a[67]), .Z(n32787) );
  XOR U37305 ( .A(n32793), .B(n32794), .Z(n32366) );
  ANDN U37306 ( .B(n32795), .A(n32796), .Z(n32793) );
  AND U37307 ( .A(b[4]), .B(a[68]), .Z(n32792) );
  XOR U37308 ( .A(n32798), .B(n32799), .Z(n32371) );
  ANDN U37309 ( .B(n32383), .A(n32384), .Z(n32798) );
  AND U37310 ( .A(b[2]), .B(a[69]), .Z(n32800) );
  XNOR U37311 ( .A(n32795), .B(n32799), .Z(n32801) );
  XOR U37312 ( .A(n32802), .B(n32803), .Z(n32799) );
  OR U37313 ( .A(n32386), .B(n32387), .Z(n32803) );
  XNOR U37314 ( .A(n32805), .B(n32806), .Z(n32804) );
  XOR U37315 ( .A(n32805), .B(n32808), .Z(n32386) );
  NAND U37316 ( .A(b[1]), .B(a[69]), .Z(n32808) );
  IV U37317 ( .A(n32802), .Z(n32805) );
  NANDN U37318 ( .A(n69), .B(n70), .Z(n32802) );
  XOR U37319 ( .A(n32809), .B(n32810), .Z(n70) );
  NAND U37320 ( .A(a[69]), .B(b[0]), .Z(n69) );
  XNOR U37321 ( .A(n32790), .B(n32794), .Z(n32811) );
  XNOR U37322 ( .A(n32785), .B(n32789), .Z(n32812) );
  XNOR U37323 ( .A(n32780), .B(n32784), .Z(n32813) );
  XNOR U37324 ( .A(n32775), .B(n32779), .Z(n32814) );
  XNOR U37325 ( .A(n32770), .B(n32774), .Z(n32815) );
  XNOR U37326 ( .A(n32765), .B(n32769), .Z(n32816) );
  XNOR U37327 ( .A(n32760), .B(n32764), .Z(n32817) );
  XNOR U37328 ( .A(n32755), .B(n32759), .Z(n32818) );
  XNOR U37329 ( .A(n32750), .B(n32754), .Z(n32819) );
  XNOR U37330 ( .A(n32745), .B(n32749), .Z(n32820) );
  XNOR U37331 ( .A(n32740), .B(n32744), .Z(n32821) );
  XNOR U37332 ( .A(n32735), .B(n32739), .Z(n32822) );
  XNOR U37333 ( .A(n32730), .B(n32734), .Z(n32823) );
  XNOR U37334 ( .A(n32725), .B(n32729), .Z(n32824) );
  XNOR U37335 ( .A(n32720), .B(n32724), .Z(n32825) );
  XNOR U37336 ( .A(n32715), .B(n32719), .Z(n32826) );
  XNOR U37337 ( .A(n32710), .B(n32714), .Z(n32827) );
  XNOR U37338 ( .A(n32705), .B(n32709), .Z(n32828) );
  XNOR U37339 ( .A(n32700), .B(n32704), .Z(n32829) );
  XNOR U37340 ( .A(n32695), .B(n32699), .Z(n32830) );
  XNOR U37341 ( .A(n32690), .B(n32694), .Z(n32831) );
  XNOR U37342 ( .A(n32685), .B(n32689), .Z(n32832) );
  XNOR U37343 ( .A(n32680), .B(n32684), .Z(n32833) );
  XNOR U37344 ( .A(n32675), .B(n32679), .Z(n32834) );
  XNOR U37345 ( .A(n32670), .B(n32674), .Z(n32835) );
  XNOR U37346 ( .A(n32665), .B(n32669), .Z(n32836) );
  XNOR U37347 ( .A(n32660), .B(n32664), .Z(n32837) );
  XNOR U37348 ( .A(n32655), .B(n32659), .Z(n32838) );
  XNOR U37349 ( .A(n32650), .B(n32654), .Z(n32839) );
  XNOR U37350 ( .A(n32645), .B(n32649), .Z(n32840) );
  XNOR U37351 ( .A(n32640), .B(n32644), .Z(n32841) );
  XNOR U37352 ( .A(n32635), .B(n32639), .Z(n32842) );
  XNOR U37353 ( .A(n32630), .B(n32634), .Z(n32843) );
  XNOR U37354 ( .A(n32625), .B(n32629), .Z(n32844) );
  XNOR U37355 ( .A(n32620), .B(n32624), .Z(n32845) );
  XNOR U37356 ( .A(n32615), .B(n32619), .Z(n32846) );
  XNOR U37357 ( .A(n32610), .B(n32614), .Z(n32847) );
  XNOR U37358 ( .A(n32605), .B(n32609), .Z(n32848) );
  XNOR U37359 ( .A(n32600), .B(n32604), .Z(n32849) );
  XNOR U37360 ( .A(n32595), .B(n32599), .Z(n32850) );
  XNOR U37361 ( .A(n32590), .B(n32594), .Z(n32851) );
  XNOR U37362 ( .A(n32585), .B(n32589), .Z(n32852) );
  XNOR U37363 ( .A(n32580), .B(n32584), .Z(n32853) );
  XNOR U37364 ( .A(n32575), .B(n32579), .Z(n32854) );
  XNOR U37365 ( .A(n32570), .B(n32574), .Z(n32855) );
  XNOR U37366 ( .A(n32565), .B(n32569), .Z(n32856) );
  XNOR U37367 ( .A(n32560), .B(n32564), .Z(n32857) );
  XNOR U37368 ( .A(n32555), .B(n32559), .Z(n32858) );
  XNOR U37369 ( .A(n32550), .B(n32554), .Z(n32859) );
  XNOR U37370 ( .A(n32545), .B(n32549), .Z(n32860) );
  XNOR U37371 ( .A(n32540), .B(n32544), .Z(n32861) );
  XNOR U37372 ( .A(n32535), .B(n32539), .Z(n32862) );
  XNOR U37373 ( .A(n32530), .B(n32534), .Z(n32863) );
  XNOR U37374 ( .A(n32525), .B(n32529), .Z(n32864) );
  XNOR U37375 ( .A(n32520), .B(n32524), .Z(n32865) );
  XNOR U37376 ( .A(n32515), .B(n32519), .Z(n32866) );
  XNOR U37377 ( .A(n32510), .B(n32514), .Z(n32867) );
  XNOR U37378 ( .A(n32505), .B(n32509), .Z(n32868) );
  XNOR U37379 ( .A(n32500), .B(n32504), .Z(n32869) );
  XNOR U37380 ( .A(n32495), .B(n32499), .Z(n32870) );
  XNOR U37381 ( .A(n32490), .B(n32494), .Z(n32871) );
  XNOR U37382 ( .A(n32485), .B(n32489), .Z(n32872) );
  XNOR U37383 ( .A(n32480), .B(n32484), .Z(n32873) );
  XNOR U37384 ( .A(n32475), .B(n32479), .Z(n32874) );
  XNOR U37385 ( .A(n32470), .B(n32474), .Z(n32875) );
  XNOR U37386 ( .A(n32465), .B(n32469), .Z(n32876) );
  XNOR U37387 ( .A(n32460), .B(n32464), .Z(n32877) );
  XNOR U37388 ( .A(n32878), .B(n32459), .Z(n32460) );
  AND U37389 ( .A(a[0]), .B(b[71]), .Z(n32878) );
  XOR U37390 ( .A(n32879), .B(n32459), .Z(n32461) );
  XNOR U37391 ( .A(n32880), .B(n32881), .Z(n32459) );
  ANDN U37392 ( .B(n32882), .A(n32883), .Z(n32880) );
  AND U37393 ( .A(a[1]), .B(b[70]), .Z(n32879) );
  XOR U37394 ( .A(n32885), .B(n32886), .Z(n32464) );
  ANDN U37395 ( .B(n32887), .A(n32888), .Z(n32885) );
  AND U37396 ( .A(a[2]), .B(b[69]), .Z(n32884) );
  XOR U37397 ( .A(n32890), .B(n32891), .Z(n32469) );
  ANDN U37398 ( .B(n32892), .A(n32893), .Z(n32890) );
  AND U37399 ( .A(a[3]), .B(b[68]), .Z(n32889) );
  XOR U37400 ( .A(n32895), .B(n32896), .Z(n32474) );
  ANDN U37401 ( .B(n32897), .A(n32898), .Z(n32895) );
  AND U37402 ( .A(a[4]), .B(b[67]), .Z(n32894) );
  XOR U37403 ( .A(n32900), .B(n32901), .Z(n32479) );
  ANDN U37404 ( .B(n32902), .A(n32903), .Z(n32900) );
  AND U37405 ( .A(a[5]), .B(b[66]), .Z(n32899) );
  XOR U37406 ( .A(n32905), .B(n32906), .Z(n32484) );
  ANDN U37407 ( .B(n32907), .A(n32908), .Z(n32905) );
  AND U37408 ( .A(a[6]), .B(b[65]), .Z(n32904) );
  XOR U37409 ( .A(n32910), .B(n32911), .Z(n32489) );
  ANDN U37410 ( .B(n32912), .A(n32913), .Z(n32910) );
  AND U37411 ( .A(a[7]), .B(b[64]), .Z(n32909) );
  XOR U37412 ( .A(n32915), .B(n32916), .Z(n32494) );
  ANDN U37413 ( .B(n32917), .A(n32918), .Z(n32915) );
  AND U37414 ( .A(a[8]), .B(b[63]), .Z(n32914) );
  XOR U37415 ( .A(n32920), .B(n32921), .Z(n32499) );
  ANDN U37416 ( .B(n32922), .A(n32923), .Z(n32920) );
  AND U37417 ( .A(a[9]), .B(b[62]), .Z(n32919) );
  XOR U37418 ( .A(n32925), .B(n32926), .Z(n32504) );
  ANDN U37419 ( .B(n32927), .A(n32928), .Z(n32925) );
  AND U37420 ( .A(a[10]), .B(b[61]), .Z(n32924) );
  XOR U37421 ( .A(n32930), .B(n32931), .Z(n32509) );
  ANDN U37422 ( .B(n32932), .A(n32933), .Z(n32930) );
  AND U37423 ( .A(a[11]), .B(b[60]), .Z(n32929) );
  XOR U37424 ( .A(n32935), .B(n32936), .Z(n32514) );
  ANDN U37425 ( .B(n32937), .A(n32938), .Z(n32935) );
  AND U37426 ( .A(a[12]), .B(b[59]), .Z(n32934) );
  XOR U37427 ( .A(n32940), .B(n32941), .Z(n32519) );
  ANDN U37428 ( .B(n32942), .A(n32943), .Z(n32940) );
  AND U37429 ( .A(a[13]), .B(b[58]), .Z(n32939) );
  XOR U37430 ( .A(n32945), .B(n32946), .Z(n32524) );
  ANDN U37431 ( .B(n32947), .A(n32948), .Z(n32945) );
  AND U37432 ( .A(a[14]), .B(b[57]), .Z(n32944) );
  XOR U37433 ( .A(n32950), .B(n32951), .Z(n32529) );
  ANDN U37434 ( .B(n32952), .A(n32953), .Z(n32950) );
  AND U37435 ( .A(a[15]), .B(b[56]), .Z(n32949) );
  XOR U37436 ( .A(n32955), .B(n32956), .Z(n32534) );
  ANDN U37437 ( .B(n32957), .A(n32958), .Z(n32955) );
  AND U37438 ( .A(a[16]), .B(b[55]), .Z(n32954) );
  XOR U37439 ( .A(n32960), .B(n32961), .Z(n32539) );
  ANDN U37440 ( .B(n32962), .A(n32963), .Z(n32960) );
  AND U37441 ( .A(a[17]), .B(b[54]), .Z(n32959) );
  XOR U37442 ( .A(n32965), .B(n32966), .Z(n32544) );
  ANDN U37443 ( .B(n32967), .A(n32968), .Z(n32965) );
  AND U37444 ( .A(a[18]), .B(b[53]), .Z(n32964) );
  XOR U37445 ( .A(n32970), .B(n32971), .Z(n32549) );
  ANDN U37446 ( .B(n32972), .A(n32973), .Z(n32970) );
  AND U37447 ( .A(a[19]), .B(b[52]), .Z(n32969) );
  XOR U37448 ( .A(n32975), .B(n32976), .Z(n32554) );
  ANDN U37449 ( .B(n32977), .A(n32978), .Z(n32975) );
  AND U37450 ( .A(a[20]), .B(b[51]), .Z(n32974) );
  XOR U37451 ( .A(n32980), .B(n32981), .Z(n32559) );
  ANDN U37452 ( .B(n32982), .A(n32983), .Z(n32980) );
  AND U37453 ( .A(a[21]), .B(b[50]), .Z(n32979) );
  XOR U37454 ( .A(n32985), .B(n32986), .Z(n32564) );
  ANDN U37455 ( .B(n32987), .A(n32988), .Z(n32985) );
  AND U37456 ( .A(a[22]), .B(b[49]), .Z(n32984) );
  XOR U37457 ( .A(n32990), .B(n32991), .Z(n32569) );
  ANDN U37458 ( .B(n32992), .A(n32993), .Z(n32990) );
  AND U37459 ( .A(a[23]), .B(b[48]), .Z(n32989) );
  XOR U37460 ( .A(n32995), .B(n32996), .Z(n32574) );
  ANDN U37461 ( .B(n32997), .A(n32998), .Z(n32995) );
  AND U37462 ( .A(a[24]), .B(b[47]), .Z(n32994) );
  XOR U37463 ( .A(n33000), .B(n33001), .Z(n32579) );
  ANDN U37464 ( .B(n33002), .A(n33003), .Z(n33000) );
  AND U37465 ( .A(a[25]), .B(b[46]), .Z(n32999) );
  XOR U37466 ( .A(n33005), .B(n33006), .Z(n32584) );
  ANDN U37467 ( .B(n33007), .A(n33008), .Z(n33005) );
  AND U37468 ( .A(a[26]), .B(b[45]), .Z(n33004) );
  XOR U37469 ( .A(n33010), .B(n33011), .Z(n32589) );
  ANDN U37470 ( .B(n33012), .A(n33013), .Z(n33010) );
  AND U37471 ( .A(a[27]), .B(b[44]), .Z(n33009) );
  XOR U37472 ( .A(n33015), .B(n33016), .Z(n32594) );
  ANDN U37473 ( .B(n33017), .A(n33018), .Z(n33015) );
  AND U37474 ( .A(a[28]), .B(b[43]), .Z(n33014) );
  XOR U37475 ( .A(n33020), .B(n33021), .Z(n32599) );
  ANDN U37476 ( .B(n33022), .A(n33023), .Z(n33020) );
  AND U37477 ( .A(a[29]), .B(b[42]), .Z(n33019) );
  XOR U37478 ( .A(n33025), .B(n33026), .Z(n32604) );
  ANDN U37479 ( .B(n33027), .A(n33028), .Z(n33025) );
  AND U37480 ( .A(a[30]), .B(b[41]), .Z(n33024) );
  XOR U37481 ( .A(n33030), .B(n33031), .Z(n32609) );
  ANDN U37482 ( .B(n33032), .A(n33033), .Z(n33030) );
  AND U37483 ( .A(a[31]), .B(b[40]), .Z(n33029) );
  XOR U37484 ( .A(n33035), .B(n33036), .Z(n32614) );
  ANDN U37485 ( .B(n33037), .A(n33038), .Z(n33035) );
  AND U37486 ( .A(a[32]), .B(b[39]), .Z(n33034) );
  XOR U37487 ( .A(n33040), .B(n33041), .Z(n32619) );
  ANDN U37488 ( .B(n33042), .A(n33043), .Z(n33040) );
  AND U37489 ( .A(a[33]), .B(b[38]), .Z(n33039) );
  XOR U37490 ( .A(n33045), .B(n33046), .Z(n32624) );
  ANDN U37491 ( .B(n33047), .A(n33048), .Z(n33045) );
  AND U37492 ( .A(a[34]), .B(b[37]), .Z(n33044) );
  XOR U37493 ( .A(n33050), .B(n33051), .Z(n32629) );
  ANDN U37494 ( .B(n33052), .A(n33053), .Z(n33050) );
  AND U37495 ( .A(a[35]), .B(b[36]), .Z(n33049) );
  XOR U37496 ( .A(n33055), .B(n33056), .Z(n32634) );
  ANDN U37497 ( .B(n33057), .A(n33058), .Z(n33055) );
  AND U37498 ( .A(a[36]), .B(b[35]), .Z(n33054) );
  XOR U37499 ( .A(n33060), .B(n33061), .Z(n32639) );
  ANDN U37500 ( .B(n33062), .A(n33063), .Z(n33060) );
  AND U37501 ( .A(a[37]), .B(b[34]), .Z(n33059) );
  XOR U37502 ( .A(n33065), .B(n33066), .Z(n32644) );
  ANDN U37503 ( .B(n33067), .A(n33068), .Z(n33065) );
  AND U37504 ( .A(a[38]), .B(b[33]), .Z(n33064) );
  XOR U37505 ( .A(n33070), .B(n33071), .Z(n32649) );
  ANDN U37506 ( .B(n33072), .A(n33073), .Z(n33070) );
  AND U37507 ( .A(a[39]), .B(b[32]), .Z(n33069) );
  XOR U37508 ( .A(n33075), .B(n33076), .Z(n32654) );
  ANDN U37509 ( .B(n33077), .A(n33078), .Z(n33075) );
  AND U37510 ( .A(a[40]), .B(b[31]), .Z(n33074) );
  XOR U37511 ( .A(n33080), .B(n33081), .Z(n32659) );
  ANDN U37512 ( .B(n33082), .A(n33083), .Z(n33080) );
  AND U37513 ( .A(a[41]), .B(b[30]), .Z(n33079) );
  XOR U37514 ( .A(n33085), .B(n33086), .Z(n32664) );
  ANDN U37515 ( .B(n33087), .A(n33088), .Z(n33085) );
  AND U37516 ( .A(a[42]), .B(b[29]), .Z(n33084) );
  XOR U37517 ( .A(n33090), .B(n33091), .Z(n32669) );
  ANDN U37518 ( .B(n33092), .A(n33093), .Z(n33090) );
  AND U37519 ( .A(a[43]), .B(b[28]), .Z(n33089) );
  XOR U37520 ( .A(n33095), .B(n33096), .Z(n32674) );
  ANDN U37521 ( .B(n33097), .A(n33098), .Z(n33095) );
  AND U37522 ( .A(a[44]), .B(b[27]), .Z(n33094) );
  XOR U37523 ( .A(n33100), .B(n33101), .Z(n32679) );
  ANDN U37524 ( .B(n33102), .A(n33103), .Z(n33100) );
  AND U37525 ( .A(a[45]), .B(b[26]), .Z(n33099) );
  XOR U37526 ( .A(n33105), .B(n33106), .Z(n32684) );
  ANDN U37527 ( .B(n33107), .A(n33108), .Z(n33105) );
  AND U37528 ( .A(a[46]), .B(b[25]), .Z(n33104) );
  XOR U37529 ( .A(n33110), .B(n33111), .Z(n32689) );
  ANDN U37530 ( .B(n33112), .A(n33113), .Z(n33110) );
  AND U37531 ( .A(a[47]), .B(b[24]), .Z(n33109) );
  XOR U37532 ( .A(n33115), .B(n33116), .Z(n32694) );
  ANDN U37533 ( .B(n33117), .A(n33118), .Z(n33115) );
  AND U37534 ( .A(a[48]), .B(b[23]), .Z(n33114) );
  XOR U37535 ( .A(n33120), .B(n33121), .Z(n32699) );
  ANDN U37536 ( .B(n33122), .A(n33123), .Z(n33120) );
  AND U37537 ( .A(a[49]), .B(b[22]), .Z(n33119) );
  XOR U37538 ( .A(n33125), .B(n33126), .Z(n32704) );
  ANDN U37539 ( .B(n33127), .A(n33128), .Z(n33125) );
  AND U37540 ( .A(a[50]), .B(b[21]), .Z(n33124) );
  XOR U37541 ( .A(n33130), .B(n33131), .Z(n32709) );
  ANDN U37542 ( .B(n33132), .A(n33133), .Z(n33130) );
  AND U37543 ( .A(a[51]), .B(b[20]), .Z(n33129) );
  XOR U37544 ( .A(n33135), .B(n33136), .Z(n32714) );
  ANDN U37545 ( .B(n33137), .A(n33138), .Z(n33135) );
  AND U37546 ( .A(a[52]), .B(b[19]), .Z(n33134) );
  XOR U37547 ( .A(n33140), .B(n33141), .Z(n32719) );
  ANDN U37548 ( .B(n33142), .A(n33143), .Z(n33140) );
  AND U37549 ( .A(a[53]), .B(b[18]), .Z(n33139) );
  XOR U37550 ( .A(n33145), .B(n33146), .Z(n32724) );
  ANDN U37551 ( .B(n33147), .A(n33148), .Z(n33145) );
  AND U37552 ( .A(a[54]), .B(b[17]), .Z(n33144) );
  XOR U37553 ( .A(n33150), .B(n33151), .Z(n32729) );
  ANDN U37554 ( .B(n33152), .A(n33153), .Z(n33150) );
  AND U37555 ( .A(a[55]), .B(b[16]), .Z(n33149) );
  XOR U37556 ( .A(n33155), .B(n33156), .Z(n32734) );
  ANDN U37557 ( .B(n33157), .A(n33158), .Z(n33155) );
  AND U37558 ( .A(a[56]), .B(b[15]), .Z(n33154) );
  XOR U37559 ( .A(n33160), .B(n33161), .Z(n32739) );
  ANDN U37560 ( .B(n33162), .A(n33163), .Z(n33160) );
  AND U37561 ( .A(a[57]), .B(b[14]), .Z(n33159) );
  XOR U37562 ( .A(n33165), .B(n33166), .Z(n32744) );
  ANDN U37563 ( .B(n33167), .A(n33168), .Z(n33165) );
  AND U37564 ( .A(a[58]), .B(b[13]), .Z(n33164) );
  XOR U37565 ( .A(n33170), .B(n33171), .Z(n32749) );
  ANDN U37566 ( .B(n33172), .A(n33173), .Z(n33170) );
  AND U37567 ( .A(a[59]), .B(b[12]), .Z(n33169) );
  XOR U37568 ( .A(n33175), .B(n33176), .Z(n32754) );
  ANDN U37569 ( .B(n33177), .A(n33178), .Z(n33175) );
  AND U37570 ( .A(a[60]), .B(b[11]), .Z(n33174) );
  XOR U37571 ( .A(n33180), .B(n33181), .Z(n32759) );
  ANDN U37572 ( .B(n33182), .A(n33183), .Z(n33180) );
  AND U37573 ( .A(a[61]), .B(b[10]), .Z(n33179) );
  XOR U37574 ( .A(n33185), .B(n33186), .Z(n32764) );
  ANDN U37575 ( .B(n33187), .A(n33188), .Z(n33185) );
  AND U37576 ( .A(b[9]), .B(a[62]), .Z(n33184) );
  XOR U37577 ( .A(n33190), .B(n33191), .Z(n32769) );
  ANDN U37578 ( .B(n33192), .A(n33193), .Z(n33190) );
  AND U37579 ( .A(b[8]), .B(a[63]), .Z(n33189) );
  XOR U37580 ( .A(n33195), .B(n33196), .Z(n32774) );
  ANDN U37581 ( .B(n33197), .A(n33198), .Z(n33195) );
  AND U37582 ( .A(b[7]), .B(a[64]), .Z(n33194) );
  XOR U37583 ( .A(n33200), .B(n33201), .Z(n32779) );
  ANDN U37584 ( .B(n33202), .A(n33203), .Z(n33200) );
  AND U37585 ( .A(b[6]), .B(a[65]), .Z(n33199) );
  XOR U37586 ( .A(n33205), .B(n33206), .Z(n32784) );
  ANDN U37587 ( .B(n33207), .A(n33208), .Z(n33205) );
  AND U37588 ( .A(b[5]), .B(a[66]), .Z(n33204) );
  XOR U37589 ( .A(n33210), .B(n33211), .Z(n32789) );
  ANDN U37590 ( .B(n33212), .A(n33213), .Z(n33210) );
  AND U37591 ( .A(b[4]), .B(a[67]), .Z(n33209) );
  XOR U37592 ( .A(n33215), .B(n33216), .Z(n32794) );
  ANDN U37593 ( .B(n32806), .A(n32807), .Z(n33215) );
  AND U37594 ( .A(b[2]), .B(a[68]), .Z(n33217) );
  XNOR U37595 ( .A(n33212), .B(n33216), .Z(n33218) );
  XOR U37596 ( .A(n33219), .B(n33220), .Z(n33216) );
  OR U37597 ( .A(n32809), .B(n32810), .Z(n33220) );
  XNOR U37598 ( .A(n33222), .B(n33223), .Z(n33221) );
  XOR U37599 ( .A(n33222), .B(n33225), .Z(n32809) );
  NAND U37600 ( .A(b[1]), .B(a[68]), .Z(n33225) );
  IV U37601 ( .A(n33219), .Z(n33222) );
  NANDN U37602 ( .A(n71), .B(n72), .Z(n33219) );
  XOR U37603 ( .A(n33226), .B(n33227), .Z(n72) );
  NAND U37604 ( .A(a[68]), .B(b[0]), .Z(n71) );
  XNOR U37605 ( .A(n33207), .B(n33211), .Z(n33228) );
  XNOR U37606 ( .A(n33202), .B(n33206), .Z(n33229) );
  XNOR U37607 ( .A(n33197), .B(n33201), .Z(n33230) );
  XNOR U37608 ( .A(n33192), .B(n33196), .Z(n33231) );
  XNOR U37609 ( .A(n33187), .B(n33191), .Z(n33232) );
  XNOR U37610 ( .A(n33182), .B(n33186), .Z(n33233) );
  XNOR U37611 ( .A(n33177), .B(n33181), .Z(n33234) );
  XNOR U37612 ( .A(n33172), .B(n33176), .Z(n33235) );
  XNOR U37613 ( .A(n33167), .B(n33171), .Z(n33236) );
  XNOR U37614 ( .A(n33162), .B(n33166), .Z(n33237) );
  XNOR U37615 ( .A(n33157), .B(n33161), .Z(n33238) );
  XNOR U37616 ( .A(n33152), .B(n33156), .Z(n33239) );
  XNOR U37617 ( .A(n33147), .B(n33151), .Z(n33240) );
  XNOR U37618 ( .A(n33142), .B(n33146), .Z(n33241) );
  XNOR U37619 ( .A(n33137), .B(n33141), .Z(n33242) );
  XNOR U37620 ( .A(n33132), .B(n33136), .Z(n33243) );
  XNOR U37621 ( .A(n33127), .B(n33131), .Z(n33244) );
  XNOR U37622 ( .A(n33122), .B(n33126), .Z(n33245) );
  XNOR U37623 ( .A(n33117), .B(n33121), .Z(n33246) );
  XNOR U37624 ( .A(n33112), .B(n33116), .Z(n33247) );
  XNOR U37625 ( .A(n33107), .B(n33111), .Z(n33248) );
  XNOR U37626 ( .A(n33102), .B(n33106), .Z(n33249) );
  XNOR U37627 ( .A(n33097), .B(n33101), .Z(n33250) );
  XNOR U37628 ( .A(n33092), .B(n33096), .Z(n33251) );
  XNOR U37629 ( .A(n33087), .B(n33091), .Z(n33252) );
  XNOR U37630 ( .A(n33082), .B(n33086), .Z(n33253) );
  XNOR U37631 ( .A(n33077), .B(n33081), .Z(n33254) );
  XNOR U37632 ( .A(n33072), .B(n33076), .Z(n33255) );
  XNOR U37633 ( .A(n33067), .B(n33071), .Z(n33256) );
  XNOR U37634 ( .A(n33062), .B(n33066), .Z(n33257) );
  XNOR U37635 ( .A(n33057), .B(n33061), .Z(n33258) );
  XNOR U37636 ( .A(n33052), .B(n33056), .Z(n33259) );
  XNOR U37637 ( .A(n33047), .B(n33051), .Z(n33260) );
  XNOR U37638 ( .A(n33042), .B(n33046), .Z(n33261) );
  XNOR U37639 ( .A(n33037), .B(n33041), .Z(n33262) );
  XNOR U37640 ( .A(n33032), .B(n33036), .Z(n33263) );
  XNOR U37641 ( .A(n33027), .B(n33031), .Z(n33264) );
  XNOR U37642 ( .A(n33022), .B(n33026), .Z(n33265) );
  XNOR U37643 ( .A(n33017), .B(n33021), .Z(n33266) );
  XNOR U37644 ( .A(n33012), .B(n33016), .Z(n33267) );
  XNOR U37645 ( .A(n33007), .B(n33011), .Z(n33268) );
  XNOR U37646 ( .A(n33002), .B(n33006), .Z(n33269) );
  XNOR U37647 ( .A(n32997), .B(n33001), .Z(n33270) );
  XNOR U37648 ( .A(n32992), .B(n32996), .Z(n33271) );
  XNOR U37649 ( .A(n32987), .B(n32991), .Z(n33272) );
  XNOR U37650 ( .A(n32982), .B(n32986), .Z(n33273) );
  XNOR U37651 ( .A(n32977), .B(n32981), .Z(n33274) );
  XNOR U37652 ( .A(n32972), .B(n32976), .Z(n33275) );
  XNOR U37653 ( .A(n32967), .B(n32971), .Z(n33276) );
  XNOR U37654 ( .A(n32962), .B(n32966), .Z(n33277) );
  XNOR U37655 ( .A(n32957), .B(n32961), .Z(n33278) );
  XNOR U37656 ( .A(n32952), .B(n32956), .Z(n33279) );
  XNOR U37657 ( .A(n32947), .B(n32951), .Z(n33280) );
  XNOR U37658 ( .A(n32942), .B(n32946), .Z(n33281) );
  XNOR U37659 ( .A(n32937), .B(n32941), .Z(n33282) );
  XNOR U37660 ( .A(n32932), .B(n32936), .Z(n33283) );
  XNOR U37661 ( .A(n32927), .B(n32931), .Z(n33284) );
  XNOR U37662 ( .A(n32922), .B(n32926), .Z(n33285) );
  XNOR U37663 ( .A(n32917), .B(n32921), .Z(n33286) );
  XNOR U37664 ( .A(n32912), .B(n32916), .Z(n33287) );
  XNOR U37665 ( .A(n32907), .B(n32911), .Z(n33288) );
  XNOR U37666 ( .A(n32902), .B(n32906), .Z(n33289) );
  XNOR U37667 ( .A(n32897), .B(n32901), .Z(n33290) );
  XNOR U37668 ( .A(n32892), .B(n32896), .Z(n33291) );
  XNOR U37669 ( .A(n32887), .B(n32891), .Z(n33292) );
  XNOR U37670 ( .A(n32882), .B(n32886), .Z(n33293) );
  XOR U37671 ( .A(n33294), .B(n32881), .Z(n32882) );
  AND U37672 ( .A(a[0]), .B(b[70]), .Z(n33294) );
  XNOR U37673 ( .A(n33295), .B(n32881), .Z(n32883) );
  XNOR U37674 ( .A(n33296), .B(n33297), .Z(n32881) );
  ANDN U37675 ( .B(n33298), .A(n33299), .Z(n33296) );
  AND U37676 ( .A(a[1]), .B(b[69]), .Z(n33295) );
  XOR U37677 ( .A(n33301), .B(n33302), .Z(n32886) );
  ANDN U37678 ( .B(n33303), .A(n33304), .Z(n33301) );
  AND U37679 ( .A(a[2]), .B(b[68]), .Z(n33300) );
  XOR U37680 ( .A(n33306), .B(n33307), .Z(n32891) );
  ANDN U37681 ( .B(n33308), .A(n33309), .Z(n33306) );
  AND U37682 ( .A(a[3]), .B(b[67]), .Z(n33305) );
  XOR U37683 ( .A(n33311), .B(n33312), .Z(n32896) );
  ANDN U37684 ( .B(n33313), .A(n33314), .Z(n33311) );
  AND U37685 ( .A(a[4]), .B(b[66]), .Z(n33310) );
  XOR U37686 ( .A(n33316), .B(n33317), .Z(n32901) );
  ANDN U37687 ( .B(n33318), .A(n33319), .Z(n33316) );
  AND U37688 ( .A(a[5]), .B(b[65]), .Z(n33315) );
  XOR U37689 ( .A(n33321), .B(n33322), .Z(n32906) );
  ANDN U37690 ( .B(n33323), .A(n33324), .Z(n33321) );
  AND U37691 ( .A(a[6]), .B(b[64]), .Z(n33320) );
  XOR U37692 ( .A(n33326), .B(n33327), .Z(n32911) );
  ANDN U37693 ( .B(n33328), .A(n33329), .Z(n33326) );
  AND U37694 ( .A(a[7]), .B(b[63]), .Z(n33325) );
  XOR U37695 ( .A(n33331), .B(n33332), .Z(n32916) );
  ANDN U37696 ( .B(n33333), .A(n33334), .Z(n33331) );
  AND U37697 ( .A(a[8]), .B(b[62]), .Z(n33330) );
  XOR U37698 ( .A(n33336), .B(n33337), .Z(n32921) );
  ANDN U37699 ( .B(n33338), .A(n33339), .Z(n33336) );
  AND U37700 ( .A(a[9]), .B(b[61]), .Z(n33335) );
  XOR U37701 ( .A(n33341), .B(n33342), .Z(n32926) );
  ANDN U37702 ( .B(n33343), .A(n33344), .Z(n33341) );
  AND U37703 ( .A(a[10]), .B(b[60]), .Z(n33340) );
  XOR U37704 ( .A(n33346), .B(n33347), .Z(n32931) );
  ANDN U37705 ( .B(n33348), .A(n33349), .Z(n33346) );
  AND U37706 ( .A(a[11]), .B(b[59]), .Z(n33345) );
  XOR U37707 ( .A(n33351), .B(n33352), .Z(n32936) );
  ANDN U37708 ( .B(n33353), .A(n33354), .Z(n33351) );
  AND U37709 ( .A(a[12]), .B(b[58]), .Z(n33350) );
  XOR U37710 ( .A(n33356), .B(n33357), .Z(n32941) );
  ANDN U37711 ( .B(n33358), .A(n33359), .Z(n33356) );
  AND U37712 ( .A(a[13]), .B(b[57]), .Z(n33355) );
  XOR U37713 ( .A(n33361), .B(n33362), .Z(n32946) );
  ANDN U37714 ( .B(n33363), .A(n33364), .Z(n33361) );
  AND U37715 ( .A(a[14]), .B(b[56]), .Z(n33360) );
  XOR U37716 ( .A(n33366), .B(n33367), .Z(n32951) );
  ANDN U37717 ( .B(n33368), .A(n33369), .Z(n33366) );
  AND U37718 ( .A(a[15]), .B(b[55]), .Z(n33365) );
  XOR U37719 ( .A(n33371), .B(n33372), .Z(n32956) );
  ANDN U37720 ( .B(n33373), .A(n33374), .Z(n33371) );
  AND U37721 ( .A(a[16]), .B(b[54]), .Z(n33370) );
  XOR U37722 ( .A(n33376), .B(n33377), .Z(n32961) );
  ANDN U37723 ( .B(n33378), .A(n33379), .Z(n33376) );
  AND U37724 ( .A(a[17]), .B(b[53]), .Z(n33375) );
  XOR U37725 ( .A(n33381), .B(n33382), .Z(n32966) );
  ANDN U37726 ( .B(n33383), .A(n33384), .Z(n33381) );
  AND U37727 ( .A(a[18]), .B(b[52]), .Z(n33380) );
  XOR U37728 ( .A(n33386), .B(n33387), .Z(n32971) );
  ANDN U37729 ( .B(n33388), .A(n33389), .Z(n33386) );
  AND U37730 ( .A(a[19]), .B(b[51]), .Z(n33385) );
  XOR U37731 ( .A(n33391), .B(n33392), .Z(n32976) );
  ANDN U37732 ( .B(n33393), .A(n33394), .Z(n33391) );
  AND U37733 ( .A(a[20]), .B(b[50]), .Z(n33390) );
  XOR U37734 ( .A(n33396), .B(n33397), .Z(n32981) );
  ANDN U37735 ( .B(n33398), .A(n33399), .Z(n33396) );
  AND U37736 ( .A(a[21]), .B(b[49]), .Z(n33395) );
  XOR U37737 ( .A(n33401), .B(n33402), .Z(n32986) );
  ANDN U37738 ( .B(n33403), .A(n33404), .Z(n33401) );
  AND U37739 ( .A(a[22]), .B(b[48]), .Z(n33400) );
  XOR U37740 ( .A(n33406), .B(n33407), .Z(n32991) );
  ANDN U37741 ( .B(n33408), .A(n33409), .Z(n33406) );
  AND U37742 ( .A(a[23]), .B(b[47]), .Z(n33405) );
  XOR U37743 ( .A(n33411), .B(n33412), .Z(n32996) );
  ANDN U37744 ( .B(n33413), .A(n33414), .Z(n33411) );
  AND U37745 ( .A(a[24]), .B(b[46]), .Z(n33410) );
  XOR U37746 ( .A(n33416), .B(n33417), .Z(n33001) );
  ANDN U37747 ( .B(n33418), .A(n33419), .Z(n33416) );
  AND U37748 ( .A(a[25]), .B(b[45]), .Z(n33415) );
  XOR U37749 ( .A(n33421), .B(n33422), .Z(n33006) );
  ANDN U37750 ( .B(n33423), .A(n33424), .Z(n33421) );
  AND U37751 ( .A(a[26]), .B(b[44]), .Z(n33420) );
  XOR U37752 ( .A(n33426), .B(n33427), .Z(n33011) );
  ANDN U37753 ( .B(n33428), .A(n33429), .Z(n33426) );
  AND U37754 ( .A(a[27]), .B(b[43]), .Z(n33425) );
  XOR U37755 ( .A(n33431), .B(n33432), .Z(n33016) );
  ANDN U37756 ( .B(n33433), .A(n33434), .Z(n33431) );
  AND U37757 ( .A(a[28]), .B(b[42]), .Z(n33430) );
  XOR U37758 ( .A(n33436), .B(n33437), .Z(n33021) );
  ANDN U37759 ( .B(n33438), .A(n33439), .Z(n33436) );
  AND U37760 ( .A(a[29]), .B(b[41]), .Z(n33435) );
  XOR U37761 ( .A(n33441), .B(n33442), .Z(n33026) );
  ANDN U37762 ( .B(n33443), .A(n33444), .Z(n33441) );
  AND U37763 ( .A(a[30]), .B(b[40]), .Z(n33440) );
  XOR U37764 ( .A(n33446), .B(n33447), .Z(n33031) );
  ANDN U37765 ( .B(n33448), .A(n33449), .Z(n33446) );
  AND U37766 ( .A(a[31]), .B(b[39]), .Z(n33445) );
  XOR U37767 ( .A(n33451), .B(n33452), .Z(n33036) );
  ANDN U37768 ( .B(n33453), .A(n33454), .Z(n33451) );
  AND U37769 ( .A(a[32]), .B(b[38]), .Z(n33450) );
  XOR U37770 ( .A(n33456), .B(n33457), .Z(n33041) );
  ANDN U37771 ( .B(n33458), .A(n33459), .Z(n33456) );
  AND U37772 ( .A(a[33]), .B(b[37]), .Z(n33455) );
  XOR U37773 ( .A(n33461), .B(n33462), .Z(n33046) );
  ANDN U37774 ( .B(n33463), .A(n33464), .Z(n33461) );
  AND U37775 ( .A(a[34]), .B(b[36]), .Z(n33460) );
  XOR U37776 ( .A(n33466), .B(n33467), .Z(n33051) );
  ANDN U37777 ( .B(n33468), .A(n33469), .Z(n33466) );
  AND U37778 ( .A(a[35]), .B(b[35]), .Z(n33465) );
  XOR U37779 ( .A(n33471), .B(n33472), .Z(n33056) );
  ANDN U37780 ( .B(n33473), .A(n33474), .Z(n33471) );
  AND U37781 ( .A(a[36]), .B(b[34]), .Z(n33470) );
  XOR U37782 ( .A(n33476), .B(n33477), .Z(n33061) );
  ANDN U37783 ( .B(n33478), .A(n33479), .Z(n33476) );
  AND U37784 ( .A(a[37]), .B(b[33]), .Z(n33475) );
  XOR U37785 ( .A(n33481), .B(n33482), .Z(n33066) );
  ANDN U37786 ( .B(n33483), .A(n33484), .Z(n33481) );
  AND U37787 ( .A(a[38]), .B(b[32]), .Z(n33480) );
  XOR U37788 ( .A(n33486), .B(n33487), .Z(n33071) );
  ANDN U37789 ( .B(n33488), .A(n33489), .Z(n33486) );
  AND U37790 ( .A(a[39]), .B(b[31]), .Z(n33485) );
  XOR U37791 ( .A(n33491), .B(n33492), .Z(n33076) );
  ANDN U37792 ( .B(n33493), .A(n33494), .Z(n33491) );
  AND U37793 ( .A(a[40]), .B(b[30]), .Z(n33490) );
  XOR U37794 ( .A(n33496), .B(n33497), .Z(n33081) );
  ANDN U37795 ( .B(n33498), .A(n33499), .Z(n33496) );
  AND U37796 ( .A(a[41]), .B(b[29]), .Z(n33495) );
  XOR U37797 ( .A(n33501), .B(n33502), .Z(n33086) );
  ANDN U37798 ( .B(n33503), .A(n33504), .Z(n33501) );
  AND U37799 ( .A(a[42]), .B(b[28]), .Z(n33500) );
  XOR U37800 ( .A(n33506), .B(n33507), .Z(n33091) );
  ANDN U37801 ( .B(n33508), .A(n33509), .Z(n33506) );
  AND U37802 ( .A(a[43]), .B(b[27]), .Z(n33505) );
  XOR U37803 ( .A(n33511), .B(n33512), .Z(n33096) );
  ANDN U37804 ( .B(n33513), .A(n33514), .Z(n33511) );
  AND U37805 ( .A(a[44]), .B(b[26]), .Z(n33510) );
  XOR U37806 ( .A(n33516), .B(n33517), .Z(n33101) );
  ANDN U37807 ( .B(n33518), .A(n33519), .Z(n33516) );
  AND U37808 ( .A(a[45]), .B(b[25]), .Z(n33515) );
  XOR U37809 ( .A(n33521), .B(n33522), .Z(n33106) );
  ANDN U37810 ( .B(n33523), .A(n33524), .Z(n33521) );
  AND U37811 ( .A(a[46]), .B(b[24]), .Z(n33520) );
  XOR U37812 ( .A(n33526), .B(n33527), .Z(n33111) );
  ANDN U37813 ( .B(n33528), .A(n33529), .Z(n33526) );
  AND U37814 ( .A(a[47]), .B(b[23]), .Z(n33525) );
  XOR U37815 ( .A(n33531), .B(n33532), .Z(n33116) );
  ANDN U37816 ( .B(n33533), .A(n33534), .Z(n33531) );
  AND U37817 ( .A(a[48]), .B(b[22]), .Z(n33530) );
  XOR U37818 ( .A(n33536), .B(n33537), .Z(n33121) );
  ANDN U37819 ( .B(n33538), .A(n33539), .Z(n33536) );
  AND U37820 ( .A(a[49]), .B(b[21]), .Z(n33535) );
  XOR U37821 ( .A(n33541), .B(n33542), .Z(n33126) );
  ANDN U37822 ( .B(n33543), .A(n33544), .Z(n33541) );
  AND U37823 ( .A(a[50]), .B(b[20]), .Z(n33540) );
  XOR U37824 ( .A(n33546), .B(n33547), .Z(n33131) );
  ANDN U37825 ( .B(n33548), .A(n33549), .Z(n33546) );
  AND U37826 ( .A(a[51]), .B(b[19]), .Z(n33545) );
  XOR U37827 ( .A(n33551), .B(n33552), .Z(n33136) );
  ANDN U37828 ( .B(n33553), .A(n33554), .Z(n33551) );
  AND U37829 ( .A(a[52]), .B(b[18]), .Z(n33550) );
  XOR U37830 ( .A(n33556), .B(n33557), .Z(n33141) );
  ANDN U37831 ( .B(n33558), .A(n33559), .Z(n33556) );
  AND U37832 ( .A(a[53]), .B(b[17]), .Z(n33555) );
  XOR U37833 ( .A(n33561), .B(n33562), .Z(n33146) );
  ANDN U37834 ( .B(n33563), .A(n33564), .Z(n33561) );
  AND U37835 ( .A(a[54]), .B(b[16]), .Z(n33560) );
  XOR U37836 ( .A(n33566), .B(n33567), .Z(n33151) );
  ANDN U37837 ( .B(n33568), .A(n33569), .Z(n33566) );
  AND U37838 ( .A(a[55]), .B(b[15]), .Z(n33565) );
  XOR U37839 ( .A(n33571), .B(n33572), .Z(n33156) );
  ANDN U37840 ( .B(n33573), .A(n33574), .Z(n33571) );
  AND U37841 ( .A(a[56]), .B(b[14]), .Z(n33570) );
  XOR U37842 ( .A(n33576), .B(n33577), .Z(n33161) );
  ANDN U37843 ( .B(n33578), .A(n33579), .Z(n33576) );
  AND U37844 ( .A(a[57]), .B(b[13]), .Z(n33575) );
  XOR U37845 ( .A(n33581), .B(n33582), .Z(n33166) );
  ANDN U37846 ( .B(n33583), .A(n33584), .Z(n33581) );
  AND U37847 ( .A(a[58]), .B(b[12]), .Z(n33580) );
  XOR U37848 ( .A(n33586), .B(n33587), .Z(n33171) );
  ANDN U37849 ( .B(n33588), .A(n33589), .Z(n33586) );
  AND U37850 ( .A(a[59]), .B(b[11]), .Z(n33585) );
  XOR U37851 ( .A(n33591), .B(n33592), .Z(n33176) );
  ANDN U37852 ( .B(n33593), .A(n33594), .Z(n33591) );
  AND U37853 ( .A(a[60]), .B(b[10]), .Z(n33590) );
  XOR U37854 ( .A(n33596), .B(n33597), .Z(n33181) );
  ANDN U37855 ( .B(n33598), .A(n33599), .Z(n33596) );
  AND U37856 ( .A(b[9]), .B(a[61]), .Z(n33595) );
  XOR U37857 ( .A(n33601), .B(n33602), .Z(n33186) );
  ANDN U37858 ( .B(n33603), .A(n33604), .Z(n33601) );
  AND U37859 ( .A(b[8]), .B(a[62]), .Z(n33600) );
  XOR U37860 ( .A(n33606), .B(n33607), .Z(n33191) );
  ANDN U37861 ( .B(n33608), .A(n33609), .Z(n33606) );
  AND U37862 ( .A(b[7]), .B(a[63]), .Z(n33605) );
  XOR U37863 ( .A(n33611), .B(n33612), .Z(n33196) );
  ANDN U37864 ( .B(n33613), .A(n33614), .Z(n33611) );
  AND U37865 ( .A(b[6]), .B(a[64]), .Z(n33610) );
  XOR U37866 ( .A(n33616), .B(n33617), .Z(n33201) );
  ANDN U37867 ( .B(n33618), .A(n33619), .Z(n33616) );
  AND U37868 ( .A(b[5]), .B(a[65]), .Z(n33615) );
  XOR U37869 ( .A(n33621), .B(n33622), .Z(n33206) );
  ANDN U37870 ( .B(n33623), .A(n33624), .Z(n33621) );
  AND U37871 ( .A(b[4]), .B(a[66]), .Z(n33620) );
  XOR U37872 ( .A(n33626), .B(n33627), .Z(n33211) );
  ANDN U37873 ( .B(n33223), .A(n33224), .Z(n33626) );
  AND U37874 ( .A(b[2]), .B(a[67]), .Z(n33628) );
  XNOR U37875 ( .A(n33623), .B(n33627), .Z(n33629) );
  XOR U37876 ( .A(n33630), .B(n33631), .Z(n33627) );
  OR U37877 ( .A(n33226), .B(n33227), .Z(n33631) );
  XNOR U37878 ( .A(n33633), .B(n33634), .Z(n33632) );
  XOR U37879 ( .A(n33633), .B(n33636), .Z(n33226) );
  NAND U37880 ( .A(b[1]), .B(a[67]), .Z(n33636) );
  IV U37881 ( .A(n33630), .Z(n33633) );
  NANDN U37882 ( .A(n73), .B(n74), .Z(n33630) );
  XOR U37883 ( .A(n33637), .B(n33638), .Z(n74) );
  NAND U37884 ( .A(a[67]), .B(b[0]), .Z(n73) );
  XNOR U37885 ( .A(n33618), .B(n33622), .Z(n33639) );
  XNOR U37886 ( .A(n33613), .B(n33617), .Z(n33640) );
  XNOR U37887 ( .A(n33608), .B(n33612), .Z(n33641) );
  XNOR U37888 ( .A(n33603), .B(n33607), .Z(n33642) );
  XNOR U37889 ( .A(n33598), .B(n33602), .Z(n33643) );
  XNOR U37890 ( .A(n33593), .B(n33597), .Z(n33644) );
  XNOR U37891 ( .A(n33588), .B(n33592), .Z(n33645) );
  XNOR U37892 ( .A(n33583), .B(n33587), .Z(n33646) );
  XNOR U37893 ( .A(n33578), .B(n33582), .Z(n33647) );
  XNOR U37894 ( .A(n33573), .B(n33577), .Z(n33648) );
  XNOR U37895 ( .A(n33568), .B(n33572), .Z(n33649) );
  XNOR U37896 ( .A(n33563), .B(n33567), .Z(n33650) );
  XNOR U37897 ( .A(n33558), .B(n33562), .Z(n33651) );
  XNOR U37898 ( .A(n33553), .B(n33557), .Z(n33652) );
  XNOR U37899 ( .A(n33548), .B(n33552), .Z(n33653) );
  XNOR U37900 ( .A(n33543), .B(n33547), .Z(n33654) );
  XNOR U37901 ( .A(n33538), .B(n33542), .Z(n33655) );
  XNOR U37902 ( .A(n33533), .B(n33537), .Z(n33656) );
  XNOR U37903 ( .A(n33528), .B(n33532), .Z(n33657) );
  XNOR U37904 ( .A(n33523), .B(n33527), .Z(n33658) );
  XNOR U37905 ( .A(n33518), .B(n33522), .Z(n33659) );
  XNOR U37906 ( .A(n33513), .B(n33517), .Z(n33660) );
  XNOR U37907 ( .A(n33508), .B(n33512), .Z(n33661) );
  XNOR U37908 ( .A(n33503), .B(n33507), .Z(n33662) );
  XNOR U37909 ( .A(n33498), .B(n33502), .Z(n33663) );
  XNOR U37910 ( .A(n33493), .B(n33497), .Z(n33664) );
  XNOR U37911 ( .A(n33488), .B(n33492), .Z(n33665) );
  XNOR U37912 ( .A(n33483), .B(n33487), .Z(n33666) );
  XNOR U37913 ( .A(n33478), .B(n33482), .Z(n33667) );
  XNOR U37914 ( .A(n33473), .B(n33477), .Z(n33668) );
  XNOR U37915 ( .A(n33468), .B(n33472), .Z(n33669) );
  XNOR U37916 ( .A(n33463), .B(n33467), .Z(n33670) );
  XNOR U37917 ( .A(n33458), .B(n33462), .Z(n33671) );
  XNOR U37918 ( .A(n33453), .B(n33457), .Z(n33672) );
  XNOR U37919 ( .A(n33448), .B(n33452), .Z(n33673) );
  XNOR U37920 ( .A(n33443), .B(n33447), .Z(n33674) );
  XNOR U37921 ( .A(n33438), .B(n33442), .Z(n33675) );
  XNOR U37922 ( .A(n33433), .B(n33437), .Z(n33676) );
  XNOR U37923 ( .A(n33428), .B(n33432), .Z(n33677) );
  XNOR U37924 ( .A(n33423), .B(n33427), .Z(n33678) );
  XNOR U37925 ( .A(n33418), .B(n33422), .Z(n33679) );
  XNOR U37926 ( .A(n33413), .B(n33417), .Z(n33680) );
  XNOR U37927 ( .A(n33408), .B(n33412), .Z(n33681) );
  XNOR U37928 ( .A(n33403), .B(n33407), .Z(n33682) );
  XNOR U37929 ( .A(n33398), .B(n33402), .Z(n33683) );
  XNOR U37930 ( .A(n33393), .B(n33397), .Z(n33684) );
  XNOR U37931 ( .A(n33388), .B(n33392), .Z(n33685) );
  XNOR U37932 ( .A(n33383), .B(n33387), .Z(n33686) );
  XNOR U37933 ( .A(n33378), .B(n33382), .Z(n33687) );
  XNOR U37934 ( .A(n33373), .B(n33377), .Z(n33688) );
  XNOR U37935 ( .A(n33368), .B(n33372), .Z(n33689) );
  XNOR U37936 ( .A(n33363), .B(n33367), .Z(n33690) );
  XNOR U37937 ( .A(n33358), .B(n33362), .Z(n33691) );
  XNOR U37938 ( .A(n33353), .B(n33357), .Z(n33692) );
  XNOR U37939 ( .A(n33348), .B(n33352), .Z(n33693) );
  XNOR U37940 ( .A(n33343), .B(n33347), .Z(n33694) );
  XNOR U37941 ( .A(n33338), .B(n33342), .Z(n33695) );
  XNOR U37942 ( .A(n33333), .B(n33337), .Z(n33696) );
  XNOR U37943 ( .A(n33328), .B(n33332), .Z(n33697) );
  XNOR U37944 ( .A(n33323), .B(n33327), .Z(n33698) );
  XNOR U37945 ( .A(n33318), .B(n33322), .Z(n33699) );
  XNOR U37946 ( .A(n33313), .B(n33317), .Z(n33700) );
  XNOR U37947 ( .A(n33308), .B(n33312), .Z(n33701) );
  XNOR U37948 ( .A(n33303), .B(n33307), .Z(n33702) );
  XNOR U37949 ( .A(n33298), .B(n33302), .Z(n33703) );
  XNOR U37950 ( .A(n33704), .B(n33297), .Z(n33298) );
  AND U37951 ( .A(a[0]), .B(b[69]), .Z(n33704) );
  XOR U37952 ( .A(n33705), .B(n33297), .Z(n33299) );
  XNOR U37953 ( .A(n33706), .B(n33707), .Z(n33297) );
  ANDN U37954 ( .B(n33708), .A(n33709), .Z(n33706) );
  AND U37955 ( .A(a[1]), .B(b[68]), .Z(n33705) );
  XOR U37956 ( .A(n33711), .B(n33712), .Z(n33302) );
  ANDN U37957 ( .B(n33713), .A(n33714), .Z(n33711) );
  AND U37958 ( .A(a[2]), .B(b[67]), .Z(n33710) );
  XOR U37959 ( .A(n33716), .B(n33717), .Z(n33307) );
  ANDN U37960 ( .B(n33718), .A(n33719), .Z(n33716) );
  AND U37961 ( .A(a[3]), .B(b[66]), .Z(n33715) );
  XOR U37962 ( .A(n33721), .B(n33722), .Z(n33312) );
  ANDN U37963 ( .B(n33723), .A(n33724), .Z(n33721) );
  AND U37964 ( .A(a[4]), .B(b[65]), .Z(n33720) );
  XOR U37965 ( .A(n33726), .B(n33727), .Z(n33317) );
  ANDN U37966 ( .B(n33728), .A(n33729), .Z(n33726) );
  AND U37967 ( .A(a[5]), .B(b[64]), .Z(n33725) );
  XOR U37968 ( .A(n33731), .B(n33732), .Z(n33322) );
  ANDN U37969 ( .B(n33733), .A(n33734), .Z(n33731) );
  AND U37970 ( .A(a[6]), .B(b[63]), .Z(n33730) );
  XOR U37971 ( .A(n33736), .B(n33737), .Z(n33327) );
  ANDN U37972 ( .B(n33738), .A(n33739), .Z(n33736) );
  AND U37973 ( .A(a[7]), .B(b[62]), .Z(n33735) );
  XOR U37974 ( .A(n33741), .B(n33742), .Z(n33332) );
  ANDN U37975 ( .B(n33743), .A(n33744), .Z(n33741) );
  AND U37976 ( .A(a[8]), .B(b[61]), .Z(n33740) );
  XOR U37977 ( .A(n33746), .B(n33747), .Z(n33337) );
  ANDN U37978 ( .B(n33748), .A(n33749), .Z(n33746) );
  AND U37979 ( .A(a[9]), .B(b[60]), .Z(n33745) );
  XOR U37980 ( .A(n33751), .B(n33752), .Z(n33342) );
  ANDN U37981 ( .B(n33753), .A(n33754), .Z(n33751) );
  AND U37982 ( .A(a[10]), .B(b[59]), .Z(n33750) );
  XOR U37983 ( .A(n33756), .B(n33757), .Z(n33347) );
  ANDN U37984 ( .B(n33758), .A(n33759), .Z(n33756) );
  AND U37985 ( .A(a[11]), .B(b[58]), .Z(n33755) );
  XOR U37986 ( .A(n33761), .B(n33762), .Z(n33352) );
  ANDN U37987 ( .B(n33763), .A(n33764), .Z(n33761) );
  AND U37988 ( .A(a[12]), .B(b[57]), .Z(n33760) );
  XOR U37989 ( .A(n33766), .B(n33767), .Z(n33357) );
  ANDN U37990 ( .B(n33768), .A(n33769), .Z(n33766) );
  AND U37991 ( .A(a[13]), .B(b[56]), .Z(n33765) );
  XOR U37992 ( .A(n33771), .B(n33772), .Z(n33362) );
  ANDN U37993 ( .B(n33773), .A(n33774), .Z(n33771) );
  AND U37994 ( .A(a[14]), .B(b[55]), .Z(n33770) );
  XOR U37995 ( .A(n33776), .B(n33777), .Z(n33367) );
  ANDN U37996 ( .B(n33778), .A(n33779), .Z(n33776) );
  AND U37997 ( .A(a[15]), .B(b[54]), .Z(n33775) );
  XOR U37998 ( .A(n33781), .B(n33782), .Z(n33372) );
  ANDN U37999 ( .B(n33783), .A(n33784), .Z(n33781) );
  AND U38000 ( .A(a[16]), .B(b[53]), .Z(n33780) );
  XOR U38001 ( .A(n33786), .B(n33787), .Z(n33377) );
  ANDN U38002 ( .B(n33788), .A(n33789), .Z(n33786) );
  AND U38003 ( .A(a[17]), .B(b[52]), .Z(n33785) );
  XOR U38004 ( .A(n33791), .B(n33792), .Z(n33382) );
  ANDN U38005 ( .B(n33793), .A(n33794), .Z(n33791) );
  AND U38006 ( .A(a[18]), .B(b[51]), .Z(n33790) );
  XOR U38007 ( .A(n33796), .B(n33797), .Z(n33387) );
  ANDN U38008 ( .B(n33798), .A(n33799), .Z(n33796) );
  AND U38009 ( .A(a[19]), .B(b[50]), .Z(n33795) );
  XOR U38010 ( .A(n33801), .B(n33802), .Z(n33392) );
  ANDN U38011 ( .B(n33803), .A(n33804), .Z(n33801) );
  AND U38012 ( .A(a[20]), .B(b[49]), .Z(n33800) );
  XOR U38013 ( .A(n33806), .B(n33807), .Z(n33397) );
  ANDN U38014 ( .B(n33808), .A(n33809), .Z(n33806) );
  AND U38015 ( .A(a[21]), .B(b[48]), .Z(n33805) );
  XOR U38016 ( .A(n33811), .B(n33812), .Z(n33402) );
  ANDN U38017 ( .B(n33813), .A(n33814), .Z(n33811) );
  AND U38018 ( .A(a[22]), .B(b[47]), .Z(n33810) );
  XOR U38019 ( .A(n33816), .B(n33817), .Z(n33407) );
  ANDN U38020 ( .B(n33818), .A(n33819), .Z(n33816) );
  AND U38021 ( .A(a[23]), .B(b[46]), .Z(n33815) );
  XOR U38022 ( .A(n33821), .B(n33822), .Z(n33412) );
  ANDN U38023 ( .B(n33823), .A(n33824), .Z(n33821) );
  AND U38024 ( .A(a[24]), .B(b[45]), .Z(n33820) );
  XOR U38025 ( .A(n33826), .B(n33827), .Z(n33417) );
  ANDN U38026 ( .B(n33828), .A(n33829), .Z(n33826) );
  AND U38027 ( .A(a[25]), .B(b[44]), .Z(n33825) );
  XOR U38028 ( .A(n33831), .B(n33832), .Z(n33422) );
  ANDN U38029 ( .B(n33833), .A(n33834), .Z(n33831) );
  AND U38030 ( .A(a[26]), .B(b[43]), .Z(n33830) );
  XOR U38031 ( .A(n33836), .B(n33837), .Z(n33427) );
  ANDN U38032 ( .B(n33838), .A(n33839), .Z(n33836) );
  AND U38033 ( .A(a[27]), .B(b[42]), .Z(n33835) );
  XOR U38034 ( .A(n33841), .B(n33842), .Z(n33432) );
  ANDN U38035 ( .B(n33843), .A(n33844), .Z(n33841) );
  AND U38036 ( .A(a[28]), .B(b[41]), .Z(n33840) );
  XOR U38037 ( .A(n33846), .B(n33847), .Z(n33437) );
  ANDN U38038 ( .B(n33848), .A(n33849), .Z(n33846) );
  AND U38039 ( .A(a[29]), .B(b[40]), .Z(n33845) );
  XOR U38040 ( .A(n33851), .B(n33852), .Z(n33442) );
  ANDN U38041 ( .B(n33853), .A(n33854), .Z(n33851) );
  AND U38042 ( .A(a[30]), .B(b[39]), .Z(n33850) );
  XOR U38043 ( .A(n33856), .B(n33857), .Z(n33447) );
  ANDN U38044 ( .B(n33858), .A(n33859), .Z(n33856) );
  AND U38045 ( .A(a[31]), .B(b[38]), .Z(n33855) );
  XOR U38046 ( .A(n33861), .B(n33862), .Z(n33452) );
  ANDN U38047 ( .B(n33863), .A(n33864), .Z(n33861) );
  AND U38048 ( .A(a[32]), .B(b[37]), .Z(n33860) );
  XOR U38049 ( .A(n33866), .B(n33867), .Z(n33457) );
  ANDN U38050 ( .B(n33868), .A(n33869), .Z(n33866) );
  AND U38051 ( .A(a[33]), .B(b[36]), .Z(n33865) );
  XOR U38052 ( .A(n33871), .B(n33872), .Z(n33462) );
  ANDN U38053 ( .B(n33873), .A(n33874), .Z(n33871) );
  AND U38054 ( .A(a[34]), .B(b[35]), .Z(n33870) );
  XOR U38055 ( .A(n33876), .B(n33877), .Z(n33467) );
  ANDN U38056 ( .B(n33878), .A(n33879), .Z(n33876) );
  AND U38057 ( .A(a[35]), .B(b[34]), .Z(n33875) );
  XOR U38058 ( .A(n33881), .B(n33882), .Z(n33472) );
  ANDN U38059 ( .B(n33883), .A(n33884), .Z(n33881) );
  AND U38060 ( .A(a[36]), .B(b[33]), .Z(n33880) );
  XOR U38061 ( .A(n33886), .B(n33887), .Z(n33477) );
  ANDN U38062 ( .B(n33888), .A(n33889), .Z(n33886) );
  AND U38063 ( .A(a[37]), .B(b[32]), .Z(n33885) );
  XOR U38064 ( .A(n33891), .B(n33892), .Z(n33482) );
  ANDN U38065 ( .B(n33893), .A(n33894), .Z(n33891) );
  AND U38066 ( .A(a[38]), .B(b[31]), .Z(n33890) );
  XOR U38067 ( .A(n33896), .B(n33897), .Z(n33487) );
  ANDN U38068 ( .B(n33898), .A(n33899), .Z(n33896) );
  AND U38069 ( .A(a[39]), .B(b[30]), .Z(n33895) );
  XOR U38070 ( .A(n33901), .B(n33902), .Z(n33492) );
  ANDN U38071 ( .B(n33903), .A(n33904), .Z(n33901) );
  AND U38072 ( .A(a[40]), .B(b[29]), .Z(n33900) );
  XOR U38073 ( .A(n33906), .B(n33907), .Z(n33497) );
  ANDN U38074 ( .B(n33908), .A(n33909), .Z(n33906) );
  AND U38075 ( .A(a[41]), .B(b[28]), .Z(n33905) );
  XOR U38076 ( .A(n33911), .B(n33912), .Z(n33502) );
  ANDN U38077 ( .B(n33913), .A(n33914), .Z(n33911) );
  AND U38078 ( .A(a[42]), .B(b[27]), .Z(n33910) );
  XOR U38079 ( .A(n33916), .B(n33917), .Z(n33507) );
  ANDN U38080 ( .B(n33918), .A(n33919), .Z(n33916) );
  AND U38081 ( .A(a[43]), .B(b[26]), .Z(n33915) );
  XOR U38082 ( .A(n33921), .B(n33922), .Z(n33512) );
  ANDN U38083 ( .B(n33923), .A(n33924), .Z(n33921) );
  AND U38084 ( .A(a[44]), .B(b[25]), .Z(n33920) );
  XOR U38085 ( .A(n33926), .B(n33927), .Z(n33517) );
  ANDN U38086 ( .B(n33928), .A(n33929), .Z(n33926) );
  AND U38087 ( .A(a[45]), .B(b[24]), .Z(n33925) );
  XOR U38088 ( .A(n33931), .B(n33932), .Z(n33522) );
  ANDN U38089 ( .B(n33933), .A(n33934), .Z(n33931) );
  AND U38090 ( .A(a[46]), .B(b[23]), .Z(n33930) );
  XOR U38091 ( .A(n33936), .B(n33937), .Z(n33527) );
  ANDN U38092 ( .B(n33938), .A(n33939), .Z(n33936) );
  AND U38093 ( .A(a[47]), .B(b[22]), .Z(n33935) );
  XOR U38094 ( .A(n33941), .B(n33942), .Z(n33532) );
  ANDN U38095 ( .B(n33943), .A(n33944), .Z(n33941) );
  AND U38096 ( .A(a[48]), .B(b[21]), .Z(n33940) );
  XOR U38097 ( .A(n33946), .B(n33947), .Z(n33537) );
  ANDN U38098 ( .B(n33948), .A(n33949), .Z(n33946) );
  AND U38099 ( .A(a[49]), .B(b[20]), .Z(n33945) );
  XOR U38100 ( .A(n33951), .B(n33952), .Z(n33542) );
  ANDN U38101 ( .B(n33953), .A(n33954), .Z(n33951) );
  AND U38102 ( .A(a[50]), .B(b[19]), .Z(n33950) );
  XOR U38103 ( .A(n33956), .B(n33957), .Z(n33547) );
  ANDN U38104 ( .B(n33958), .A(n33959), .Z(n33956) );
  AND U38105 ( .A(a[51]), .B(b[18]), .Z(n33955) );
  XOR U38106 ( .A(n33961), .B(n33962), .Z(n33552) );
  ANDN U38107 ( .B(n33963), .A(n33964), .Z(n33961) );
  AND U38108 ( .A(a[52]), .B(b[17]), .Z(n33960) );
  XOR U38109 ( .A(n33966), .B(n33967), .Z(n33557) );
  ANDN U38110 ( .B(n33968), .A(n33969), .Z(n33966) );
  AND U38111 ( .A(a[53]), .B(b[16]), .Z(n33965) );
  XOR U38112 ( .A(n33971), .B(n33972), .Z(n33562) );
  ANDN U38113 ( .B(n33973), .A(n33974), .Z(n33971) );
  AND U38114 ( .A(a[54]), .B(b[15]), .Z(n33970) );
  XOR U38115 ( .A(n33976), .B(n33977), .Z(n33567) );
  ANDN U38116 ( .B(n33978), .A(n33979), .Z(n33976) );
  AND U38117 ( .A(a[55]), .B(b[14]), .Z(n33975) );
  XOR U38118 ( .A(n33981), .B(n33982), .Z(n33572) );
  ANDN U38119 ( .B(n33983), .A(n33984), .Z(n33981) );
  AND U38120 ( .A(a[56]), .B(b[13]), .Z(n33980) );
  XOR U38121 ( .A(n33986), .B(n33987), .Z(n33577) );
  ANDN U38122 ( .B(n33988), .A(n33989), .Z(n33986) );
  AND U38123 ( .A(a[57]), .B(b[12]), .Z(n33985) );
  XOR U38124 ( .A(n33991), .B(n33992), .Z(n33582) );
  ANDN U38125 ( .B(n33993), .A(n33994), .Z(n33991) );
  AND U38126 ( .A(a[58]), .B(b[11]), .Z(n33990) );
  XOR U38127 ( .A(n33996), .B(n33997), .Z(n33587) );
  ANDN U38128 ( .B(n33998), .A(n33999), .Z(n33996) );
  AND U38129 ( .A(a[59]), .B(b[10]), .Z(n33995) );
  XOR U38130 ( .A(n34001), .B(n34002), .Z(n33592) );
  ANDN U38131 ( .B(n34003), .A(n34004), .Z(n34001) );
  AND U38132 ( .A(b[9]), .B(a[60]), .Z(n34000) );
  XOR U38133 ( .A(n34006), .B(n34007), .Z(n33597) );
  ANDN U38134 ( .B(n34008), .A(n34009), .Z(n34006) );
  AND U38135 ( .A(b[8]), .B(a[61]), .Z(n34005) );
  XOR U38136 ( .A(n34011), .B(n34012), .Z(n33602) );
  ANDN U38137 ( .B(n34013), .A(n34014), .Z(n34011) );
  AND U38138 ( .A(b[7]), .B(a[62]), .Z(n34010) );
  XOR U38139 ( .A(n34016), .B(n34017), .Z(n33607) );
  ANDN U38140 ( .B(n34018), .A(n34019), .Z(n34016) );
  AND U38141 ( .A(b[6]), .B(a[63]), .Z(n34015) );
  XOR U38142 ( .A(n34021), .B(n34022), .Z(n33612) );
  ANDN U38143 ( .B(n34023), .A(n34024), .Z(n34021) );
  AND U38144 ( .A(b[5]), .B(a[64]), .Z(n34020) );
  XOR U38145 ( .A(n34026), .B(n34027), .Z(n33617) );
  ANDN U38146 ( .B(n34028), .A(n34029), .Z(n34026) );
  AND U38147 ( .A(b[4]), .B(a[65]), .Z(n34025) );
  XOR U38148 ( .A(n34031), .B(n34032), .Z(n33622) );
  ANDN U38149 ( .B(n33634), .A(n33635), .Z(n34031) );
  AND U38150 ( .A(b[2]), .B(a[66]), .Z(n34033) );
  XNOR U38151 ( .A(n34028), .B(n34032), .Z(n34034) );
  XOR U38152 ( .A(n34035), .B(n34036), .Z(n34032) );
  OR U38153 ( .A(n33637), .B(n33638), .Z(n34036) );
  XNOR U38154 ( .A(n34038), .B(n34039), .Z(n34037) );
  XOR U38155 ( .A(n34038), .B(n34041), .Z(n33637) );
  NAND U38156 ( .A(b[1]), .B(a[66]), .Z(n34041) );
  IV U38157 ( .A(n34035), .Z(n34038) );
  NANDN U38158 ( .A(n75), .B(n76), .Z(n34035) );
  XOR U38159 ( .A(n34042), .B(n34043), .Z(n76) );
  NAND U38160 ( .A(a[66]), .B(b[0]), .Z(n75) );
  XNOR U38161 ( .A(n34023), .B(n34027), .Z(n34044) );
  XNOR U38162 ( .A(n34018), .B(n34022), .Z(n34045) );
  XNOR U38163 ( .A(n34013), .B(n34017), .Z(n34046) );
  XNOR U38164 ( .A(n34008), .B(n34012), .Z(n34047) );
  XNOR U38165 ( .A(n34003), .B(n34007), .Z(n34048) );
  XNOR U38166 ( .A(n33998), .B(n34002), .Z(n34049) );
  XNOR U38167 ( .A(n33993), .B(n33997), .Z(n34050) );
  XNOR U38168 ( .A(n33988), .B(n33992), .Z(n34051) );
  XNOR U38169 ( .A(n33983), .B(n33987), .Z(n34052) );
  XNOR U38170 ( .A(n33978), .B(n33982), .Z(n34053) );
  XNOR U38171 ( .A(n33973), .B(n33977), .Z(n34054) );
  XNOR U38172 ( .A(n33968), .B(n33972), .Z(n34055) );
  XNOR U38173 ( .A(n33963), .B(n33967), .Z(n34056) );
  XNOR U38174 ( .A(n33958), .B(n33962), .Z(n34057) );
  XNOR U38175 ( .A(n33953), .B(n33957), .Z(n34058) );
  XNOR U38176 ( .A(n33948), .B(n33952), .Z(n34059) );
  XNOR U38177 ( .A(n33943), .B(n33947), .Z(n34060) );
  XNOR U38178 ( .A(n33938), .B(n33942), .Z(n34061) );
  XNOR U38179 ( .A(n33933), .B(n33937), .Z(n34062) );
  XNOR U38180 ( .A(n33928), .B(n33932), .Z(n34063) );
  XNOR U38181 ( .A(n33923), .B(n33927), .Z(n34064) );
  XNOR U38182 ( .A(n33918), .B(n33922), .Z(n34065) );
  XNOR U38183 ( .A(n33913), .B(n33917), .Z(n34066) );
  XNOR U38184 ( .A(n33908), .B(n33912), .Z(n34067) );
  XNOR U38185 ( .A(n33903), .B(n33907), .Z(n34068) );
  XNOR U38186 ( .A(n33898), .B(n33902), .Z(n34069) );
  XNOR U38187 ( .A(n33893), .B(n33897), .Z(n34070) );
  XNOR U38188 ( .A(n33888), .B(n33892), .Z(n34071) );
  XNOR U38189 ( .A(n33883), .B(n33887), .Z(n34072) );
  XNOR U38190 ( .A(n33878), .B(n33882), .Z(n34073) );
  XNOR U38191 ( .A(n33873), .B(n33877), .Z(n34074) );
  XNOR U38192 ( .A(n33868), .B(n33872), .Z(n34075) );
  XNOR U38193 ( .A(n33863), .B(n33867), .Z(n34076) );
  XNOR U38194 ( .A(n33858), .B(n33862), .Z(n34077) );
  XNOR U38195 ( .A(n33853), .B(n33857), .Z(n34078) );
  XNOR U38196 ( .A(n33848), .B(n33852), .Z(n34079) );
  XNOR U38197 ( .A(n33843), .B(n33847), .Z(n34080) );
  XNOR U38198 ( .A(n33838), .B(n33842), .Z(n34081) );
  XNOR U38199 ( .A(n33833), .B(n33837), .Z(n34082) );
  XNOR U38200 ( .A(n33828), .B(n33832), .Z(n34083) );
  XNOR U38201 ( .A(n33823), .B(n33827), .Z(n34084) );
  XNOR U38202 ( .A(n33818), .B(n33822), .Z(n34085) );
  XNOR U38203 ( .A(n33813), .B(n33817), .Z(n34086) );
  XNOR U38204 ( .A(n33808), .B(n33812), .Z(n34087) );
  XNOR U38205 ( .A(n33803), .B(n33807), .Z(n34088) );
  XNOR U38206 ( .A(n33798), .B(n33802), .Z(n34089) );
  XNOR U38207 ( .A(n33793), .B(n33797), .Z(n34090) );
  XNOR U38208 ( .A(n33788), .B(n33792), .Z(n34091) );
  XNOR U38209 ( .A(n33783), .B(n33787), .Z(n34092) );
  XNOR U38210 ( .A(n33778), .B(n33782), .Z(n34093) );
  XNOR U38211 ( .A(n33773), .B(n33777), .Z(n34094) );
  XNOR U38212 ( .A(n33768), .B(n33772), .Z(n34095) );
  XNOR U38213 ( .A(n33763), .B(n33767), .Z(n34096) );
  XNOR U38214 ( .A(n33758), .B(n33762), .Z(n34097) );
  XNOR U38215 ( .A(n33753), .B(n33757), .Z(n34098) );
  XNOR U38216 ( .A(n33748), .B(n33752), .Z(n34099) );
  XNOR U38217 ( .A(n33743), .B(n33747), .Z(n34100) );
  XNOR U38218 ( .A(n33738), .B(n33742), .Z(n34101) );
  XNOR U38219 ( .A(n33733), .B(n33737), .Z(n34102) );
  XNOR U38220 ( .A(n33728), .B(n33732), .Z(n34103) );
  XNOR U38221 ( .A(n33723), .B(n33727), .Z(n34104) );
  XNOR U38222 ( .A(n33718), .B(n33722), .Z(n34105) );
  XNOR U38223 ( .A(n33713), .B(n33717), .Z(n34106) );
  XNOR U38224 ( .A(n33708), .B(n33712), .Z(n34107) );
  XOR U38225 ( .A(n34108), .B(n33707), .Z(n33708) );
  AND U38226 ( .A(a[0]), .B(b[68]), .Z(n34108) );
  XNOR U38227 ( .A(n34109), .B(n33707), .Z(n33709) );
  XNOR U38228 ( .A(n34110), .B(n34111), .Z(n33707) );
  ANDN U38229 ( .B(n34112), .A(n34113), .Z(n34110) );
  AND U38230 ( .A(a[1]), .B(b[67]), .Z(n34109) );
  XOR U38231 ( .A(n34115), .B(n34116), .Z(n33712) );
  ANDN U38232 ( .B(n34117), .A(n34118), .Z(n34115) );
  AND U38233 ( .A(a[2]), .B(b[66]), .Z(n34114) );
  XOR U38234 ( .A(n34120), .B(n34121), .Z(n33717) );
  ANDN U38235 ( .B(n34122), .A(n34123), .Z(n34120) );
  AND U38236 ( .A(a[3]), .B(b[65]), .Z(n34119) );
  XOR U38237 ( .A(n34125), .B(n34126), .Z(n33722) );
  ANDN U38238 ( .B(n34127), .A(n34128), .Z(n34125) );
  AND U38239 ( .A(a[4]), .B(b[64]), .Z(n34124) );
  XOR U38240 ( .A(n34130), .B(n34131), .Z(n33727) );
  ANDN U38241 ( .B(n34132), .A(n34133), .Z(n34130) );
  AND U38242 ( .A(a[5]), .B(b[63]), .Z(n34129) );
  XOR U38243 ( .A(n34135), .B(n34136), .Z(n33732) );
  ANDN U38244 ( .B(n34137), .A(n34138), .Z(n34135) );
  AND U38245 ( .A(a[6]), .B(b[62]), .Z(n34134) );
  XOR U38246 ( .A(n34140), .B(n34141), .Z(n33737) );
  ANDN U38247 ( .B(n34142), .A(n34143), .Z(n34140) );
  AND U38248 ( .A(a[7]), .B(b[61]), .Z(n34139) );
  XOR U38249 ( .A(n34145), .B(n34146), .Z(n33742) );
  ANDN U38250 ( .B(n34147), .A(n34148), .Z(n34145) );
  AND U38251 ( .A(a[8]), .B(b[60]), .Z(n34144) );
  XOR U38252 ( .A(n34150), .B(n34151), .Z(n33747) );
  ANDN U38253 ( .B(n34152), .A(n34153), .Z(n34150) );
  AND U38254 ( .A(a[9]), .B(b[59]), .Z(n34149) );
  XOR U38255 ( .A(n34155), .B(n34156), .Z(n33752) );
  ANDN U38256 ( .B(n34157), .A(n34158), .Z(n34155) );
  AND U38257 ( .A(a[10]), .B(b[58]), .Z(n34154) );
  XOR U38258 ( .A(n34160), .B(n34161), .Z(n33757) );
  ANDN U38259 ( .B(n34162), .A(n34163), .Z(n34160) );
  AND U38260 ( .A(a[11]), .B(b[57]), .Z(n34159) );
  XOR U38261 ( .A(n34165), .B(n34166), .Z(n33762) );
  ANDN U38262 ( .B(n34167), .A(n34168), .Z(n34165) );
  AND U38263 ( .A(a[12]), .B(b[56]), .Z(n34164) );
  XOR U38264 ( .A(n34170), .B(n34171), .Z(n33767) );
  ANDN U38265 ( .B(n34172), .A(n34173), .Z(n34170) );
  AND U38266 ( .A(a[13]), .B(b[55]), .Z(n34169) );
  XOR U38267 ( .A(n34175), .B(n34176), .Z(n33772) );
  ANDN U38268 ( .B(n34177), .A(n34178), .Z(n34175) );
  AND U38269 ( .A(a[14]), .B(b[54]), .Z(n34174) );
  XOR U38270 ( .A(n34180), .B(n34181), .Z(n33777) );
  ANDN U38271 ( .B(n34182), .A(n34183), .Z(n34180) );
  AND U38272 ( .A(a[15]), .B(b[53]), .Z(n34179) );
  XOR U38273 ( .A(n34185), .B(n34186), .Z(n33782) );
  ANDN U38274 ( .B(n34187), .A(n34188), .Z(n34185) );
  AND U38275 ( .A(a[16]), .B(b[52]), .Z(n34184) );
  XOR U38276 ( .A(n34190), .B(n34191), .Z(n33787) );
  ANDN U38277 ( .B(n34192), .A(n34193), .Z(n34190) );
  AND U38278 ( .A(a[17]), .B(b[51]), .Z(n34189) );
  XOR U38279 ( .A(n34195), .B(n34196), .Z(n33792) );
  ANDN U38280 ( .B(n34197), .A(n34198), .Z(n34195) );
  AND U38281 ( .A(a[18]), .B(b[50]), .Z(n34194) );
  XOR U38282 ( .A(n34200), .B(n34201), .Z(n33797) );
  ANDN U38283 ( .B(n34202), .A(n34203), .Z(n34200) );
  AND U38284 ( .A(a[19]), .B(b[49]), .Z(n34199) );
  XOR U38285 ( .A(n34205), .B(n34206), .Z(n33802) );
  ANDN U38286 ( .B(n34207), .A(n34208), .Z(n34205) );
  AND U38287 ( .A(a[20]), .B(b[48]), .Z(n34204) );
  XOR U38288 ( .A(n34210), .B(n34211), .Z(n33807) );
  ANDN U38289 ( .B(n34212), .A(n34213), .Z(n34210) );
  AND U38290 ( .A(a[21]), .B(b[47]), .Z(n34209) );
  XOR U38291 ( .A(n34215), .B(n34216), .Z(n33812) );
  ANDN U38292 ( .B(n34217), .A(n34218), .Z(n34215) );
  AND U38293 ( .A(a[22]), .B(b[46]), .Z(n34214) );
  XOR U38294 ( .A(n34220), .B(n34221), .Z(n33817) );
  ANDN U38295 ( .B(n34222), .A(n34223), .Z(n34220) );
  AND U38296 ( .A(a[23]), .B(b[45]), .Z(n34219) );
  XOR U38297 ( .A(n34225), .B(n34226), .Z(n33822) );
  ANDN U38298 ( .B(n34227), .A(n34228), .Z(n34225) );
  AND U38299 ( .A(a[24]), .B(b[44]), .Z(n34224) );
  XOR U38300 ( .A(n34230), .B(n34231), .Z(n33827) );
  ANDN U38301 ( .B(n34232), .A(n34233), .Z(n34230) );
  AND U38302 ( .A(a[25]), .B(b[43]), .Z(n34229) );
  XOR U38303 ( .A(n34235), .B(n34236), .Z(n33832) );
  ANDN U38304 ( .B(n34237), .A(n34238), .Z(n34235) );
  AND U38305 ( .A(a[26]), .B(b[42]), .Z(n34234) );
  XOR U38306 ( .A(n34240), .B(n34241), .Z(n33837) );
  ANDN U38307 ( .B(n34242), .A(n34243), .Z(n34240) );
  AND U38308 ( .A(a[27]), .B(b[41]), .Z(n34239) );
  XOR U38309 ( .A(n34245), .B(n34246), .Z(n33842) );
  ANDN U38310 ( .B(n34247), .A(n34248), .Z(n34245) );
  AND U38311 ( .A(a[28]), .B(b[40]), .Z(n34244) );
  XOR U38312 ( .A(n34250), .B(n34251), .Z(n33847) );
  ANDN U38313 ( .B(n34252), .A(n34253), .Z(n34250) );
  AND U38314 ( .A(a[29]), .B(b[39]), .Z(n34249) );
  XOR U38315 ( .A(n34255), .B(n34256), .Z(n33852) );
  ANDN U38316 ( .B(n34257), .A(n34258), .Z(n34255) );
  AND U38317 ( .A(a[30]), .B(b[38]), .Z(n34254) );
  XOR U38318 ( .A(n34260), .B(n34261), .Z(n33857) );
  ANDN U38319 ( .B(n34262), .A(n34263), .Z(n34260) );
  AND U38320 ( .A(a[31]), .B(b[37]), .Z(n34259) );
  XOR U38321 ( .A(n34265), .B(n34266), .Z(n33862) );
  ANDN U38322 ( .B(n34267), .A(n34268), .Z(n34265) );
  AND U38323 ( .A(a[32]), .B(b[36]), .Z(n34264) );
  XOR U38324 ( .A(n34270), .B(n34271), .Z(n33867) );
  ANDN U38325 ( .B(n34272), .A(n34273), .Z(n34270) );
  AND U38326 ( .A(a[33]), .B(b[35]), .Z(n34269) );
  XOR U38327 ( .A(n34275), .B(n34276), .Z(n33872) );
  ANDN U38328 ( .B(n34277), .A(n34278), .Z(n34275) );
  AND U38329 ( .A(a[34]), .B(b[34]), .Z(n34274) );
  XOR U38330 ( .A(n34280), .B(n34281), .Z(n33877) );
  ANDN U38331 ( .B(n34282), .A(n34283), .Z(n34280) );
  AND U38332 ( .A(a[35]), .B(b[33]), .Z(n34279) );
  XOR U38333 ( .A(n34285), .B(n34286), .Z(n33882) );
  ANDN U38334 ( .B(n34287), .A(n34288), .Z(n34285) );
  AND U38335 ( .A(a[36]), .B(b[32]), .Z(n34284) );
  XOR U38336 ( .A(n34290), .B(n34291), .Z(n33887) );
  ANDN U38337 ( .B(n34292), .A(n34293), .Z(n34290) );
  AND U38338 ( .A(a[37]), .B(b[31]), .Z(n34289) );
  XOR U38339 ( .A(n34295), .B(n34296), .Z(n33892) );
  ANDN U38340 ( .B(n34297), .A(n34298), .Z(n34295) );
  AND U38341 ( .A(a[38]), .B(b[30]), .Z(n34294) );
  XOR U38342 ( .A(n34300), .B(n34301), .Z(n33897) );
  ANDN U38343 ( .B(n34302), .A(n34303), .Z(n34300) );
  AND U38344 ( .A(a[39]), .B(b[29]), .Z(n34299) );
  XOR U38345 ( .A(n34305), .B(n34306), .Z(n33902) );
  ANDN U38346 ( .B(n34307), .A(n34308), .Z(n34305) );
  AND U38347 ( .A(a[40]), .B(b[28]), .Z(n34304) );
  XOR U38348 ( .A(n34310), .B(n34311), .Z(n33907) );
  ANDN U38349 ( .B(n34312), .A(n34313), .Z(n34310) );
  AND U38350 ( .A(a[41]), .B(b[27]), .Z(n34309) );
  XOR U38351 ( .A(n34315), .B(n34316), .Z(n33912) );
  ANDN U38352 ( .B(n34317), .A(n34318), .Z(n34315) );
  AND U38353 ( .A(a[42]), .B(b[26]), .Z(n34314) );
  XOR U38354 ( .A(n34320), .B(n34321), .Z(n33917) );
  ANDN U38355 ( .B(n34322), .A(n34323), .Z(n34320) );
  AND U38356 ( .A(a[43]), .B(b[25]), .Z(n34319) );
  XOR U38357 ( .A(n34325), .B(n34326), .Z(n33922) );
  ANDN U38358 ( .B(n34327), .A(n34328), .Z(n34325) );
  AND U38359 ( .A(a[44]), .B(b[24]), .Z(n34324) );
  XOR U38360 ( .A(n34330), .B(n34331), .Z(n33927) );
  ANDN U38361 ( .B(n34332), .A(n34333), .Z(n34330) );
  AND U38362 ( .A(a[45]), .B(b[23]), .Z(n34329) );
  XOR U38363 ( .A(n34335), .B(n34336), .Z(n33932) );
  ANDN U38364 ( .B(n34337), .A(n34338), .Z(n34335) );
  AND U38365 ( .A(a[46]), .B(b[22]), .Z(n34334) );
  XOR U38366 ( .A(n34340), .B(n34341), .Z(n33937) );
  ANDN U38367 ( .B(n34342), .A(n34343), .Z(n34340) );
  AND U38368 ( .A(a[47]), .B(b[21]), .Z(n34339) );
  XOR U38369 ( .A(n34345), .B(n34346), .Z(n33942) );
  ANDN U38370 ( .B(n34347), .A(n34348), .Z(n34345) );
  AND U38371 ( .A(a[48]), .B(b[20]), .Z(n34344) );
  XOR U38372 ( .A(n34350), .B(n34351), .Z(n33947) );
  ANDN U38373 ( .B(n34352), .A(n34353), .Z(n34350) );
  AND U38374 ( .A(a[49]), .B(b[19]), .Z(n34349) );
  XOR U38375 ( .A(n34355), .B(n34356), .Z(n33952) );
  ANDN U38376 ( .B(n34357), .A(n34358), .Z(n34355) );
  AND U38377 ( .A(a[50]), .B(b[18]), .Z(n34354) );
  XOR U38378 ( .A(n34360), .B(n34361), .Z(n33957) );
  ANDN U38379 ( .B(n34362), .A(n34363), .Z(n34360) );
  AND U38380 ( .A(a[51]), .B(b[17]), .Z(n34359) );
  XOR U38381 ( .A(n34365), .B(n34366), .Z(n33962) );
  ANDN U38382 ( .B(n34367), .A(n34368), .Z(n34365) );
  AND U38383 ( .A(a[52]), .B(b[16]), .Z(n34364) );
  XOR U38384 ( .A(n34370), .B(n34371), .Z(n33967) );
  ANDN U38385 ( .B(n34372), .A(n34373), .Z(n34370) );
  AND U38386 ( .A(a[53]), .B(b[15]), .Z(n34369) );
  XOR U38387 ( .A(n34375), .B(n34376), .Z(n33972) );
  ANDN U38388 ( .B(n34377), .A(n34378), .Z(n34375) );
  AND U38389 ( .A(a[54]), .B(b[14]), .Z(n34374) );
  XOR U38390 ( .A(n34380), .B(n34381), .Z(n33977) );
  ANDN U38391 ( .B(n34382), .A(n34383), .Z(n34380) );
  AND U38392 ( .A(a[55]), .B(b[13]), .Z(n34379) );
  XOR U38393 ( .A(n34385), .B(n34386), .Z(n33982) );
  ANDN U38394 ( .B(n34387), .A(n34388), .Z(n34385) );
  AND U38395 ( .A(a[56]), .B(b[12]), .Z(n34384) );
  XOR U38396 ( .A(n34390), .B(n34391), .Z(n33987) );
  ANDN U38397 ( .B(n34392), .A(n34393), .Z(n34390) );
  AND U38398 ( .A(a[57]), .B(b[11]), .Z(n34389) );
  XOR U38399 ( .A(n34395), .B(n34396), .Z(n33992) );
  ANDN U38400 ( .B(n34397), .A(n34398), .Z(n34395) );
  AND U38401 ( .A(a[58]), .B(b[10]), .Z(n34394) );
  XOR U38402 ( .A(n34400), .B(n34401), .Z(n33997) );
  ANDN U38403 ( .B(n34402), .A(n34403), .Z(n34400) );
  AND U38404 ( .A(b[9]), .B(a[59]), .Z(n34399) );
  XOR U38405 ( .A(n34405), .B(n34406), .Z(n34002) );
  ANDN U38406 ( .B(n34407), .A(n34408), .Z(n34405) );
  AND U38407 ( .A(b[8]), .B(a[60]), .Z(n34404) );
  XOR U38408 ( .A(n34410), .B(n34411), .Z(n34007) );
  ANDN U38409 ( .B(n34412), .A(n34413), .Z(n34410) );
  AND U38410 ( .A(b[7]), .B(a[61]), .Z(n34409) );
  XOR U38411 ( .A(n34415), .B(n34416), .Z(n34012) );
  ANDN U38412 ( .B(n34417), .A(n34418), .Z(n34415) );
  AND U38413 ( .A(b[6]), .B(a[62]), .Z(n34414) );
  XOR U38414 ( .A(n34420), .B(n34421), .Z(n34017) );
  ANDN U38415 ( .B(n34422), .A(n34423), .Z(n34420) );
  AND U38416 ( .A(b[5]), .B(a[63]), .Z(n34419) );
  XOR U38417 ( .A(n34425), .B(n34426), .Z(n34022) );
  ANDN U38418 ( .B(n34427), .A(n34428), .Z(n34425) );
  AND U38419 ( .A(b[4]), .B(a[64]), .Z(n34424) );
  XOR U38420 ( .A(n34430), .B(n34431), .Z(n34027) );
  ANDN U38421 ( .B(n34039), .A(n34040), .Z(n34430) );
  AND U38422 ( .A(b[2]), .B(a[65]), .Z(n34432) );
  XNOR U38423 ( .A(n34427), .B(n34431), .Z(n34433) );
  XOR U38424 ( .A(n34434), .B(n34435), .Z(n34431) );
  OR U38425 ( .A(n34042), .B(n34043), .Z(n34435) );
  XNOR U38426 ( .A(n34437), .B(n34438), .Z(n34436) );
  XOR U38427 ( .A(n34437), .B(n34440), .Z(n34042) );
  NAND U38428 ( .A(b[1]), .B(a[65]), .Z(n34440) );
  IV U38429 ( .A(n34434), .Z(n34437) );
  NANDN U38430 ( .A(n77), .B(n78), .Z(n34434) );
  XOR U38431 ( .A(n34441), .B(n34442), .Z(n78) );
  NAND U38432 ( .A(a[65]), .B(b[0]), .Z(n77) );
  XNOR U38433 ( .A(n34422), .B(n34426), .Z(n34443) );
  XNOR U38434 ( .A(n34417), .B(n34421), .Z(n34444) );
  XNOR U38435 ( .A(n34412), .B(n34416), .Z(n34445) );
  XNOR U38436 ( .A(n34407), .B(n34411), .Z(n34446) );
  XNOR U38437 ( .A(n34402), .B(n34406), .Z(n34447) );
  XNOR U38438 ( .A(n34397), .B(n34401), .Z(n34448) );
  XNOR U38439 ( .A(n34392), .B(n34396), .Z(n34449) );
  XNOR U38440 ( .A(n34387), .B(n34391), .Z(n34450) );
  XNOR U38441 ( .A(n34382), .B(n34386), .Z(n34451) );
  XNOR U38442 ( .A(n34377), .B(n34381), .Z(n34452) );
  XNOR U38443 ( .A(n34372), .B(n34376), .Z(n34453) );
  XNOR U38444 ( .A(n34367), .B(n34371), .Z(n34454) );
  XNOR U38445 ( .A(n34362), .B(n34366), .Z(n34455) );
  XNOR U38446 ( .A(n34357), .B(n34361), .Z(n34456) );
  XNOR U38447 ( .A(n34352), .B(n34356), .Z(n34457) );
  XNOR U38448 ( .A(n34347), .B(n34351), .Z(n34458) );
  XNOR U38449 ( .A(n34342), .B(n34346), .Z(n34459) );
  XNOR U38450 ( .A(n34337), .B(n34341), .Z(n34460) );
  XNOR U38451 ( .A(n34332), .B(n34336), .Z(n34461) );
  XNOR U38452 ( .A(n34327), .B(n34331), .Z(n34462) );
  XNOR U38453 ( .A(n34322), .B(n34326), .Z(n34463) );
  XNOR U38454 ( .A(n34317), .B(n34321), .Z(n34464) );
  XNOR U38455 ( .A(n34312), .B(n34316), .Z(n34465) );
  XNOR U38456 ( .A(n34307), .B(n34311), .Z(n34466) );
  XNOR U38457 ( .A(n34302), .B(n34306), .Z(n34467) );
  XNOR U38458 ( .A(n34297), .B(n34301), .Z(n34468) );
  XNOR U38459 ( .A(n34292), .B(n34296), .Z(n34469) );
  XNOR U38460 ( .A(n34287), .B(n34291), .Z(n34470) );
  XNOR U38461 ( .A(n34282), .B(n34286), .Z(n34471) );
  XNOR U38462 ( .A(n34277), .B(n34281), .Z(n34472) );
  XNOR U38463 ( .A(n34272), .B(n34276), .Z(n34473) );
  XNOR U38464 ( .A(n34267), .B(n34271), .Z(n34474) );
  XNOR U38465 ( .A(n34262), .B(n34266), .Z(n34475) );
  XNOR U38466 ( .A(n34257), .B(n34261), .Z(n34476) );
  XNOR U38467 ( .A(n34252), .B(n34256), .Z(n34477) );
  XNOR U38468 ( .A(n34247), .B(n34251), .Z(n34478) );
  XNOR U38469 ( .A(n34242), .B(n34246), .Z(n34479) );
  XNOR U38470 ( .A(n34237), .B(n34241), .Z(n34480) );
  XNOR U38471 ( .A(n34232), .B(n34236), .Z(n34481) );
  XNOR U38472 ( .A(n34227), .B(n34231), .Z(n34482) );
  XNOR U38473 ( .A(n34222), .B(n34226), .Z(n34483) );
  XNOR U38474 ( .A(n34217), .B(n34221), .Z(n34484) );
  XNOR U38475 ( .A(n34212), .B(n34216), .Z(n34485) );
  XNOR U38476 ( .A(n34207), .B(n34211), .Z(n34486) );
  XNOR U38477 ( .A(n34202), .B(n34206), .Z(n34487) );
  XNOR U38478 ( .A(n34197), .B(n34201), .Z(n34488) );
  XNOR U38479 ( .A(n34192), .B(n34196), .Z(n34489) );
  XNOR U38480 ( .A(n34187), .B(n34191), .Z(n34490) );
  XNOR U38481 ( .A(n34182), .B(n34186), .Z(n34491) );
  XNOR U38482 ( .A(n34177), .B(n34181), .Z(n34492) );
  XNOR U38483 ( .A(n34172), .B(n34176), .Z(n34493) );
  XNOR U38484 ( .A(n34167), .B(n34171), .Z(n34494) );
  XNOR U38485 ( .A(n34162), .B(n34166), .Z(n34495) );
  XNOR U38486 ( .A(n34157), .B(n34161), .Z(n34496) );
  XNOR U38487 ( .A(n34152), .B(n34156), .Z(n34497) );
  XNOR U38488 ( .A(n34147), .B(n34151), .Z(n34498) );
  XNOR U38489 ( .A(n34142), .B(n34146), .Z(n34499) );
  XNOR U38490 ( .A(n34137), .B(n34141), .Z(n34500) );
  XNOR U38491 ( .A(n34132), .B(n34136), .Z(n34501) );
  XNOR U38492 ( .A(n34127), .B(n34131), .Z(n34502) );
  XNOR U38493 ( .A(n34122), .B(n34126), .Z(n34503) );
  XNOR U38494 ( .A(n34117), .B(n34121), .Z(n34504) );
  XNOR U38495 ( .A(n34112), .B(n34116), .Z(n34505) );
  XNOR U38496 ( .A(n34506), .B(n34111), .Z(n34112) );
  AND U38497 ( .A(a[0]), .B(b[67]), .Z(n34506) );
  XOR U38498 ( .A(n34507), .B(n34111), .Z(n34113) );
  XNOR U38499 ( .A(n34508), .B(n34509), .Z(n34111) );
  ANDN U38500 ( .B(n34510), .A(n34511), .Z(n34508) );
  AND U38501 ( .A(a[1]), .B(b[66]), .Z(n34507) );
  XOR U38502 ( .A(n34513), .B(n34514), .Z(n34116) );
  ANDN U38503 ( .B(n34515), .A(n34516), .Z(n34513) );
  AND U38504 ( .A(a[2]), .B(b[65]), .Z(n34512) );
  XOR U38505 ( .A(n34518), .B(n34519), .Z(n34121) );
  ANDN U38506 ( .B(n34520), .A(n34521), .Z(n34518) );
  AND U38507 ( .A(a[3]), .B(b[64]), .Z(n34517) );
  XOR U38508 ( .A(n34523), .B(n34524), .Z(n34126) );
  ANDN U38509 ( .B(n34525), .A(n34526), .Z(n34523) );
  AND U38510 ( .A(a[4]), .B(b[63]), .Z(n34522) );
  XOR U38511 ( .A(n34528), .B(n34529), .Z(n34131) );
  ANDN U38512 ( .B(n34530), .A(n34531), .Z(n34528) );
  AND U38513 ( .A(a[5]), .B(b[62]), .Z(n34527) );
  XOR U38514 ( .A(n34533), .B(n34534), .Z(n34136) );
  ANDN U38515 ( .B(n34535), .A(n34536), .Z(n34533) );
  AND U38516 ( .A(a[6]), .B(b[61]), .Z(n34532) );
  XOR U38517 ( .A(n34538), .B(n34539), .Z(n34141) );
  ANDN U38518 ( .B(n34540), .A(n34541), .Z(n34538) );
  AND U38519 ( .A(a[7]), .B(b[60]), .Z(n34537) );
  XOR U38520 ( .A(n34543), .B(n34544), .Z(n34146) );
  ANDN U38521 ( .B(n34545), .A(n34546), .Z(n34543) );
  AND U38522 ( .A(a[8]), .B(b[59]), .Z(n34542) );
  XOR U38523 ( .A(n34548), .B(n34549), .Z(n34151) );
  ANDN U38524 ( .B(n34550), .A(n34551), .Z(n34548) );
  AND U38525 ( .A(a[9]), .B(b[58]), .Z(n34547) );
  XOR U38526 ( .A(n34553), .B(n34554), .Z(n34156) );
  ANDN U38527 ( .B(n34555), .A(n34556), .Z(n34553) );
  AND U38528 ( .A(a[10]), .B(b[57]), .Z(n34552) );
  XOR U38529 ( .A(n34558), .B(n34559), .Z(n34161) );
  ANDN U38530 ( .B(n34560), .A(n34561), .Z(n34558) );
  AND U38531 ( .A(a[11]), .B(b[56]), .Z(n34557) );
  XOR U38532 ( .A(n34563), .B(n34564), .Z(n34166) );
  ANDN U38533 ( .B(n34565), .A(n34566), .Z(n34563) );
  AND U38534 ( .A(a[12]), .B(b[55]), .Z(n34562) );
  XOR U38535 ( .A(n34568), .B(n34569), .Z(n34171) );
  ANDN U38536 ( .B(n34570), .A(n34571), .Z(n34568) );
  AND U38537 ( .A(a[13]), .B(b[54]), .Z(n34567) );
  XOR U38538 ( .A(n34573), .B(n34574), .Z(n34176) );
  ANDN U38539 ( .B(n34575), .A(n34576), .Z(n34573) );
  AND U38540 ( .A(a[14]), .B(b[53]), .Z(n34572) );
  XOR U38541 ( .A(n34578), .B(n34579), .Z(n34181) );
  ANDN U38542 ( .B(n34580), .A(n34581), .Z(n34578) );
  AND U38543 ( .A(a[15]), .B(b[52]), .Z(n34577) );
  XOR U38544 ( .A(n34583), .B(n34584), .Z(n34186) );
  ANDN U38545 ( .B(n34585), .A(n34586), .Z(n34583) );
  AND U38546 ( .A(a[16]), .B(b[51]), .Z(n34582) );
  XOR U38547 ( .A(n34588), .B(n34589), .Z(n34191) );
  ANDN U38548 ( .B(n34590), .A(n34591), .Z(n34588) );
  AND U38549 ( .A(a[17]), .B(b[50]), .Z(n34587) );
  XOR U38550 ( .A(n34593), .B(n34594), .Z(n34196) );
  ANDN U38551 ( .B(n34595), .A(n34596), .Z(n34593) );
  AND U38552 ( .A(a[18]), .B(b[49]), .Z(n34592) );
  XOR U38553 ( .A(n34598), .B(n34599), .Z(n34201) );
  ANDN U38554 ( .B(n34600), .A(n34601), .Z(n34598) );
  AND U38555 ( .A(a[19]), .B(b[48]), .Z(n34597) );
  XOR U38556 ( .A(n34603), .B(n34604), .Z(n34206) );
  ANDN U38557 ( .B(n34605), .A(n34606), .Z(n34603) );
  AND U38558 ( .A(a[20]), .B(b[47]), .Z(n34602) );
  XOR U38559 ( .A(n34608), .B(n34609), .Z(n34211) );
  ANDN U38560 ( .B(n34610), .A(n34611), .Z(n34608) );
  AND U38561 ( .A(a[21]), .B(b[46]), .Z(n34607) );
  XOR U38562 ( .A(n34613), .B(n34614), .Z(n34216) );
  ANDN U38563 ( .B(n34615), .A(n34616), .Z(n34613) );
  AND U38564 ( .A(a[22]), .B(b[45]), .Z(n34612) );
  XOR U38565 ( .A(n34618), .B(n34619), .Z(n34221) );
  ANDN U38566 ( .B(n34620), .A(n34621), .Z(n34618) );
  AND U38567 ( .A(a[23]), .B(b[44]), .Z(n34617) );
  XOR U38568 ( .A(n34623), .B(n34624), .Z(n34226) );
  ANDN U38569 ( .B(n34625), .A(n34626), .Z(n34623) );
  AND U38570 ( .A(a[24]), .B(b[43]), .Z(n34622) );
  XOR U38571 ( .A(n34628), .B(n34629), .Z(n34231) );
  ANDN U38572 ( .B(n34630), .A(n34631), .Z(n34628) );
  AND U38573 ( .A(a[25]), .B(b[42]), .Z(n34627) );
  XOR U38574 ( .A(n34633), .B(n34634), .Z(n34236) );
  ANDN U38575 ( .B(n34635), .A(n34636), .Z(n34633) );
  AND U38576 ( .A(a[26]), .B(b[41]), .Z(n34632) );
  XOR U38577 ( .A(n34638), .B(n34639), .Z(n34241) );
  ANDN U38578 ( .B(n34640), .A(n34641), .Z(n34638) );
  AND U38579 ( .A(a[27]), .B(b[40]), .Z(n34637) );
  XOR U38580 ( .A(n34643), .B(n34644), .Z(n34246) );
  ANDN U38581 ( .B(n34645), .A(n34646), .Z(n34643) );
  AND U38582 ( .A(a[28]), .B(b[39]), .Z(n34642) );
  XOR U38583 ( .A(n34648), .B(n34649), .Z(n34251) );
  ANDN U38584 ( .B(n34650), .A(n34651), .Z(n34648) );
  AND U38585 ( .A(a[29]), .B(b[38]), .Z(n34647) );
  XOR U38586 ( .A(n34653), .B(n34654), .Z(n34256) );
  ANDN U38587 ( .B(n34655), .A(n34656), .Z(n34653) );
  AND U38588 ( .A(a[30]), .B(b[37]), .Z(n34652) );
  XOR U38589 ( .A(n34658), .B(n34659), .Z(n34261) );
  ANDN U38590 ( .B(n34660), .A(n34661), .Z(n34658) );
  AND U38591 ( .A(a[31]), .B(b[36]), .Z(n34657) );
  XOR U38592 ( .A(n34663), .B(n34664), .Z(n34266) );
  ANDN U38593 ( .B(n34665), .A(n34666), .Z(n34663) );
  AND U38594 ( .A(a[32]), .B(b[35]), .Z(n34662) );
  XOR U38595 ( .A(n34668), .B(n34669), .Z(n34271) );
  ANDN U38596 ( .B(n34670), .A(n34671), .Z(n34668) );
  AND U38597 ( .A(a[33]), .B(b[34]), .Z(n34667) );
  XOR U38598 ( .A(n34673), .B(n34674), .Z(n34276) );
  ANDN U38599 ( .B(n34675), .A(n34676), .Z(n34673) );
  AND U38600 ( .A(a[34]), .B(b[33]), .Z(n34672) );
  XOR U38601 ( .A(n34678), .B(n34679), .Z(n34281) );
  ANDN U38602 ( .B(n34680), .A(n34681), .Z(n34678) );
  AND U38603 ( .A(a[35]), .B(b[32]), .Z(n34677) );
  XOR U38604 ( .A(n34683), .B(n34684), .Z(n34286) );
  ANDN U38605 ( .B(n34685), .A(n34686), .Z(n34683) );
  AND U38606 ( .A(a[36]), .B(b[31]), .Z(n34682) );
  XOR U38607 ( .A(n34688), .B(n34689), .Z(n34291) );
  ANDN U38608 ( .B(n34690), .A(n34691), .Z(n34688) );
  AND U38609 ( .A(a[37]), .B(b[30]), .Z(n34687) );
  XOR U38610 ( .A(n34693), .B(n34694), .Z(n34296) );
  ANDN U38611 ( .B(n34695), .A(n34696), .Z(n34693) );
  AND U38612 ( .A(a[38]), .B(b[29]), .Z(n34692) );
  XOR U38613 ( .A(n34698), .B(n34699), .Z(n34301) );
  ANDN U38614 ( .B(n34700), .A(n34701), .Z(n34698) );
  AND U38615 ( .A(a[39]), .B(b[28]), .Z(n34697) );
  XOR U38616 ( .A(n34703), .B(n34704), .Z(n34306) );
  ANDN U38617 ( .B(n34705), .A(n34706), .Z(n34703) );
  AND U38618 ( .A(a[40]), .B(b[27]), .Z(n34702) );
  XOR U38619 ( .A(n34708), .B(n34709), .Z(n34311) );
  ANDN U38620 ( .B(n34710), .A(n34711), .Z(n34708) );
  AND U38621 ( .A(a[41]), .B(b[26]), .Z(n34707) );
  XOR U38622 ( .A(n34713), .B(n34714), .Z(n34316) );
  ANDN U38623 ( .B(n34715), .A(n34716), .Z(n34713) );
  AND U38624 ( .A(a[42]), .B(b[25]), .Z(n34712) );
  XOR U38625 ( .A(n34718), .B(n34719), .Z(n34321) );
  ANDN U38626 ( .B(n34720), .A(n34721), .Z(n34718) );
  AND U38627 ( .A(a[43]), .B(b[24]), .Z(n34717) );
  XOR U38628 ( .A(n34723), .B(n34724), .Z(n34326) );
  ANDN U38629 ( .B(n34725), .A(n34726), .Z(n34723) );
  AND U38630 ( .A(a[44]), .B(b[23]), .Z(n34722) );
  XOR U38631 ( .A(n34728), .B(n34729), .Z(n34331) );
  ANDN U38632 ( .B(n34730), .A(n34731), .Z(n34728) );
  AND U38633 ( .A(a[45]), .B(b[22]), .Z(n34727) );
  XOR U38634 ( .A(n34733), .B(n34734), .Z(n34336) );
  ANDN U38635 ( .B(n34735), .A(n34736), .Z(n34733) );
  AND U38636 ( .A(a[46]), .B(b[21]), .Z(n34732) );
  XOR U38637 ( .A(n34738), .B(n34739), .Z(n34341) );
  ANDN U38638 ( .B(n34740), .A(n34741), .Z(n34738) );
  AND U38639 ( .A(a[47]), .B(b[20]), .Z(n34737) );
  XOR U38640 ( .A(n34743), .B(n34744), .Z(n34346) );
  ANDN U38641 ( .B(n34745), .A(n34746), .Z(n34743) );
  AND U38642 ( .A(a[48]), .B(b[19]), .Z(n34742) );
  XOR U38643 ( .A(n34748), .B(n34749), .Z(n34351) );
  ANDN U38644 ( .B(n34750), .A(n34751), .Z(n34748) );
  AND U38645 ( .A(a[49]), .B(b[18]), .Z(n34747) );
  XOR U38646 ( .A(n34753), .B(n34754), .Z(n34356) );
  ANDN U38647 ( .B(n34755), .A(n34756), .Z(n34753) );
  AND U38648 ( .A(a[50]), .B(b[17]), .Z(n34752) );
  XOR U38649 ( .A(n34758), .B(n34759), .Z(n34361) );
  ANDN U38650 ( .B(n34760), .A(n34761), .Z(n34758) );
  AND U38651 ( .A(a[51]), .B(b[16]), .Z(n34757) );
  XOR U38652 ( .A(n34763), .B(n34764), .Z(n34366) );
  ANDN U38653 ( .B(n34765), .A(n34766), .Z(n34763) );
  AND U38654 ( .A(a[52]), .B(b[15]), .Z(n34762) );
  XOR U38655 ( .A(n34768), .B(n34769), .Z(n34371) );
  ANDN U38656 ( .B(n34770), .A(n34771), .Z(n34768) );
  AND U38657 ( .A(a[53]), .B(b[14]), .Z(n34767) );
  XOR U38658 ( .A(n34773), .B(n34774), .Z(n34376) );
  ANDN U38659 ( .B(n34775), .A(n34776), .Z(n34773) );
  AND U38660 ( .A(a[54]), .B(b[13]), .Z(n34772) );
  XOR U38661 ( .A(n34778), .B(n34779), .Z(n34381) );
  ANDN U38662 ( .B(n34780), .A(n34781), .Z(n34778) );
  AND U38663 ( .A(a[55]), .B(b[12]), .Z(n34777) );
  XOR U38664 ( .A(n34783), .B(n34784), .Z(n34386) );
  ANDN U38665 ( .B(n34785), .A(n34786), .Z(n34783) );
  AND U38666 ( .A(a[56]), .B(b[11]), .Z(n34782) );
  XOR U38667 ( .A(n34788), .B(n34789), .Z(n34391) );
  ANDN U38668 ( .B(n34790), .A(n34791), .Z(n34788) );
  AND U38669 ( .A(a[57]), .B(b[10]), .Z(n34787) );
  XOR U38670 ( .A(n34793), .B(n34794), .Z(n34396) );
  ANDN U38671 ( .B(n34795), .A(n34796), .Z(n34793) );
  AND U38672 ( .A(b[9]), .B(a[58]), .Z(n34792) );
  XOR U38673 ( .A(n34798), .B(n34799), .Z(n34401) );
  ANDN U38674 ( .B(n34800), .A(n34801), .Z(n34798) );
  AND U38675 ( .A(b[8]), .B(a[59]), .Z(n34797) );
  XOR U38676 ( .A(n34803), .B(n34804), .Z(n34406) );
  ANDN U38677 ( .B(n34805), .A(n34806), .Z(n34803) );
  AND U38678 ( .A(b[7]), .B(a[60]), .Z(n34802) );
  XOR U38679 ( .A(n34808), .B(n34809), .Z(n34411) );
  ANDN U38680 ( .B(n34810), .A(n34811), .Z(n34808) );
  AND U38681 ( .A(b[6]), .B(a[61]), .Z(n34807) );
  XOR U38682 ( .A(n34813), .B(n34814), .Z(n34416) );
  ANDN U38683 ( .B(n34815), .A(n34816), .Z(n34813) );
  AND U38684 ( .A(b[5]), .B(a[62]), .Z(n34812) );
  XOR U38685 ( .A(n34818), .B(n34819), .Z(n34421) );
  ANDN U38686 ( .B(n34820), .A(n34821), .Z(n34818) );
  AND U38687 ( .A(b[4]), .B(a[63]), .Z(n34817) );
  XOR U38688 ( .A(n34823), .B(n34824), .Z(n34426) );
  ANDN U38689 ( .B(n34438), .A(n34439), .Z(n34823) );
  AND U38690 ( .A(b[2]), .B(a[64]), .Z(n34825) );
  XNOR U38691 ( .A(n34820), .B(n34824), .Z(n34826) );
  XOR U38692 ( .A(n34827), .B(n34828), .Z(n34824) );
  OR U38693 ( .A(n34441), .B(n34442), .Z(n34828) );
  XNOR U38694 ( .A(n34830), .B(n34831), .Z(n34829) );
  XOR U38695 ( .A(n34830), .B(n34833), .Z(n34441) );
  NAND U38696 ( .A(b[1]), .B(a[64]), .Z(n34833) );
  IV U38697 ( .A(n34827), .Z(n34830) );
  NANDN U38698 ( .A(n79), .B(n80), .Z(n34827) );
  XOR U38699 ( .A(n34834), .B(n34835), .Z(n80) );
  NAND U38700 ( .A(a[64]), .B(b[0]), .Z(n79) );
  XNOR U38701 ( .A(n34815), .B(n34819), .Z(n34836) );
  XNOR U38702 ( .A(n34810), .B(n34814), .Z(n34837) );
  XNOR U38703 ( .A(n34805), .B(n34809), .Z(n34838) );
  XNOR U38704 ( .A(n34800), .B(n34804), .Z(n34839) );
  XNOR U38705 ( .A(n34795), .B(n34799), .Z(n34840) );
  XNOR U38706 ( .A(n34790), .B(n34794), .Z(n34841) );
  XNOR U38707 ( .A(n34785), .B(n34789), .Z(n34842) );
  XNOR U38708 ( .A(n34780), .B(n34784), .Z(n34843) );
  XNOR U38709 ( .A(n34775), .B(n34779), .Z(n34844) );
  XNOR U38710 ( .A(n34770), .B(n34774), .Z(n34845) );
  XNOR U38711 ( .A(n34765), .B(n34769), .Z(n34846) );
  XNOR U38712 ( .A(n34760), .B(n34764), .Z(n34847) );
  XNOR U38713 ( .A(n34755), .B(n34759), .Z(n34848) );
  XNOR U38714 ( .A(n34750), .B(n34754), .Z(n34849) );
  XNOR U38715 ( .A(n34745), .B(n34749), .Z(n34850) );
  XNOR U38716 ( .A(n34740), .B(n34744), .Z(n34851) );
  XNOR U38717 ( .A(n34735), .B(n34739), .Z(n34852) );
  XNOR U38718 ( .A(n34730), .B(n34734), .Z(n34853) );
  XNOR U38719 ( .A(n34725), .B(n34729), .Z(n34854) );
  XNOR U38720 ( .A(n34720), .B(n34724), .Z(n34855) );
  XNOR U38721 ( .A(n34715), .B(n34719), .Z(n34856) );
  XNOR U38722 ( .A(n34710), .B(n34714), .Z(n34857) );
  XNOR U38723 ( .A(n34705), .B(n34709), .Z(n34858) );
  XNOR U38724 ( .A(n34700), .B(n34704), .Z(n34859) );
  XNOR U38725 ( .A(n34695), .B(n34699), .Z(n34860) );
  XNOR U38726 ( .A(n34690), .B(n34694), .Z(n34861) );
  XNOR U38727 ( .A(n34685), .B(n34689), .Z(n34862) );
  XNOR U38728 ( .A(n34680), .B(n34684), .Z(n34863) );
  XNOR U38729 ( .A(n34675), .B(n34679), .Z(n34864) );
  XNOR U38730 ( .A(n34670), .B(n34674), .Z(n34865) );
  XNOR U38731 ( .A(n34665), .B(n34669), .Z(n34866) );
  XNOR U38732 ( .A(n34660), .B(n34664), .Z(n34867) );
  XNOR U38733 ( .A(n34655), .B(n34659), .Z(n34868) );
  XNOR U38734 ( .A(n34650), .B(n34654), .Z(n34869) );
  XNOR U38735 ( .A(n34645), .B(n34649), .Z(n34870) );
  XNOR U38736 ( .A(n34640), .B(n34644), .Z(n34871) );
  XNOR U38737 ( .A(n34635), .B(n34639), .Z(n34872) );
  XNOR U38738 ( .A(n34630), .B(n34634), .Z(n34873) );
  XNOR U38739 ( .A(n34625), .B(n34629), .Z(n34874) );
  XNOR U38740 ( .A(n34620), .B(n34624), .Z(n34875) );
  XNOR U38741 ( .A(n34615), .B(n34619), .Z(n34876) );
  XNOR U38742 ( .A(n34610), .B(n34614), .Z(n34877) );
  XNOR U38743 ( .A(n34605), .B(n34609), .Z(n34878) );
  XNOR U38744 ( .A(n34600), .B(n34604), .Z(n34879) );
  XNOR U38745 ( .A(n34595), .B(n34599), .Z(n34880) );
  XNOR U38746 ( .A(n34590), .B(n34594), .Z(n34881) );
  XNOR U38747 ( .A(n34585), .B(n34589), .Z(n34882) );
  XNOR U38748 ( .A(n34580), .B(n34584), .Z(n34883) );
  XNOR U38749 ( .A(n34575), .B(n34579), .Z(n34884) );
  XNOR U38750 ( .A(n34570), .B(n34574), .Z(n34885) );
  XNOR U38751 ( .A(n34565), .B(n34569), .Z(n34886) );
  XNOR U38752 ( .A(n34560), .B(n34564), .Z(n34887) );
  XNOR U38753 ( .A(n34555), .B(n34559), .Z(n34888) );
  XNOR U38754 ( .A(n34550), .B(n34554), .Z(n34889) );
  XNOR U38755 ( .A(n34545), .B(n34549), .Z(n34890) );
  XNOR U38756 ( .A(n34540), .B(n34544), .Z(n34891) );
  XNOR U38757 ( .A(n34535), .B(n34539), .Z(n34892) );
  XNOR U38758 ( .A(n34530), .B(n34534), .Z(n34893) );
  XNOR U38759 ( .A(n34525), .B(n34529), .Z(n34894) );
  XNOR U38760 ( .A(n34520), .B(n34524), .Z(n34895) );
  XNOR U38761 ( .A(n34515), .B(n34519), .Z(n34896) );
  XNOR U38762 ( .A(n34510), .B(n34514), .Z(n34897) );
  XOR U38763 ( .A(n34898), .B(n34509), .Z(n34510) );
  AND U38764 ( .A(a[0]), .B(b[66]), .Z(n34898) );
  XNOR U38765 ( .A(n34899), .B(n34509), .Z(n34511) );
  XNOR U38766 ( .A(n34900), .B(n34901), .Z(n34509) );
  ANDN U38767 ( .B(n34902), .A(n34903), .Z(n34900) );
  AND U38768 ( .A(a[1]), .B(b[65]), .Z(n34899) );
  XOR U38769 ( .A(n34905), .B(n34906), .Z(n34514) );
  ANDN U38770 ( .B(n34907), .A(n34908), .Z(n34905) );
  AND U38771 ( .A(a[2]), .B(b[64]), .Z(n34904) );
  XOR U38772 ( .A(n34910), .B(n34911), .Z(n34519) );
  ANDN U38773 ( .B(n34912), .A(n34913), .Z(n34910) );
  AND U38774 ( .A(a[3]), .B(b[63]), .Z(n34909) );
  XOR U38775 ( .A(n34915), .B(n34916), .Z(n34524) );
  ANDN U38776 ( .B(n34917), .A(n34918), .Z(n34915) );
  AND U38777 ( .A(a[4]), .B(b[62]), .Z(n34914) );
  XOR U38778 ( .A(n34920), .B(n34921), .Z(n34529) );
  ANDN U38779 ( .B(n34922), .A(n34923), .Z(n34920) );
  AND U38780 ( .A(a[5]), .B(b[61]), .Z(n34919) );
  XOR U38781 ( .A(n34925), .B(n34926), .Z(n34534) );
  ANDN U38782 ( .B(n34927), .A(n34928), .Z(n34925) );
  AND U38783 ( .A(a[6]), .B(b[60]), .Z(n34924) );
  XOR U38784 ( .A(n34930), .B(n34931), .Z(n34539) );
  ANDN U38785 ( .B(n34932), .A(n34933), .Z(n34930) );
  AND U38786 ( .A(a[7]), .B(b[59]), .Z(n34929) );
  XOR U38787 ( .A(n34935), .B(n34936), .Z(n34544) );
  ANDN U38788 ( .B(n34937), .A(n34938), .Z(n34935) );
  AND U38789 ( .A(a[8]), .B(b[58]), .Z(n34934) );
  XOR U38790 ( .A(n34940), .B(n34941), .Z(n34549) );
  ANDN U38791 ( .B(n34942), .A(n34943), .Z(n34940) );
  AND U38792 ( .A(a[9]), .B(b[57]), .Z(n34939) );
  XOR U38793 ( .A(n34945), .B(n34946), .Z(n34554) );
  ANDN U38794 ( .B(n34947), .A(n34948), .Z(n34945) );
  AND U38795 ( .A(a[10]), .B(b[56]), .Z(n34944) );
  XOR U38796 ( .A(n34950), .B(n34951), .Z(n34559) );
  ANDN U38797 ( .B(n34952), .A(n34953), .Z(n34950) );
  AND U38798 ( .A(a[11]), .B(b[55]), .Z(n34949) );
  XOR U38799 ( .A(n34955), .B(n34956), .Z(n34564) );
  ANDN U38800 ( .B(n34957), .A(n34958), .Z(n34955) );
  AND U38801 ( .A(a[12]), .B(b[54]), .Z(n34954) );
  XOR U38802 ( .A(n34960), .B(n34961), .Z(n34569) );
  ANDN U38803 ( .B(n34962), .A(n34963), .Z(n34960) );
  AND U38804 ( .A(a[13]), .B(b[53]), .Z(n34959) );
  XOR U38805 ( .A(n34965), .B(n34966), .Z(n34574) );
  ANDN U38806 ( .B(n34967), .A(n34968), .Z(n34965) );
  AND U38807 ( .A(a[14]), .B(b[52]), .Z(n34964) );
  XOR U38808 ( .A(n34970), .B(n34971), .Z(n34579) );
  ANDN U38809 ( .B(n34972), .A(n34973), .Z(n34970) );
  AND U38810 ( .A(a[15]), .B(b[51]), .Z(n34969) );
  XOR U38811 ( .A(n34975), .B(n34976), .Z(n34584) );
  ANDN U38812 ( .B(n34977), .A(n34978), .Z(n34975) );
  AND U38813 ( .A(a[16]), .B(b[50]), .Z(n34974) );
  XOR U38814 ( .A(n34980), .B(n34981), .Z(n34589) );
  ANDN U38815 ( .B(n34982), .A(n34983), .Z(n34980) );
  AND U38816 ( .A(a[17]), .B(b[49]), .Z(n34979) );
  XOR U38817 ( .A(n34985), .B(n34986), .Z(n34594) );
  ANDN U38818 ( .B(n34987), .A(n34988), .Z(n34985) );
  AND U38819 ( .A(a[18]), .B(b[48]), .Z(n34984) );
  XOR U38820 ( .A(n34990), .B(n34991), .Z(n34599) );
  ANDN U38821 ( .B(n34992), .A(n34993), .Z(n34990) );
  AND U38822 ( .A(a[19]), .B(b[47]), .Z(n34989) );
  XOR U38823 ( .A(n34995), .B(n34996), .Z(n34604) );
  ANDN U38824 ( .B(n34997), .A(n34998), .Z(n34995) );
  AND U38825 ( .A(a[20]), .B(b[46]), .Z(n34994) );
  XOR U38826 ( .A(n35000), .B(n35001), .Z(n34609) );
  ANDN U38827 ( .B(n35002), .A(n35003), .Z(n35000) );
  AND U38828 ( .A(a[21]), .B(b[45]), .Z(n34999) );
  XOR U38829 ( .A(n35005), .B(n35006), .Z(n34614) );
  ANDN U38830 ( .B(n35007), .A(n35008), .Z(n35005) );
  AND U38831 ( .A(a[22]), .B(b[44]), .Z(n35004) );
  XOR U38832 ( .A(n35010), .B(n35011), .Z(n34619) );
  ANDN U38833 ( .B(n35012), .A(n35013), .Z(n35010) );
  AND U38834 ( .A(a[23]), .B(b[43]), .Z(n35009) );
  XOR U38835 ( .A(n35015), .B(n35016), .Z(n34624) );
  ANDN U38836 ( .B(n35017), .A(n35018), .Z(n35015) );
  AND U38837 ( .A(a[24]), .B(b[42]), .Z(n35014) );
  XOR U38838 ( .A(n35020), .B(n35021), .Z(n34629) );
  ANDN U38839 ( .B(n35022), .A(n35023), .Z(n35020) );
  AND U38840 ( .A(a[25]), .B(b[41]), .Z(n35019) );
  XOR U38841 ( .A(n35025), .B(n35026), .Z(n34634) );
  ANDN U38842 ( .B(n35027), .A(n35028), .Z(n35025) );
  AND U38843 ( .A(a[26]), .B(b[40]), .Z(n35024) );
  XOR U38844 ( .A(n35030), .B(n35031), .Z(n34639) );
  ANDN U38845 ( .B(n35032), .A(n35033), .Z(n35030) );
  AND U38846 ( .A(a[27]), .B(b[39]), .Z(n35029) );
  XOR U38847 ( .A(n35035), .B(n35036), .Z(n34644) );
  ANDN U38848 ( .B(n35037), .A(n35038), .Z(n35035) );
  AND U38849 ( .A(a[28]), .B(b[38]), .Z(n35034) );
  XOR U38850 ( .A(n35040), .B(n35041), .Z(n34649) );
  ANDN U38851 ( .B(n35042), .A(n35043), .Z(n35040) );
  AND U38852 ( .A(a[29]), .B(b[37]), .Z(n35039) );
  XOR U38853 ( .A(n35045), .B(n35046), .Z(n34654) );
  ANDN U38854 ( .B(n35047), .A(n35048), .Z(n35045) );
  AND U38855 ( .A(a[30]), .B(b[36]), .Z(n35044) );
  XOR U38856 ( .A(n35050), .B(n35051), .Z(n34659) );
  ANDN U38857 ( .B(n35052), .A(n35053), .Z(n35050) );
  AND U38858 ( .A(a[31]), .B(b[35]), .Z(n35049) );
  XOR U38859 ( .A(n35055), .B(n35056), .Z(n34664) );
  ANDN U38860 ( .B(n35057), .A(n35058), .Z(n35055) );
  AND U38861 ( .A(a[32]), .B(b[34]), .Z(n35054) );
  XOR U38862 ( .A(n35060), .B(n35061), .Z(n34669) );
  ANDN U38863 ( .B(n35062), .A(n35063), .Z(n35060) );
  AND U38864 ( .A(a[33]), .B(b[33]), .Z(n35059) );
  XOR U38865 ( .A(n35065), .B(n35066), .Z(n34674) );
  ANDN U38866 ( .B(n35067), .A(n35068), .Z(n35065) );
  AND U38867 ( .A(a[34]), .B(b[32]), .Z(n35064) );
  XOR U38868 ( .A(n35070), .B(n35071), .Z(n34679) );
  ANDN U38869 ( .B(n35072), .A(n35073), .Z(n35070) );
  AND U38870 ( .A(a[35]), .B(b[31]), .Z(n35069) );
  XOR U38871 ( .A(n35075), .B(n35076), .Z(n34684) );
  ANDN U38872 ( .B(n35077), .A(n35078), .Z(n35075) );
  AND U38873 ( .A(a[36]), .B(b[30]), .Z(n35074) );
  XOR U38874 ( .A(n35080), .B(n35081), .Z(n34689) );
  ANDN U38875 ( .B(n35082), .A(n35083), .Z(n35080) );
  AND U38876 ( .A(a[37]), .B(b[29]), .Z(n35079) );
  XOR U38877 ( .A(n35085), .B(n35086), .Z(n34694) );
  ANDN U38878 ( .B(n35087), .A(n35088), .Z(n35085) );
  AND U38879 ( .A(a[38]), .B(b[28]), .Z(n35084) );
  XOR U38880 ( .A(n35090), .B(n35091), .Z(n34699) );
  ANDN U38881 ( .B(n35092), .A(n35093), .Z(n35090) );
  AND U38882 ( .A(a[39]), .B(b[27]), .Z(n35089) );
  XOR U38883 ( .A(n35095), .B(n35096), .Z(n34704) );
  ANDN U38884 ( .B(n35097), .A(n35098), .Z(n35095) );
  AND U38885 ( .A(a[40]), .B(b[26]), .Z(n35094) );
  XOR U38886 ( .A(n35100), .B(n35101), .Z(n34709) );
  ANDN U38887 ( .B(n35102), .A(n35103), .Z(n35100) );
  AND U38888 ( .A(a[41]), .B(b[25]), .Z(n35099) );
  XOR U38889 ( .A(n35105), .B(n35106), .Z(n34714) );
  ANDN U38890 ( .B(n35107), .A(n35108), .Z(n35105) );
  AND U38891 ( .A(a[42]), .B(b[24]), .Z(n35104) );
  XOR U38892 ( .A(n35110), .B(n35111), .Z(n34719) );
  ANDN U38893 ( .B(n35112), .A(n35113), .Z(n35110) );
  AND U38894 ( .A(a[43]), .B(b[23]), .Z(n35109) );
  XOR U38895 ( .A(n35115), .B(n35116), .Z(n34724) );
  ANDN U38896 ( .B(n35117), .A(n35118), .Z(n35115) );
  AND U38897 ( .A(a[44]), .B(b[22]), .Z(n35114) );
  XOR U38898 ( .A(n35120), .B(n35121), .Z(n34729) );
  ANDN U38899 ( .B(n35122), .A(n35123), .Z(n35120) );
  AND U38900 ( .A(a[45]), .B(b[21]), .Z(n35119) );
  XOR U38901 ( .A(n35125), .B(n35126), .Z(n34734) );
  ANDN U38902 ( .B(n35127), .A(n35128), .Z(n35125) );
  AND U38903 ( .A(a[46]), .B(b[20]), .Z(n35124) );
  XOR U38904 ( .A(n35130), .B(n35131), .Z(n34739) );
  ANDN U38905 ( .B(n35132), .A(n35133), .Z(n35130) );
  AND U38906 ( .A(a[47]), .B(b[19]), .Z(n35129) );
  XOR U38907 ( .A(n35135), .B(n35136), .Z(n34744) );
  ANDN U38908 ( .B(n35137), .A(n35138), .Z(n35135) );
  AND U38909 ( .A(a[48]), .B(b[18]), .Z(n35134) );
  XOR U38910 ( .A(n35140), .B(n35141), .Z(n34749) );
  ANDN U38911 ( .B(n35142), .A(n35143), .Z(n35140) );
  AND U38912 ( .A(a[49]), .B(b[17]), .Z(n35139) );
  XOR U38913 ( .A(n35145), .B(n35146), .Z(n34754) );
  ANDN U38914 ( .B(n35147), .A(n35148), .Z(n35145) );
  AND U38915 ( .A(a[50]), .B(b[16]), .Z(n35144) );
  XOR U38916 ( .A(n35150), .B(n35151), .Z(n34759) );
  ANDN U38917 ( .B(n35152), .A(n35153), .Z(n35150) );
  AND U38918 ( .A(a[51]), .B(b[15]), .Z(n35149) );
  XOR U38919 ( .A(n35155), .B(n35156), .Z(n34764) );
  ANDN U38920 ( .B(n35157), .A(n35158), .Z(n35155) );
  AND U38921 ( .A(a[52]), .B(b[14]), .Z(n35154) );
  XOR U38922 ( .A(n35160), .B(n35161), .Z(n34769) );
  ANDN U38923 ( .B(n35162), .A(n35163), .Z(n35160) );
  AND U38924 ( .A(a[53]), .B(b[13]), .Z(n35159) );
  XOR U38925 ( .A(n35165), .B(n35166), .Z(n34774) );
  ANDN U38926 ( .B(n35167), .A(n35168), .Z(n35165) );
  AND U38927 ( .A(a[54]), .B(b[12]), .Z(n35164) );
  XOR U38928 ( .A(n35170), .B(n35171), .Z(n34779) );
  ANDN U38929 ( .B(n35172), .A(n35173), .Z(n35170) );
  AND U38930 ( .A(a[55]), .B(b[11]), .Z(n35169) );
  XOR U38931 ( .A(n35175), .B(n35176), .Z(n34784) );
  ANDN U38932 ( .B(n35177), .A(n35178), .Z(n35175) );
  AND U38933 ( .A(a[56]), .B(b[10]), .Z(n35174) );
  XOR U38934 ( .A(n35180), .B(n35181), .Z(n34789) );
  ANDN U38935 ( .B(n35182), .A(n35183), .Z(n35180) );
  AND U38936 ( .A(b[9]), .B(a[57]), .Z(n35179) );
  XOR U38937 ( .A(n35185), .B(n35186), .Z(n34794) );
  ANDN U38938 ( .B(n35187), .A(n35188), .Z(n35185) );
  AND U38939 ( .A(b[8]), .B(a[58]), .Z(n35184) );
  XOR U38940 ( .A(n35190), .B(n35191), .Z(n34799) );
  ANDN U38941 ( .B(n35192), .A(n35193), .Z(n35190) );
  AND U38942 ( .A(b[7]), .B(a[59]), .Z(n35189) );
  XOR U38943 ( .A(n35195), .B(n35196), .Z(n34804) );
  ANDN U38944 ( .B(n35197), .A(n35198), .Z(n35195) );
  AND U38945 ( .A(b[6]), .B(a[60]), .Z(n35194) );
  XOR U38946 ( .A(n35200), .B(n35201), .Z(n34809) );
  ANDN U38947 ( .B(n35202), .A(n35203), .Z(n35200) );
  AND U38948 ( .A(b[5]), .B(a[61]), .Z(n35199) );
  XOR U38949 ( .A(n35205), .B(n35206), .Z(n34814) );
  ANDN U38950 ( .B(n35207), .A(n35208), .Z(n35205) );
  AND U38951 ( .A(b[4]), .B(a[62]), .Z(n35204) );
  XOR U38952 ( .A(n35210), .B(n35211), .Z(n34819) );
  ANDN U38953 ( .B(n34831), .A(n34832), .Z(n35210) );
  AND U38954 ( .A(b[2]), .B(a[63]), .Z(n35212) );
  XNOR U38955 ( .A(n35207), .B(n35211), .Z(n35213) );
  XOR U38956 ( .A(n35214), .B(n35215), .Z(n35211) );
  OR U38957 ( .A(n34834), .B(n34835), .Z(n35215) );
  XNOR U38958 ( .A(n35217), .B(n35218), .Z(n35216) );
  XOR U38959 ( .A(n35217), .B(n35220), .Z(n34834) );
  NAND U38960 ( .A(b[1]), .B(a[63]), .Z(n35220) );
  IV U38961 ( .A(n35214), .Z(n35217) );
  NANDN U38962 ( .A(n81), .B(n82), .Z(n35214) );
  XOR U38963 ( .A(n35221), .B(n35222), .Z(n82) );
  NAND U38964 ( .A(a[63]), .B(b[0]), .Z(n81) );
  XNOR U38965 ( .A(n35202), .B(n35206), .Z(n35223) );
  XNOR U38966 ( .A(n35197), .B(n35201), .Z(n35224) );
  XNOR U38967 ( .A(n35192), .B(n35196), .Z(n35225) );
  XNOR U38968 ( .A(n35187), .B(n35191), .Z(n35226) );
  XNOR U38969 ( .A(n35182), .B(n35186), .Z(n35227) );
  XNOR U38970 ( .A(n35177), .B(n35181), .Z(n35228) );
  XNOR U38971 ( .A(n35172), .B(n35176), .Z(n35229) );
  XNOR U38972 ( .A(n35167), .B(n35171), .Z(n35230) );
  XNOR U38973 ( .A(n35162), .B(n35166), .Z(n35231) );
  XNOR U38974 ( .A(n35157), .B(n35161), .Z(n35232) );
  XNOR U38975 ( .A(n35152), .B(n35156), .Z(n35233) );
  XNOR U38976 ( .A(n35147), .B(n35151), .Z(n35234) );
  XNOR U38977 ( .A(n35142), .B(n35146), .Z(n35235) );
  XNOR U38978 ( .A(n35137), .B(n35141), .Z(n35236) );
  XNOR U38979 ( .A(n35132), .B(n35136), .Z(n35237) );
  XNOR U38980 ( .A(n35127), .B(n35131), .Z(n35238) );
  XNOR U38981 ( .A(n35122), .B(n35126), .Z(n35239) );
  XNOR U38982 ( .A(n35117), .B(n35121), .Z(n35240) );
  XNOR U38983 ( .A(n35112), .B(n35116), .Z(n35241) );
  XNOR U38984 ( .A(n35107), .B(n35111), .Z(n35242) );
  XNOR U38985 ( .A(n35102), .B(n35106), .Z(n35243) );
  XNOR U38986 ( .A(n35097), .B(n35101), .Z(n35244) );
  XNOR U38987 ( .A(n35092), .B(n35096), .Z(n35245) );
  XNOR U38988 ( .A(n35087), .B(n35091), .Z(n35246) );
  XNOR U38989 ( .A(n35082), .B(n35086), .Z(n35247) );
  XNOR U38990 ( .A(n35077), .B(n35081), .Z(n35248) );
  XNOR U38991 ( .A(n35072), .B(n35076), .Z(n35249) );
  XNOR U38992 ( .A(n35067), .B(n35071), .Z(n35250) );
  XNOR U38993 ( .A(n35062), .B(n35066), .Z(n35251) );
  XNOR U38994 ( .A(n35057), .B(n35061), .Z(n35252) );
  XNOR U38995 ( .A(n35052), .B(n35056), .Z(n35253) );
  XNOR U38996 ( .A(n35047), .B(n35051), .Z(n35254) );
  XNOR U38997 ( .A(n35042), .B(n35046), .Z(n35255) );
  XNOR U38998 ( .A(n35037), .B(n35041), .Z(n35256) );
  XNOR U38999 ( .A(n35032), .B(n35036), .Z(n35257) );
  XNOR U39000 ( .A(n35027), .B(n35031), .Z(n35258) );
  XNOR U39001 ( .A(n35022), .B(n35026), .Z(n35259) );
  XNOR U39002 ( .A(n35017), .B(n35021), .Z(n35260) );
  XNOR U39003 ( .A(n35012), .B(n35016), .Z(n35261) );
  XNOR U39004 ( .A(n35007), .B(n35011), .Z(n35262) );
  XNOR U39005 ( .A(n35002), .B(n35006), .Z(n35263) );
  XNOR U39006 ( .A(n34997), .B(n35001), .Z(n35264) );
  XNOR U39007 ( .A(n34992), .B(n34996), .Z(n35265) );
  XNOR U39008 ( .A(n34987), .B(n34991), .Z(n35266) );
  XNOR U39009 ( .A(n34982), .B(n34986), .Z(n35267) );
  XNOR U39010 ( .A(n34977), .B(n34981), .Z(n35268) );
  XNOR U39011 ( .A(n34972), .B(n34976), .Z(n35269) );
  XNOR U39012 ( .A(n34967), .B(n34971), .Z(n35270) );
  XNOR U39013 ( .A(n34962), .B(n34966), .Z(n35271) );
  XNOR U39014 ( .A(n34957), .B(n34961), .Z(n35272) );
  XNOR U39015 ( .A(n34952), .B(n34956), .Z(n35273) );
  XNOR U39016 ( .A(n34947), .B(n34951), .Z(n35274) );
  XNOR U39017 ( .A(n34942), .B(n34946), .Z(n35275) );
  XNOR U39018 ( .A(n34937), .B(n34941), .Z(n35276) );
  XNOR U39019 ( .A(n34932), .B(n34936), .Z(n35277) );
  XNOR U39020 ( .A(n34927), .B(n34931), .Z(n35278) );
  XNOR U39021 ( .A(n34922), .B(n34926), .Z(n35279) );
  XNOR U39022 ( .A(n34917), .B(n34921), .Z(n35280) );
  XNOR U39023 ( .A(n34912), .B(n34916), .Z(n35281) );
  XNOR U39024 ( .A(n34907), .B(n34911), .Z(n35282) );
  XNOR U39025 ( .A(n34902), .B(n34906), .Z(n35283) );
  XNOR U39026 ( .A(n35284), .B(n34901), .Z(n34902) );
  AND U39027 ( .A(a[0]), .B(b[65]), .Z(n35284) );
  XOR U39028 ( .A(n35285), .B(n34901), .Z(n34903) );
  XNOR U39029 ( .A(n35286), .B(n35287), .Z(n34901) );
  ANDN U39030 ( .B(n35288), .A(n35289), .Z(n35286) );
  AND U39031 ( .A(a[1]), .B(b[64]), .Z(n35285) );
  XOR U39032 ( .A(n35291), .B(n35292), .Z(n34906) );
  ANDN U39033 ( .B(n35293), .A(n35294), .Z(n35291) );
  AND U39034 ( .A(a[2]), .B(b[63]), .Z(n35290) );
  XOR U39035 ( .A(n35296), .B(n35297), .Z(n34911) );
  ANDN U39036 ( .B(n35298), .A(n35299), .Z(n35296) );
  AND U39037 ( .A(a[3]), .B(b[62]), .Z(n35295) );
  XOR U39038 ( .A(n35301), .B(n35302), .Z(n34916) );
  ANDN U39039 ( .B(n35303), .A(n35304), .Z(n35301) );
  AND U39040 ( .A(a[4]), .B(b[61]), .Z(n35300) );
  XOR U39041 ( .A(n35306), .B(n35307), .Z(n34921) );
  ANDN U39042 ( .B(n35308), .A(n35309), .Z(n35306) );
  AND U39043 ( .A(a[5]), .B(b[60]), .Z(n35305) );
  XOR U39044 ( .A(n35311), .B(n35312), .Z(n34926) );
  ANDN U39045 ( .B(n35313), .A(n35314), .Z(n35311) );
  AND U39046 ( .A(a[6]), .B(b[59]), .Z(n35310) );
  XOR U39047 ( .A(n35316), .B(n35317), .Z(n34931) );
  ANDN U39048 ( .B(n35318), .A(n35319), .Z(n35316) );
  AND U39049 ( .A(a[7]), .B(b[58]), .Z(n35315) );
  XOR U39050 ( .A(n35321), .B(n35322), .Z(n34936) );
  ANDN U39051 ( .B(n35323), .A(n35324), .Z(n35321) );
  AND U39052 ( .A(a[8]), .B(b[57]), .Z(n35320) );
  XOR U39053 ( .A(n35326), .B(n35327), .Z(n34941) );
  ANDN U39054 ( .B(n35328), .A(n35329), .Z(n35326) );
  AND U39055 ( .A(a[9]), .B(b[56]), .Z(n35325) );
  XOR U39056 ( .A(n35331), .B(n35332), .Z(n34946) );
  ANDN U39057 ( .B(n35333), .A(n35334), .Z(n35331) );
  AND U39058 ( .A(a[10]), .B(b[55]), .Z(n35330) );
  XOR U39059 ( .A(n35336), .B(n35337), .Z(n34951) );
  ANDN U39060 ( .B(n35338), .A(n35339), .Z(n35336) );
  AND U39061 ( .A(a[11]), .B(b[54]), .Z(n35335) );
  XOR U39062 ( .A(n35341), .B(n35342), .Z(n34956) );
  ANDN U39063 ( .B(n35343), .A(n35344), .Z(n35341) );
  AND U39064 ( .A(a[12]), .B(b[53]), .Z(n35340) );
  XOR U39065 ( .A(n35346), .B(n35347), .Z(n34961) );
  ANDN U39066 ( .B(n35348), .A(n35349), .Z(n35346) );
  AND U39067 ( .A(a[13]), .B(b[52]), .Z(n35345) );
  XOR U39068 ( .A(n35351), .B(n35352), .Z(n34966) );
  ANDN U39069 ( .B(n35353), .A(n35354), .Z(n35351) );
  AND U39070 ( .A(a[14]), .B(b[51]), .Z(n35350) );
  XOR U39071 ( .A(n35356), .B(n35357), .Z(n34971) );
  ANDN U39072 ( .B(n35358), .A(n35359), .Z(n35356) );
  AND U39073 ( .A(a[15]), .B(b[50]), .Z(n35355) );
  XOR U39074 ( .A(n35361), .B(n35362), .Z(n34976) );
  ANDN U39075 ( .B(n35363), .A(n35364), .Z(n35361) );
  AND U39076 ( .A(a[16]), .B(b[49]), .Z(n35360) );
  XOR U39077 ( .A(n35366), .B(n35367), .Z(n34981) );
  ANDN U39078 ( .B(n35368), .A(n35369), .Z(n35366) );
  AND U39079 ( .A(a[17]), .B(b[48]), .Z(n35365) );
  XOR U39080 ( .A(n35371), .B(n35372), .Z(n34986) );
  ANDN U39081 ( .B(n35373), .A(n35374), .Z(n35371) );
  AND U39082 ( .A(a[18]), .B(b[47]), .Z(n35370) );
  XOR U39083 ( .A(n35376), .B(n35377), .Z(n34991) );
  ANDN U39084 ( .B(n35378), .A(n35379), .Z(n35376) );
  AND U39085 ( .A(a[19]), .B(b[46]), .Z(n35375) );
  XOR U39086 ( .A(n35381), .B(n35382), .Z(n34996) );
  ANDN U39087 ( .B(n35383), .A(n35384), .Z(n35381) );
  AND U39088 ( .A(a[20]), .B(b[45]), .Z(n35380) );
  XOR U39089 ( .A(n35386), .B(n35387), .Z(n35001) );
  ANDN U39090 ( .B(n35388), .A(n35389), .Z(n35386) );
  AND U39091 ( .A(a[21]), .B(b[44]), .Z(n35385) );
  XOR U39092 ( .A(n35391), .B(n35392), .Z(n35006) );
  ANDN U39093 ( .B(n35393), .A(n35394), .Z(n35391) );
  AND U39094 ( .A(a[22]), .B(b[43]), .Z(n35390) );
  XOR U39095 ( .A(n35396), .B(n35397), .Z(n35011) );
  ANDN U39096 ( .B(n35398), .A(n35399), .Z(n35396) );
  AND U39097 ( .A(a[23]), .B(b[42]), .Z(n35395) );
  XOR U39098 ( .A(n35401), .B(n35402), .Z(n35016) );
  ANDN U39099 ( .B(n35403), .A(n35404), .Z(n35401) );
  AND U39100 ( .A(a[24]), .B(b[41]), .Z(n35400) );
  XOR U39101 ( .A(n35406), .B(n35407), .Z(n35021) );
  ANDN U39102 ( .B(n35408), .A(n35409), .Z(n35406) );
  AND U39103 ( .A(a[25]), .B(b[40]), .Z(n35405) );
  XOR U39104 ( .A(n35411), .B(n35412), .Z(n35026) );
  ANDN U39105 ( .B(n35413), .A(n35414), .Z(n35411) );
  AND U39106 ( .A(a[26]), .B(b[39]), .Z(n35410) );
  XOR U39107 ( .A(n35416), .B(n35417), .Z(n35031) );
  ANDN U39108 ( .B(n35418), .A(n35419), .Z(n35416) );
  AND U39109 ( .A(a[27]), .B(b[38]), .Z(n35415) );
  XOR U39110 ( .A(n35421), .B(n35422), .Z(n35036) );
  ANDN U39111 ( .B(n35423), .A(n35424), .Z(n35421) );
  AND U39112 ( .A(a[28]), .B(b[37]), .Z(n35420) );
  XOR U39113 ( .A(n35426), .B(n35427), .Z(n35041) );
  ANDN U39114 ( .B(n35428), .A(n35429), .Z(n35426) );
  AND U39115 ( .A(a[29]), .B(b[36]), .Z(n35425) );
  XOR U39116 ( .A(n35431), .B(n35432), .Z(n35046) );
  ANDN U39117 ( .B(n35433), .A(n35434), .Z(n35431) );
  AND U39118 ( .A(a[30]), .B(b[35]), .Z(n35430) );
  XOR U39119 ( .A(n35436), .B(n35437), .Z(n35051) );
  ANDN U39120 ( .B(n35438), .A(n35439), .Z(n35436) );
  AND U39121 ( .A(a[31]), .B(b[34]), .Z(n35435) );
  XOR U39122 ( .A(n35441), .B(n35442), .Z(n35056) );
  ANDN U39123 ( .B(n35443), .A(n35444), .Z(n35441) );
  AND U39124 ( .A(a[32]), .B(b[33]), .Z(n35440) );
  XOR U39125 ( .A(n35446), .B(n35447), .Z(n35061) );
  ANDN U39126 ( .B(n35448), .A(n35449), .Z(n35446) );
  AND U39127 ( .A(a[33]), .B(b[32]), .Z(n35445) );
  XOR U39128 ( .A(n35451), .B(n35452), .Z(n35066) );
  ANDN U39129 ( .B(n35453), .A(n35454), .Z(n35451) );
  AND U39130 ( .A(a[34]), .B(b[31]), .Z(n35450) );
  XOR U39131 ( .A(n35456), .B(n35457), .Z(n35071) );
  ANDN U39132 ( .B(n35458), .A(n35459), .Z(n35456) );
  AND U39133 ( .A(a[35]), .B(b[30]), .Z(n35455) );
  XOR U39134 ( .A(n35461), .B(n35462), .Z(n35076) );
  ANDN U39135 ( .B(n35463), .A(n35464), .Z(n35461) );
  AND U39136 ( .A(a[36]), .B(b[29]), .Z(n35460) );
  XOR U39137 ( .A(n35466), .B(n35467), .Z(n35081) );
  ANDN U39138 ( .B(n35468), .A(n35469), .Z(n35466) );
  AND U39139 ( .A(a[37]), .B(b[28]), .Z(n35465) );
  XOR U39140 ( .A(n35471), .B(n35472), .Z(n35086) );
  ANDN U39141 ( .B(n35473), .A(n35474), .Z(n35471) );
  AND U39142 ( .A(a[38]), .B(b[27]), .Z(n35470) );
  XOR U39143 ( .A(n35476), .B(n35477), .Z(n35091) );
  ANDN U39144 ( .B(n35478), .A(n35479), .Z(n35476) );
  AND U39145 ( .A(a[39]), .B(b[26]), .Z(n35475) );
  XOR U39146 ( .A(n35481), .B(n35482), .Z(n35096) );
  ANDN U39147 ( .B(n35483), .A(n35484), .Z(n35481) );
  AND U39148 ( .A(a[40]), .B(b[25]), .Z(n35480) );
  XOR U39149 ( .A(n35486), .B(n35487), .Z(n35101) );
  ANDN U39150 ( .B(n35488), .A(n35489), .Z(n35486) );
  AND U39151 ( .A(a[41]), .B(b[24]), .Z(n35485) );
  XOR U39152 ( .A(n35491), .B(n35492), .Z(n35106) );
  ANDN U39153 ( .B(n35493), .A(n35494), .Z(n35491) );
  AND U39154 ( .A(a[42]), .B(b[23]), .Z(n35490) );
  XOR U39155 ( .A(n35496), .B(n35497), .Z(n35111) );
  ANDN U39156 ( .B(n35498), .A(n35499), .Z(n35496) );
  AND U39157 ( .A(a[43]), .B(b[22]), .Z(n35495) );
  XOR U39158 ( .A(n35501), .B(n35502), .Z(n35116) );
  ANDN U39159 ( .B(n35503), .A(n35504), .Z(n35501) );
  AND U39160 ( .A(a[44]), .B(b[21]), .Z(n35500) );
  XOR U39161 ( .A(n35506), .B(n35507), .Z(n35121) );
  ANDN U39162 ( .B(n35508), .A(n35509), .Z(n35506) );
  AND U39163 ( .A(a[45]), .B(b[20]), .Z(n35505) );
  XOR U39164 ( .A(n35511), .B(n35512), .Z(n35126) );
  ANDN U39165 ( .B(n35513), .A(n35514), .Z(n35511) );
  AND U39166 ( .A(a[46]), .B(b[19]), .Z(n35510) );
  XOR U39167 ( .A(n35516), .B(n35517), .Z(n35131) );
  ANDN U39168 ( .B(n35518), .A(n35519), .Z(n35516) );
  AND U39169 ( .A(a[47]), .B(b[18]), .Z(n35515) );
  XOR U39170 ( .A(n35521), .B(n35522), .Z(n35136) );
  ANDN U39171 ( .B(n35523), .A(n35524), .Z(n35521) );
  AND U39172 ( .A(a[48]), .B(b[17]), .Z(n35520) );
  XOR U39173 ( .A(n35526), .B(n35527), .Z(n35141) );
  ANDN U39174 ( .B(n35528), .A(n35529), .Z(n35526) );
  AND U39175 ( .A(a[49]), .B(b[16]), .Z(n35525) );
  XOR U39176 ( .A(n35531), .B(n35532), .Z(n35146) );
  ANDN U39177 ( .B(n35533), .A(n35534), .Z(n35531) );
  AND U39178 ( .A(a[50]), .B(b[15]), .Z(n35530) );
  XOR U39179 ( .A(n35536), .B(n35537), .Z(n35151) );
  ANDN U39180 ( .B(n35538), .A(n35539), .Z(n35536) );
  AND U39181 ( .A(a[51]), .B(b[14]), .Z(n35535) );
  XOR U39182 ( .A(n35541), .B(n35542), .Z(n35156) );
  ANDN U39183 ( .B(n35543), .A(n35544), .Z(n35541) );
  AND U39184 ( .A(a[52]), .B(b[13]), .Z(n35540) );
  XOR U39185 ( .A(n35546), .B(n35547), .Z(n35161) );
  ANDN U39186 ( .B(n35548), .A(n35549), .Z(n35546) );
  AND U39187 ( .A(a[53]), .B(b[12]), .Z(n35545) );
  XOR U39188 ( .A(n35551), .B(n35552), .Z(n35166) );
  ANDN U39189 ( .B(n35553), .A(n35554), .Z(n35551) );
  AND U39190 ( .A(a[54]), .B(b[11]), .Z(n35550) );
  XOR U39191 ( .A(n35556), .B(n35557), .Z(n35171) );
  ANDN U39192 ( .B(n35558), .A(n35559), .Z(n35556) );
  AND U39193 ( .A(a[55]), .B(b[10]), .Z(n35555) );
  XOR U39194 ( .A(n35561), .B(n35562), .Z(n35176) );
  ANDN U39195 ( .B(n35563), .A(n35564), .Z(n35561) );
  AND U39196 ( .A(b[9]), .B(a[56]), .Z(n35560) );
  XOR U39197 ( .A(n35566), .B(n35567), .Z(n35181) );
  ANDN U39198 ( .B(n35568), .A(n35569), .Z(n35566) );
  AND U39199 ( .A(b[8]), .B(a[57]), .Z(n35565) );
  XOR U39200 ( .A(n35571), .B(n35572), .Z(n35186) );
  ANDN U39201 ( .B(n35573), .A(n35574), .Z(n35571) );
  AND U39202 ( .A(b[7]), .B(a[58]), .Z(n35570) );
  XOR U39203 ( .A(n35576), .B(n35577), .Z(n35191) );
  ANDN U39204 ( .B(n35578), .A(n35579), .Z(n35576) );
  AND U39205 ( .A(b[6]), .B(a[59]), .Z(n35575) );
  XOR U39206 ( .A(n35581), .B(n35582), .Z(n35196) );
  ANDN U39207 ( .B(n35583), .A(n35584), .Z(n35581) );
  AND U39208 ( .A(b[5]), .B(a[60]), .Z(n35580) );
  XOR U39209 ( .A(n35586), .B(n35587), .Z(n35201) );
  ANDN U39210 ( .B(n35588), .A(n35589), .Z(n35586) );
  AND U39211 ( .A(b[4]), .B(a[61]), .Z(n35585) );
  XOR U39212 ( .A(n35591), .B(n35592), .Z(n35206) );
  ANDN U39213 ( .B(n35218), .A(n35219), .Z(n35591) );
  AND U39214 ( .A(b[2]), .B(a[62]), .Z(n35593) );
  XNOR U39215 ( .A(n35588), .B(n35592), .Z(n35594) );
  XOR U39216 ( .A(n35595), .B(n35596), .Z(n35592) );
  OR U39217 ( .A(n35221), .B(n35222), .Z(n35596) );
  XNOR U39218 ( .A(n35598), .B(n35599), .Z(n35597) );
  XOR U39219 ( .A(n35598), .B(n35601), .Z(n35221) );
  NAND U39220 ( .A(b[1]), .B(a[62]), .Z(n35601) );
  IV U39221 ( .A(n35595), .Z(n35598) );
  NANDN U39222 ( .A(n83), .B(n84), .Z(n35595) );
  XOR U39223 ( .A(n35602), .B(n35603), .Z(n84) );
  NAND U39224 ( .A(a[62]), .B(b[0]), .Z(n83) );
  XNOR U39225 ( .A(n35583), .B(n35587), .Z(n35604) );
  XNOR U39226 ( .A(n35578), .B(n35582), .Z(n35605) );
  XNOR U39227 ( .A(n35573), .B(n35577), .Z(n35606) );
  XNOR U39228 ( .A(n35568), .B(n35572), .Z(n35607) );
  XNOR U39229 ( .A(n35563), .B(n35567), .Z(n35608) );
  XNOR U39230 ( .A(n35558), .B(n35562), .Z(n35609) );
  XNOR U39231 ( .A(n35553), .B(n35557), .Z(n35610) );
  XNOR U39232 ( .A(n35548), .B(n35552), .Z(n35611) );
  XNOR U39233 ( .A(n35543), .B(n35547), .Z(n35612) );
  XNOR U39234 ( .A(n35538), .B(n35542), .Z(n35613) );
  XNOR U39235 ( .A(n35533), .B(n35537), .Z(n35614) );
  XNOR U39236 ( .A(n35528), .B(n35532), .Z(n35615) );
  XNOR U39237 ( .A(n35523), .B(n35527), .Z(n35616) );
  XNOR U39238 ( .A(n35518), .B(n35522), .Z(n35617) );
  XNOR U39239 ( .A(n35513), .B(n35517), .Z(n35618) );
  XNOR U39240 ( .A(n35508), .B(n35512), .Z(n35619) );
  XNOR U39241 ( .A(n35503), .B(n35507), .Z(n35620) );
  XNOR U39242 ( .A(n35498), .B(n35502), .Z(n35621) );
  XNOR U39243 ( .A(n35493), .B(n35497), .Z(n35622) );
  XNOR U39244 ( .A(n35488), .B(n35492), .Z(n35623) );
  XNOR U39245 ( .A(n35483), .B(n35487), .Z(n35624) );
  XNOR U39246 ( .A(n35478), .B(n35482), .Z(n35625) );
  XNOR U39247 ( .A(n35473), .B(n35477), .Z(n35626) );
  XNOR U39248 ( .A(n35468), .B(n35472), .Z(n35627) );
  XNOR U39249 ( .A(n35463), .B(n35467), .Z(n35628) );
  XNOR U39250 ( .A(n35458), .B(n35462), .Z(n35629) );
  XNOR U39251 ( .A(n35453), .B(n35457), .Z(n35630) );
  XNOR U39252 ( .A(n35448), .B(n35452), .Z(n35631) );
  XNOR U39253 ( .A(n35443), .B(n35447), .Z(n35632) );
  XNOR U39254 ( .A(n35438), .B(n35442), .Z(n35633) );
  XNOR U39255 ( .A(n35433), .B(n35437), .Z(n35634) );
  XNOR U39256 ( .A(n35428), .B(n35432), .Z(n35635) );
  XNOR U39257 ( .A(n35423), .B(n35427), .Z(n35636) );
  XNOR U39258 ( .A(n35418), .B(n35422), .Z(n35637) );
  XNOR U39259 ( .A(n35413), .B(n35417), .Z(n35638) );
  XNOR U39260 ( .A(n35408), .B(n35412), .Z(n35639) );
  XNOR U39261 ( .A(n35403), .B(n35407), .Z(n35640) );
  XNOR U39262 ( .A(n35398), .B(n35402), .Z(n35641) );
  XNOR U39263 ( .A(n35393), .B(n35397), .Z(n35642) );
  XNOR U39264 ( .A(n35388), .B(n35392), .Z(n35643) );
  XNOR U39265 ( .A(n35383), .B(n35387), .Z(n35644) );
  XNOR U39266 ( .A(n35378), .B(n35382), .Z(n35645) );
  XNOR U39267 ( .A(n35373), .B(n35377), .Z(n35646) );
  XNOR U39268 ( .A(n35368), .B(n35372), .Z(n35647) );
  XNOR U39269 ( .A(n35363), .B(n35367), .Z(n35648) );
  XNOR U39270 ( .A(n35358), .B(n35362), .Z(n35649) );
  XNOR U39271 ( .A(n35353), .B(n35357), .Z(n35650) );
  XNOR U39272 ( .A(n35348), .B(n35352), .Z(n35651) );
  XNOR U39273 ( .A(n35343), .B(n35347), .Z(n35652) );
  XNOR U39274 ( .A(n35338), .B(n35342), .Z(n35653) );
  XNOR U39275 ( .A(n35333), .B(n35337), .Z(n35654) );
  XNOR U39276 ( .A(n35328), .B(n35332), .Z(n35655) );
  XNOR U39277 ( .A(n35323), .B(n35327), .Z(n35656) );
  XNOR U39278 ( .A(n35318), .B(n35322), .Z(n35657) );
  XNOR U39279 ( .A(n35313), .B(n35317), .Z(n35658) );
  XNOR U39280 ( .A(n35308), .B(n35312), .Z(n35659) );
  XNOR U39281 ( .A(n35303), .B(n35307), .Z(n35660) );
  XNOR U39282 ( .A(n35298), .B(n35302), .Z(n35661) );
  XNOR U39283 ( .A(n35293), .B(n35297), .Z(n35662) );
  XNOR U39284 ( .A(n35288), .B(n35292), .Z(n35663) );
  XOR U39285 ( .A(n35664), .B(n35287), .Z(n35288) );
  AND U39286 ( .A(a[0]), .B(b[64]), .Z(n35664) );
  XNOR U39287 ( .A(n35665), .B(n35287), .Z(n35289) );
  XNOR U39288 ( .A(n35666), .B(n35667), .Z(n35287) );
  ANDN U39289 ( .B(n35668), .A(n35669), .Z(n35666) );
  AND U39290 ( .A(a[1]), .B(b[63]), .Z(n35665) );
  XOR U39291 ( .A(n35671), .B(n35672), .Z(n35292) );
  ANDN U39292 ( .B(n35673), .A(n35674), .Z(n35671) );
  AND U39293 ( .A(a[2]), .B(b[62]), .Z(n35670) );
  XOR U39294 ( .A(n35676), .B(n35677), .Z(n35297) );
  ANDN U39295 ( .B(n35678), .A(n35679), .Z(n35676) );
  AND U39296 ( .A(a[3]), .B(b[61]), .Z(n35675) );
  XOR U39297 ( .A(n35681), .B(n35682), .Z(n35302) );
  ANDN U39298 ( .B(n35683), .A(n35684), .Z(n35681) );
  AND U39299 ( .A(a[4]), .B(b[60]), .Z(n35680) );
  XOR U39300 ( .A(n35686), .B(n35687), .Z(n35307) );
  ANDN U39301 ( .B(n35688), .A(n35689), .Z(n35686) );
  AND U39302 ( .A(a[5]), .B(b[59]), .Z(n35685) );
  XOR U39303 ( .A(n35691), .B(n35692), .Z(n35312) );
  ANDN U39304 ( .B(n35693), .A(n35694), .Z(n35691) );
  AND U39305 ( .A(a[6]), .B(b[58]), .Z(n35690) );
  XOR U39306 ( .A(n35696), .B(n35697), .Z(n35317) );
  ANDN U39307 ( .B(n35698), .A(n35699), .Z(n35696) );
  AND U39308 ( .A(a[7]), .B(b[57]), .Z(n35695) );
  XOR U39309 ( .A(n35701), .B(n35702), .Z(n35322) );
  ANDN U39310 ( .B(n35703), .A(n35704), .Z(n35701) );
  AND U39311 ( .A(a[8]), .B(b[56]), .Z(n35700) );
  XOR U39312 ( .A(n35706), .B(n35707), .Z(n35327) );
  ANDN U39313 ( .B(n35708), .A(n35709), .Z(n35706) );
  AND U39314 ( .A(a[9]), .B(b[55]), .Z(n35705) );
  XOR U39315 ( .A(n35711), .B(n35712), .Z(n35332) );
  ANDN U39316 ( .B(n35713), .A(n35714), .Z(n35711) );
  AND U39317 ( .A(a[10]), .B(b[54]), .Z(n35710) );
  XOR U39318 ( .A(n35716), .B(n35717), .Z(n35337) );
  ANDN U39319 ( .B(n35718), .A(n35719), .Z(n35716) );
  AND U39320 ( .A(a[11]), .B(b[53]), .Z(n35715) );
  XOR U39321 ( .A(n35721), .B(n35722), .Z(n35342) );
  ANDN U39322 ( .B(n35723), .A(n35724), .Z(n35721) );
  AND U39323 ( .A(a[12]), .B(b[52]), .Z(n35720) );
  XOR U39324 ( .A(n35726), .B(n35727), .Z(n35347) );
  ANDN U39325 ( .B(n35728), .A(n35729), .Z(n35726) );
  AND U39326 ( .A(a[13]), .B(b[51]), .Z(n35725) );
  XOR U39327 ( .A(n35731), .B(n35732), .Z(n35352) );
  ANDN U39328 ( .B(n35733), .A(n35734), .Z(n35731) );
  AND U39329 ( .A(a[14]), .B(b[50]), .Z(n35730) );
  XOR U39330 ( .A(n35736), .B(n35737), .Z(n35357) );
  ANDN U39331 ( .B(n35738), .A(n35739), .Z(n35736) );
  AND U39332 ( .A(a[15]), .B(b[49]), .Z(n35735) );
  XOR U39333 ( .A(n35741), .B(n35742), .Z(n35362) );
  ANDN U39334 ( .B(n35743), .A(n35744), .Z(n35741) );
  AND U39335 ( .A(a[16]), .B(b[48]), .Z(n35740) );
  XOR U39336 ( .A(n35746), .B(n35747), .Z(n35367) );
  ANDN U39337 ( .B(n35748), .A(n35749), .Z(n35746) );
  AND U39338 ( .A(a[17]), .B(b[47]), .Z(n35745) );
  XOR U39339 ( .A(n35751), .B(n35752), .Z(n35372) );
  ANDN U39340 ( .B(n35753), .A(n35754), .Z(n35751) );
  AND U39341 ( .A(a[18]), .B(b[46]), .Z(n35750) );
  XOR U39342 ( .A(n35756), .B(n35757), .Z(n35377) );
  ANDN U39343 ( .B(n35758), .A(n35759), .Z(n35756) );
  AND U39344 ( .A(a[19]), .B(b[45]), .Z(n35755) );
  XOR U39345 ( .A(n35761), .B(n35762), .Z(n35382) );
  ANDN U39346 ( .B(n35763), .A(n35764), .Z(n35761) );
  AND U39347 ( .A(a[20]), .B(b[44]), .Z(n35760) );
  XOR U39348 ( .A(n35766), .B(n35767), .Z(n35387) );
  ANDN U39349 ( .B(n35768), .A(n35769), .Z(n35766) );
  AND U39350 ( .A(a[21]), .B(b[43]), .Z(n35765) );
  XOR U39351 ( .A(n35771), .B(n35772), .Z(n35392) );
  ANDN U39352 ( .B(n35773), .A(n35774), .Z(n35771) );
  AND U39353 ( .A(a[22]), .B(b[42]), .Z(n35770) );
  XOR U39354 ( .A(n35776), .B(n35777), .Z(n35397) );
  ANDN U39355 ( .B(n35778), .A(n35779), .Z(n35776) );
  AND U39356 ( .A(a[23]), .B(b[41]), .Z(n35775) );
  XOR U39357 ( .A(n35781), .B(n35782), .Z(n35402) );
  ANDN U39358 ( .B(n35783), .A(n35784), .Z(n35781) );
  AND U39359 ( .A(a[24]), .B(b[40]), .Z(n35780) );
  XOR U39360 ( .A(n35786), .B(n35787), .Z(n35407) );
  ANDN U39361 ( .B(n35788), .A(n35789), .Z(n35786) );
  AND U39362 ( .A(a[25]), .B(b[39]), .Z(n35785) );
  XOR U39363 ( .A(n35791), .B(n35792), .Z(n35412) );
  ANDN U39364 ( .B(n35793), .A(n35794), .Z(n35791) );
  AND U39365 ( .A(a[26]), .B(b[38]), .Z(n35790) );
  XOR U39366 ( .A(n35796), .B(n35797), .Z(n35417) );
  ANDN U39367 ( .B(n35798), .A(n35799), .Z(n35796) );
  AND U39368 ( .A(a[27]), .B(b[37]), .Z(n35795) );
  XOR U39369 ( .A(n35801), .B(n35802), .Z(n35422) );
  ANDN U39370 ( .B(n35803), .A(n35804), .Z(n35801) );
  AND U39371 ( .A(a[28]), .B(b[36]), .Z(n35800) );
  XOR U39372 ( .A(n35806), .B(n35807), .Z(n35427) );
  ANDN U39373 ( .B(n35808), .A(n35809), .Z(n35806) );
  AND U39374 ( .A(a[29]), .B(b[35]), .Z(n35805) );
  XOR U39375 ( .A(n35811), .B(n35812), .Z(n35432) );
  ANDN U39376 ( .B(n35813), .A(n35814), .Z(n35811) );
  AND U39377 ( .A(a[30]), .B(b[34]), .Z(n35810) );
  XOR U39378 ( .A(n35816), .B(n35817), .Z(n35437) );
  ANDN U39379 ( .B(n35818), .A(n35819), .Z(n35816) );
  AND U39380 ( .A(a[31]), .B(b[33]), .Z(n35815) );
  XOR U39381 ( .A(n35821), .B(n35822), .Z(n35442) );
  ANDN U39382 ( .B(n35823), .A(n35824), .Z(n35821) );
  AND U39383 ( .A(a[32]), .B(b[32]), .Z(n35820) );
  XOR U39384 ( .A(n35826), .B(n35827), .Z(n35447) );
  ANDN U39385 ( .B(n35828), .A(n35829), .Z(n35826) );
  AND U39386 ( .A(a[33]), .B(b[31]), .Z(n35825) );
  XOR U39387 ( .A(n35831), .B(n35832), .Z(n35452) );
  ANDN U39388 ( .B(n35833), .A(n35834), .Z(n35831) );
  AND U39389 ( .A(a[34]), .B(b[30]), .Z(n35830) );
  XOR U39390 ( .A(n35836), .B(n35837), .Z(n35457) );
  ANDN U39391 ( .B(n35838), .A(n35839), .Z(n35836) );
  AND U39392 ( .A(a[35]), .B(b[29]), .Z(n35835) );
  XOR U39393 ( .A(n35841), .B(n35842), .Z(n35462) );
  ANDN U39394 ( .B(n35843), .A(n35844), .Z(n35841) );
  AND U39395 ( .A(a[36]), .B(b[28]), .Z(n35840) );
  XOR U39396 ( .A(n35846), .B(n35847), .Z(n35467) );
  ANDN U39397 ( .B(n35848), .A(n35849), .Z(n35846) );
  AND U39398 ( .A(a[37]), .B(b[27]), .Z(n35845) );
  XOR U39399 ( .A(n35851), .B(n35852), .Z(n35472) );
  ANDN U39400 ( .B(n35853), .A(n35854), .Z(n35851) );
  AND U39401 ( .A(a[38]), .B(b[26]), .Z(n35850) );
  XOR U39402 ( .A(n35856), .B(n35857), .Z(n35477) );
  ANDN U39403 ( .B(n35858), .A(n35859), .Z(n35856) );
  AND U39404 ( .A(a[39]), .B(b[25]), .Z(n35855) );
  XOR U39405 ( .A(n35861), .B(n35862), .Z(n35482) );
  ANDN U39406 ( .B(n35863), .A(n35864), .Z(n35861) );
  AND U39407 ( .A(a[40]), .B(b[24]), .Z(n35860) );
  XOR U39408 ( .A(n35866), .B(n35867), .Z(n35487) );
  ANDN U39409 ( .B(n35868), .A(n35869), .Z(n35866) );
  AND U39410 ( .A(a[41]), .B(b[23]), .Z(n35865) );
  XOR U39411 ( .A(n35871), .B(n35872), .Z(n35492) );
  ANDN U39412 ( .B(n35873), .A(n35874), .Z(n35871) );
  AND U39413 ( .A(a[42]), .B(b[22]), .Z(n35870) );
  XOR U39414 ( .A(n35876), .B(n35877), .Z(n35497) );
  ANDN U39415 ( .B(n35878), .A(n35879), .Z(n35876) );
  AND U39416 ( .A(a[43]), .B(b[21]), .Z(n35875) );
  XOR U39417 ( .A(n35881), .B(n35882), .Z(n35502) );
  ANDN U39418 ( .B(n35883), .A(n35884), .Z(n35881) );
  AND U39419 ( .A(a[44]), .B(b[20]), .Z(n35880) );
  XOR U39420 ( .A(n35886), .B(n35887), .Z(n35507) );
  ANDN U39421 ( .B(n35888), .A(n35889), .Z(n35886) );
  AND U39422 ( .A(a[45]), .B(b[19]), .Z(n35885) );
  XOR U39423 ( .A(n35891), .B(n35892), .Z(n35512) );
  ANDN U39424 ( .B(n35893), .A(n35894), .Z(n35891) );
  AND U39425 ( .A(a[46]), .B(b[18]), .Z(n35890) );
  XOR U39426 ( .A(n35896), .B(n35897), .Z(n35517) );
  ANDN U39427 ( .B(n35898), .A(n35899), .Z(n35896) );
  AND U39428 ( .A(a[47]), .B(b[17]), .Z(n35895) );
  XOR U39429 ( .A(n35901), .B(n35902), .Z(n35522) );
  ANDN U39430 ( .B(n35903), .A(n35904), .Z(n35901) );
  AND U39431 ( .A(a[48]), .B(b[16]), .Z(n35900) );
  XOR U39432 ( .A(n35906), .B(n35907), .Z(n35527) );
  ANDN U39433 ( .B(n35908), .A(n35909), .Z(n35906) );
  AND U39434 ( .A(a[49]), .B(b[15]), .Z(n35905) );
  XOR U39435 ( .A(n35911), .B(n35912), .Z(n35532) );
  ANDN U39436 ( .B(n35913), .A(n35914), .Z(n35911) );
  AND U39437 ( .A(a[50]), .B(b[14]), .Z(n35910) );
  XOR U39438 ( .A(n35916), .B(n35917), .Z(n35537) );
  ANDN U39439 ( .B(n35918), .A(n35919), .Z(n35916) );
  AND U39440 ( .A(a[51]), .B(b[13]), .Z(n35915) );
  XOR U39441 ( .A(n35921), .B(n35922), .Z(n35542) );
  ANDN U39442 ( .B(n35923), .A(n35924), .Z(n35921) );
  AND U39443 ( .A(a[52]), .B(b[12]), .Z(n35920) );
  XOR U39444 ( .A(n35926), .B(n35927), .Z(n35547) );
  ANDN U39445 ( .B(n35928), .A(n35929), .Z(n35926) );
  AND U39446 ( .A(a[53]), .B(b[11]), .Z(n35925) );
  XOR U39447 ( .A(n35931), .B(n35932), .Z(n35552) );
  ANDN U39448 ( .B(n35933), .A(n35934), .Z(n35931) );
  AND U39449 ( .A(a[54]), .B(b[10]), .Z(n35930) );
  XOR U39450 ( .A(n35936), .B(n35937), .Z(n35557) );
  ANDN U39451 ( .B(n35938), .A(n35939), .Z(n35936) );
  AND U39452 ( .A(b[9]), .B(a[55]), .Z(n35935) );
  XOR U39453 ( .A(n35941), .B(n35942), .Z(n35562) );
  ANDN U39454 ( .B(n35943), .A(n35944), .Z(n35941) );
  AND U39455 ( .A(b[8]), .B(a[56]), .Z(n35940) );
  XOR U39456 ( .A(n35946), .B(n35947), .Z(n35567) );
  ANDN U39457 ( .B(n35948), .A(n35949), .Z(n35946) );
  AND U39458 ( .A(b[7]), .B(a[57]), .Z(n35945) );
  XOR U39459 ( .A(n35951), .B(n35952), .Z(n35572) );
  ANDN U39460 ( .B(n35953), .A(n35954), .Z(n35951) );
  AND U39461 ( .A(b[6]), .B(a[58]), .Z(n35950) );
  XOR U39462 ( .A(n35956), .B(n35957), .Z(n35577) );
  ANDN U39463 ( .B(n35958), .A(n35959), .Z(n35956) );
  AND U39464 ( .A(b[5]), .B(a[59]), .Z(n35955) );
  XOR U39465 ( .A(n35961), .B(n35962), .Z(n35582) );
  ANDN U39466 ( .B(n35963), .A(n35964), .Z(n35961) );
  AND U39467 ( .A(b[4]), .B(a[60]), .Z(n35960) );
  XOR U39468 ( .A(n35966), .B(n35967), .Z(n35587) );
  ANDN U39469 ( .B(n35599), .A(n35600), .Z(n35966) );
  AND U39470 ( .A(b[2]), .B(a[61]), .Z(n35968) );
  XNOR U39471 ( .A(n35963), .B(n35967), .Z(n35969) );
  XOR U39472 ( .A(n35970), .B(n35971), .Z(n35967) );
  OR U39473 ( .A(n35602), .B(n35603), .Z(n35971) );
  XNOR U39474 ( .A(n35973), .B(n35974), .Z(n35972) );
  XOR U39475 ( .A(n35973), .B(n35976), .Z(n35602) );
  NAND U39476 ( .A(b[1]), .B(a[61]), .Z(n35976) );
  IV U39477 ( .A(n35970), .Z(n35973) );
  NANDN U39478 ( .A(n85), .B(n86), .Z(n35970) );
  XOR U39479 ( .A(n35977), .B(n35978), .Z(n86) );
  NAND U39480 ( .A(a[61]), .B(b[0]), .Z(n85) );
  XNOR U39481 ( .A(n35958), .B(n35962), .Z(n35979) );
  XNOR U39482 ( .A(n35953), .B(n35957), .Z(n35980) );
  XNOR U39483 ( .A(n35948), .B(n35952), .Z(n35981) );
  XNOR U39484 ( .A(n35943), .B(n35947), .Z(n35982) );
  XNOR U39485 ( .A(n35938), .B(n35942), .Z(n35983) );
  XNOR U39486 ( .A(n35933), .B(n35937), .Z(n35984) );
  XNOR U39487 ( .A(n35928), .B(n35932), .Z(n35985) );
  XNOR U39488 ( .A(n35923), .B(n35927), .Z(n35986) );
  XNOR U39489 ( .A(n35918), .B(n35922), .Z(n35987) );
  XNOR U39490 ( .A(n35913), .B(n35917), .Z(n35988) );
  XNOR U39491 ( .A(n35908), .B(n35912), .Z(n35989) );
  XNOR U39492 ( .A(n35903), .B(n35907), .Z(n35990) );
  XNOR U39493 ( .A(n35898), .B(n35902), .Z(n35991) );
  XNOR U39494 ( .A(n35893), .B(n35897), .Z(n35992) );
  XNOR U39495 ( .A(n35888), .B(n35892), .Z(n35993) );
  XNOR U39496 ( .A(n35883), .B(n35887), .Z(n35994) );
  XNOR U39497 ( .A(n35878), .B(n35882), .Z(n35995) );
  XNOR U39498 ( .A(n35873), .B(n35877), .Z(n35996) );
  XNOR U39499 ( .A(n35868), .B(n35872), .Z(n35997) );
  XNOR U39500 ( .A(n35863), .B(n35867), .Z(n35998) );
  XNOR U39501 ( .A(n35858), .B(n35862), .Z(n35999) );
  XNOR U39502 ( .A(n35853), .B(n35857), .Z(n36000) );
  XNOR U39503 ( .A(n35848), .B(n35852), .Z(n36001) );
  XNOR U39504 ( .A(n35843), .B(n35847), .Z(n36002) );
  XNOR U39505 ( .A(n35838), .B(n35842), .Z(n36003) );
  XNOR U39506 ( .A(n35833), .B(n35837), .Z(n36004) );
  XNOR U39507 ( .A(n35828), .B(n35832), .Z(n36005) );
  XNOR U39508 ( .A(n35823), .B(n35827), .Z(n36006) );
  XNOR U39509 ( .A(n35818), .B(n35822), .Z(n36007) );
  XNOR U39510 ( .A(n35813), .B(n35817), .Z(n36008) );
  XNOR U39511 ( .A(n35808), .B(n35812), .Z(n36009) );
  XNOR U39512 ( .A(n35803), .B(n35807), .Z(n36010) );
  XNOR U39513 ( .A(n35798), .B(n35802), .Z(n36011) );
  XNOR U39514 ( .A(n35793), .B(n35797), .Z(n36012) );
  XNOR U39515 ( .A(n35788), .B(n35792), .Z(n36013) );
  XNOR U39516 ( .A(n35783), .B(n35787), .Z(n36014) );
  XNOR U39517 ( .A(n35778), .B(n35782), .Z(n36015) );
  XNOR U39518 ( .A(n35773), .B(n35777), .Z(n36016) );
  XNOR U39519 ( .A(n35768), .B(n35772), .Z(n36017) );
  XNOR U39520 ( .A(n35763), .B(n35767), .Z(n36018) );
  XNOR U39521 ( .A(n35758), .B(n35762), .Z(n36019) );
  XNOR U39522 ( .A(n35753), .B(n35757), .Z(n36020) );
  XNOR U39523 ( .A(n35748), .B(n35752), .Z(n36021) );
  XNOR U39524 ( .A(n35743), .B(n35747), .Z(n36022) );
  XNOR U39525 ( .A(n35738), .B(n35742), .Z(n36023) );
  XNOR U39526 ( .A(n35733), .B(n35737), .Z(n36024) );
  XNOR U39527 ( .A(n35728), .B(n35732), .Z(n36025) );
  XNOR U39528 ( .A(n35723), .B(n35727), .Z(n36026) );
  XNOR U39529 ( .A(n35718), .B(n35722), .Z(n36027) );
  XNOR U39530 ( .A(n35713), .B(n35717), .Z(n36028) );
  XNOR U39531 ( .A(n35708), .B(n35712), .Z(n36029) );
  XNOR U39532 ( .A(n35703), .B(n35707), .Z(n36030) );
  XNOR U39533 ( .A(n35698), .B(n35702), .Z(n36031) );
  XNOR U39534 ( .A(n35693), .B(n35697), .Z(n36032) );
  XNOR U39535 ( .A(n35688), .B(n35692), .Z(n36033) );
  XNOR U39536 ( .A(n35683), .B(n35687), .Z(n36034) );
  XNOR U39537 ( .A(n35678), .B(n35682), .Z(n36035) );
  XNOR U39538 ( .A(n35673), .B(n35677), .Z(n36036) );
  XNOR U39539 ( .A(n35668), .B(n35672), .Z(n36037) );
  XNOR U39540 ( .A(n36038), .B(n35667), .Z(n35668) );
  AND U39541 ( .A(a[0]), .B(b[63]), .Z(n36038) );
  XOR U39542 ( .A(n36039), .B(n35667), .Z(n35669) );
  XNOR U39543 ( .A(n36040), .B(n36041), .Z(n35667) );
  ANDN U39544 ( .B(n36042), .A(n36043), .Z(n36040) );
  AND U39545 ( .A(a[1]), .B(b[62]), .Z(n36039) );
  XOR U39546 ( .A(n36045), .B(n36046), .Z(n35672) );
  ANDN U39547 ( .B(n36047), .A(n36048), .Z(n36045) );
  AND U39548 ( .A(a[2]), .B(b[61]), .Z(n36044) );
  XOR U39549 ( .A(n36050), .B(n36051), .Z(n35677) );
  ANDN U39550 ( .B(n36052), .A(n36053), .Z(n36050) );
  AND U39551 ( .A(a[3]), .B(b[60]), .Z(n36049) );
  XOR U39552 ( .A(n36055), .B(n36056), .Z(n35682) );
  ANDN U39553 ( .B(n36057), .A(n36058), .Z(n36055) );
  AND U39554 ( .A(a[4]), .B(b[59]), .Z(n36054) );
  XOR U39555 ( .A(n36060), .B(n36061), .Z(n35687) );
  ANDN U39556 ( .B(n36062), .A(n36063), .Z(n36060) );
  AND U39557 ( .A(a[5]), .B(b[58]), .Z(n36059) );
  XOR U39558 ( .A(n36065), .B(n36066), .Z(n35692) );
  ANDN U39559 ( .B(n36067), .A(n36068), .Z(n36065) );
  AND U39560 ( .A(a[6]), .B(b[57]), .Z(n36064) );
  XOR U39561 ( .A(n36070), .B(n36071), .Z(n35697) );
  ANDN U39562 ( .B(n36072), .A(n36073), .Z(n36070) );
  AND U39563 ( .A(a[7]), .B(b[56]), .Z(n36069) );
  XOR U39564 ( .A(n36075), .B(n36076), .Z(n35702) );
  ANDN U39565 ( .B(n36077), .A(n36078), .Z(n36075) );
  AND U39566 ( .A(a[8]), .B(b[55]), .Z(n36074) );
  XOR U39567 ( .A(n36080), .B(n36081), .Z(n35707) );
  ANDN U39568 ( .B(n36082), .A(n36083), .Z(n36080) );
  AND U39569 ( .A(a[9]), .B(b[54]), .Z(n36079) );
  XOR U39570 ( .A(n36085), .B(n36086), .Z(n35712) );
  ANDN U39571 ( .B(n36087), .A(n36088), .Z(n36085) );
  AND U39572 ( .A(a[10]), .B(b[53]), .Z(n36084) );
  XOR U39573 ( .A(n36090), .B(n36091), .Z(n35717) );
  ANDN U39574 ( .B(n36092), .A(n36093), .Z(n36090) );
  AND U39575 ( .A(a[11]), .B(b[52]), .Z(n36089) );
  XOR U39576 ( .A(n36095), .B(n36096), .Z(n35722) );
  ANDN U39577 ( .B(n36097), .A(n36098), .Z(n36095) );
  AND U39578 ( .A(a[12]), .B(b[51]), .Z(n36094) );
  XOR U39579 ( .A(n36100), .B(n36101), .Z(n35727) );
  ANDN U39580 ( .B(n36102), .A(n36103), .Z(n36100) );
  AND U39581 ( .A(a[13]), .B(b[50]), .Z(n36099) );
  XOR U39582 ( .A(n36105), .B(n36106), .Z(n35732) );
  ANDN U39583 ( .B(n36107), .A(n36108), .Z(n36105) );
  AND U39584 ( .A(a[14]), .B(b[49]), .Z(n36104) );
  XOR U39585 ( .A(n36110), .B(n36111), .Z(n35737) );
  ANDN U39586 ( .B(n36112), .A(n36113), .Z(n36110) );
  AND U39587 ( .A(a[15]), .B(b[48]), .Z(n36109) );
  XOR U39588 ( .A(n36115), .B(n36116), .Z(n35742) );
  ANDN U39589 ( .B(n36117), .A(n36118), .Z(n36115) );
  AND U39590 ( .A(a[16]), .B(b[47]), .Z(n36114) );
  XOR U39591 ( .A(n36120), .B(n36121), .Z(n35747) );
  ANDN U39592 ( .B(n36122), .A(n36123), .Z(n36120) );
  AND U39593 ( .A(a[17]), .B(b[46]), .Z(n36119) );
  XOR U39594 ( .A(n36125), .B(n36126), .Z(n35752) );
  ANDN U39595 ( .B(n36127), .A(n36128), .Z(n36125) );
  AND U39596 ( .A(a[18]), .B(b[45]), .Z(n36124) );
  XOR U39597 ( .A(n36130), .B(n36131), .Z(n35757) );
  ANDN U39598 ( .B(n36132), .A(n36133), .Z(n36130) );
  AND U39599 ( .A(a[19]), .B(b[44]), .Z(n36129) );
  XOR U39600 ( .A(n36135), .B(n36136), .Z(n35762) );
  ANDN U39601 ( .B(n36137), .A(n36138), .Z(n36135) );
  AND U39602 ( .A(a[20]), .B(b[43]), .Z(n36134) );
  XOR U39603 ( .A(n36140), .B(n36141), .Z(n35767) );
  ANDN U39604 ( .B(n36142), .A(n36143), .Z(n36140) );
  AND U39605 ( .A(a[21]), .B(b[42]), .Z(n36139) );
  XOR U39606 ( .A(n36145), .B(n36146), .Z(n35772) );
  ANDN U39607 ( .B(n36147), .A(n36148), .Z(n36145) );
  AND U39608 ( .A(a[22]), .B(b[41]), .Z(n36144) );
  XOR U39609 ( .A(n36150), .B(n36151), .Z(n35777) );
  ANDN U39610 ( .B(n36152), .A(n36153), .Z(n36150) );
  AND U39611 ( .A(a[23]), .B(b[40]), .Z(n36149) );
  XOR U39612 ( .A(n36155), .B(n36156), .Z(n35782) );
  ANDN U39613 ( .B(n36157), .A(n36158), .Z(n36155) );
  AND U39614 ( .A(a[24]), .B(b[39]), .Z(n36154) );
  XOR U39615 ( .A(n36160), .B(n36161), .Z(n35787) );
  ANDN U39616 ( .B(n36162), .A(n36163), .Z(n36160) );
  AND U39617 ( .A(a[25]), .B(b[38]), .Z(n36159) );
  XOR U39618 ( .A(n36165), .B(n36166), .Z(n35792) );
  ANDN U39619 ( .B(n36167), .A(n36168), .Z(n36165) );
  AND U39620 ( .A(a[26]), .B(b[37]), .Z(n36164) );
  XOR U39621 ( .A(n36170), .B(n36171), .Z(n35797) );
  ANDN U39622 ( .B(n36172), .A(n36173), .Z(n36170) );
  AND U39623 ( .A(a[27]), .B(b[36]), .Z(n36169) );
  XOR U39624 ( .A(n36175), .B(n36176), .Z(n35802) );
  ANDN U39625 ( .B(n36177), .A(n36178), .Z(n36175) );
  AND U39626 ( .A(a[28]), .B(b[35]), .Z(n36174) );
  XOR U39627 ( .A(n36180), .B(n36181), .Z(n35807) );
  ANDN U39628 ( .B(n36182), .A(n36183), .Z(n36180) );
  AND U39629 ( .A(a[29]), .B(b[34]), .Z(n36179) );
  XOR U39630 ( .A(n36185), .B(n36186), .Z(n35812) );
  ANDN U39631 ( .B(n36187), .A(n36188), .Z(n36185) );
  AND U39632 ( .A(a[30]), .B(b[33]), .Z(n36184) );
  XOR U39633 ( .A(n36190), .B(n36191), .Z(n35817) );
  ANDN U39634 ( .B(n36192), .A(n36193), .Z(n36190) );
  AND U39635 ( .A(a[31]), .B(b[32]), .Z(n36189) );
  XOR U39636 ( .A(n36195), .B(n36196), .Z(n35822) );
  ANDN U39637 ( .B(n36197), .A(n36198), .Z(n36195) );
  AND U39638 ( .A(a[32]), .B(b[31]), .Z(n36194) );
  XOR U39639 ( .A(n36200), .B(n36201), .Z(n35827) );
  ANDN U39640 ( .B(n36202), .A(n36203), .Z(n36200) );
  AND U39641 ( .A(a[33]), .B(b[30]), .Z(n36199) );
  XOR U39642 ( .A(n36205), .B(n36206), .Z(n35832) );
  ANDN U39643 ( .B(n36207), .A(n36208), .Z(n36205) );
  AND U39644 ( .A(a[34]), .B(b[29]), .Z(n36204) );
  XOR U39645 ( .A(n36210), .B(n36211), .Z(n35837) );
  ANDN U39646 ( .B(n36212), .A(n36213), .Z(n36210) );
  AND U39647 ( .A(a[35]), .B(b[28]), .Z(n36209) );
  XOR U39648 ( .A(n36215), .B(n36216), .Z(n35842) );
  ANDN U39649 ( .B(n36217), .A(n36218), .Z(n36215) );
  AND U39650 ( .A(a[36]), .B(b[27]), .Z(n36214) );
  XOR U39651 ( .A(n36220), .B(n36221), .Z(n35847) );
  ANDN U39652 ( .B(n36222), .A(n36223), .Z(n36220) );
  AND U39653 ( .A(a[37]), .B(b[26]), .Z(n36219) );
  XOR U39654 ( .A(n36225), .B(n36226), .Z(n35852) );
  ANDN U39655 ( .B(n36227), .A(n36228), .Z(n36225) );
  AND U39656 ( .A(a[38]), .B(b[25]), .Z(n36224) );
  XOR U39657 ( .A(n36230), .B(n36231), .Z(n35857) );
  ANDN U39658 ( .B(n36232), .A(n36233), .Z(n36230) );
  AND U39659 ( .A(a[39]), .B(b[24]), .Z(n36229) );
  XOR U39660 ( .A(n36235), .B(n36236), .Z(n35862) );
  ANDN U39661 ( .B(n36237), .A(n36238), .Z(n36235) );
  AND U39662 ( .A(a[40]), .B(b[23]), .Z(n36234) );
  XOR U39663 ( .A(n36240), .B(n36241), .Z(n35867) );
  ANDN U39664 ( .B(n36242), .A(n36243), .Z(n36240) );
  AND U39665 ( .A(a[41]), .B(b[22]), .Z(n36239) );
  XOR U39666 ( .A(n36245), .B(n36246), .Z(n35872) );
  ANDN U39667 ( .B(n36247), .A(n36248), .Z(n36245) );
  AND U39668 ( .A(a[42]), .B(b[21]), .Z(n36244) );
  XOR U39669 ( .A(n36250), .B(n36251), .Z(n35877) );
  ANDN U39670 ( .B(n36252), .A(n36253), .Z(n36250) );
  AND U39671 ( .A(a[43]), .B(b[20]), .Z(n36249) );
  XOR U39672 ( .A(n36255), .B(n36256), .Z(n35882) );
  ANDN U39673 ( .B(n36257), .A(n36258), .Z(n36255) );
  AND U39674 ( .A(a[44]), .B(b[19]), .Z(n36254) );
  XOR U39675 ( .A(n36260), .B(n36261), .Z(n35887) );
  ANDN U39676 ( .B(n36262), .A(n36263), .Z(n36260) );
  AND U39677 ( .A(a[45]), .B(b[18]), .Z(n36259) );
  XOR U39678 ( .A(n36265), .B(n36266), .Z(n35892) );
  ANDN U39679 ( .B(n36267), .A(n36268), .Z(n36265) );
  AND U39680 ( .A(a[46]), .B(b[17]), .Z(n36264) );
  XOR U39681 ( .A(n36270), .B(n36271), .Z(n35897) );
  ANDN U39682 ( .B(n36272), .A(n36273), .Z(n36270) );
  AND U39683 ( .A(a[47]), .B(b[16]), .Z(n36269) );
  XOR U39684 ( .A(n36275), .B(n36276), .Z(n35902) );
  ANDN U39685 ( .B(n36277), .A(n36278), .Z(n36275) );
  AND U39686 ( .A(a[48]), .B(b[15]), .Z(n36274) );
  XOR U39687 ( .A(n36280), .B(n36281), .Z(n35907) );
  ANDN U39688 ( .B(n36282), .A(n36283), .Z(n36280) );
  AND U39689 ( .A(a[49]), .B(b[14]), .Z(n36279) );
  XOR U39690 ( .A(n36285), .B(n36286), .Z(n35912) );
  ANDN U39691 ( .B(n36287), .A(n36288), .Z(n36285) );
  AND U39692 ( .A(a[50]), .B(b[13]), .Z(n36284) );
  XOR U39693 ( .A(n36290), .B(n36291), .Z(n35917) );
  ANDN U39694 ( .B(n36292), .A(n36293), .Z(n36290) );
  AND U39695 ( .A(a[51]), .B(b[12]), .Z(n36289) );
  XOR U39696 ( .A(n36295), .B(n36296), .Z(n35922) );
  ANDN U39697 ( .B(n36297), .A(n36298), .Z(n36295) );
  AND U39698 ( .A(a[52]), .B(b[11]), .Z(n36294) );
  XOR U39699 ( .A(n36300), .B(n36301), .Z(n35927) );
  ANDN U39700 ( .B(n36302), .A(n36303), .Z(n36300) );
  AND U39701 ( .A(a[53]), .B(b[10]), .Z(n36299) );
  XOR U39702 ( .A(n36305), .B(n36306), .Z(n35932) );
  ANDN U39703 ( .B(n36307), .A(n36308), .Z(n36305) );
  AND U39704 ( .A(b[9]), .B(a[54]), .Z(n36304) );
  XOR U39705 ( .A(n36310), .B(n36311), .Z(n35937) );
  ANDN U39706 ( .B(n36312), .A(n36313), .Z(n36310) );
  AND U39707 ( .A(b[8]), .B(a[55]), .Z(n36309) );
  XOR U39708 ( .A(n36315), .B(n36316), .Z(n35942) );
  ANDN U39709 ( .B(n36317), .A(n36318), .Z(n36315) );
  AND U39710 ( .A(b[7]), .B(a[56]), .Z(n36314) );
  XOR U39711 ( .A(n36320), .B(n36321), .Z(n35947) );
  ANDN U39712 ( .B(n36322), .A(n36323), .Z(n36320) );
  AND U39713 ( .A(b[6]), .B(a[57]), .Z(n36319) );
  XOR U39714 ( .A(n36325), .B(n36326), .Z(n35952) );
  ANDN U39715 ( .B(n36327), .A(n36328), .Z(n36325) );
  AND U39716 ( .A(b[5]), .B(a[58]), .Z(n36324) );
  XOR U39717 ( .A(n36330), .B(n36331), .Z(n35957) );
  ANDN U39718 ( .B(n36332), .A(n36333), .Z(n36330) );
  AND U39719 ( .A(b[4]), .B(a[59]), .Z(n36329) );
  XOR U39720 ( .A(n36335), .B(n36336), .Z(n35962) );
  ANDN U39721 ( .B(n35974), .A(n35975), .Z(n36335) );
  AND U39722 ( .A(b[2]), .B(a[60]), .Z(n36337) );
  XNOR U39723 ( .A(n36332), .B(n36336), .Z(n36338) );
  XOR U39724 ( .A(n36339), .B(n36340), .Z(n36336) );
  OR U39725 ( .A(n35977), .B(n35978), .Z(n36340) );
  XNOR U39726 ( .A(n36342), .B(n36343), .Z(n36341) );
  XOR U39727 ( .A(n36342), .B(n36345), .Z(n35977) );
  NAND U39728 ( .A(b[1]), .B(a[60]), .Z(n36345) );
  IV U39729 ( .A(n36339), .Z(n36342) );
  NANDN U39730 ( .A(n87), .B(n88), .Z(n36339) );
  XOR U39731 ( .A(n36346), .B(n36347), .Z(n88) );
  NAND U39732 ( .A(a[60]), .B(b[0]), .Z(n87) );
  XNOR U39733 ( .A(n36327), .B(n36331), .Z(n36348) );
  XNOR U39734 ( .A(n36322), .B(n36326), .Z(n36349) );
  XNOR U39735 ( .A(n36317), .B(n36321), .Z(n36350) );
  XNOR U39736 ( .A(n36312), .B(n36316), .Z(n36351) );
  XNOR U39737 ( .A(n36307), .B(n36311), .Z(n36352) );
  XNOR U39738 ( .A(n36302), .B(n36306), .Z(n36353) );
  XNOR U39739 ( .A(n36297), .B(n36301), .Z(n36354) );
  XNOR U39740 ( .A(n36292), .B(n36296), .Z(n36355) );
  XNOR U39741 ( .A(n36287), .B(n36291), .Z(n36356) );
  XNOR U39742 ( .A(n36282), .B(n36286), .Z(n36357) );
  XNOR U39743 ( .A(n36277), .B(n36281), .Z(n36358) );
  XNOR U39744 ( .A(n36272), .B(n36276), .Z(n36359) );
  XNOR U39745 ( .A(n36267), .B(n36271), .Z(n36360) );
  XNOR U39746 ( .A(n36262), .B(n36266), .Z(n36361) );
  XNOR U39747 ( .A(n36257), .B(n36261), .Z(n36362) );
  XNOR U39748 ( .A(n36252), .B(n36256), .Z(n36363) );
  XNOR U39749 ( .A(n36247), .B(n36251), .Z(n36364) );
  XNOR U39750 ( .A(n36242), .B(n36246), .Z(n36365) );
  XNOR U39751 ( .A(n36237), .B(n36241), .Z(n36366) );
  XNOR U39752 ( .A(n36232), .B(n36236), .Z(n36367) );
  XNOR U39753 ( .A(n36227), .B(n36231), .Z(n36368) );
  XNOR U39754 ( .A(n36222), .B(n36226), .Z(n36369) );
  XNOR U39755 ( .A(n36217), .B(n36221), .Z(n36370) );
  XNOR U39756 ( .A(n36212), .B(n36216), .Z(n36371) );
  XNOR U39757 ( .A(n36207), .B(n36211), .Z(n36372) );
  XNOR U39758 ( .A(n36202), .B(n36206), .Z(n36373) );
  XNOR U39759 ( .A(n36197), .B(n36201), .Z(n36374) );
  XNOR U39760 ( .A(n36192), .B(n36196), .Z(n36375) );
  XNOR U39761 ( .A(n36187), .B(n36191), .Z(n36376) );
  XNOR U39762 ( .A(n36182), .B(n36186), .Z(n36377) );
  XNOR U39763 ( .A(n36177), .B(n36181), .Z(n36378) );
  XNOR U39764 ( .A(n36172), .B(n36176), .Z(n36379) );
  XNOR U39765 ( .A(n36167), .B(n36171), .Z(n36380) );
  XNOR U39766 ( .A(n36162), .B(n36166), .Z(n36381) );
  XNOR U39767 ( .A(n36157), .B(n36161), .Z(n36382) );
  XNOR U39768 ( .A(n36152), .B(n36156), .Z(n36383) );
  XNOR U39769 ( .A(n36147), .B(n36151), .Z(n36384) );
  XNOR U39770 ( .A(n36142), .B(n36146), .Z(n36385) );
  XNOR U39771 ( .A(n36137), .B(n36141), .Z(n36386) );
  XNOR U39772 ( .A(n36132), .B(n36136), .Z(n36387) );
  XNOR U39773 ( .A(n36127), .B(n36131), .Z(n36388) );
  XNOR U39774 ( .A(n36122), .B(n36126), .Z(n36389) );
  XNOR U39775 ( .A(n36117), .B(n36121), .Z(n36390) );
  XNOR U39776 ( .A(n36112), .B(n36116), .Z(n36391) );
  XNOR U39777 ( .A(n36107), .B(n36111), .Z(n36392) );
  XNOR U39778 ( .A(n36102), .B(n36106), .Z(n36393) );
  XNOR U39779 ( .A(n36097), .B(n36101), .Z(n36394) );
  XNOR U39780 ( .A(n36092), .B(n36096), .Z(n36395) );
  XNOR U39781 ( .A(n36087), .B(n36091), .Z(n36396) );
  XNOR U39782 ( .A(n36082), .B(n36086), .Z(n36397) );
  XNOR U39783 ( .A(n36077), .B(n36081), .Z(n36398) );
  XNOR U39784 ( .A(n36072), .B(n36076), .Z(n36399) );
  XNOR U39785 ( .A(n36067), .B(n36071), .Z(n36400) );
  XNOR U39786 ( .A(n36062), .B(n36066), .Z(n36401) );
  XNOR U39787 ( .A(n36057), .B(n36061), .Z(n36402) );
  XNOR U39788 ( .A(n36052), .B(n36056), .Z(n36403) );
  XNOR U39789 ( .A(n36047), .B(n36051), .Z(n36404) );
  XNOR U39790 ( .A(n36042), .B(n36046), .Z(n36405) );
  XOR U39791 ( .A(n36406), .B(n36041), .Z(n36042) );
  AND U39792 ( .A(a[0]), .B(b[62]), .Z(n36406) );
  XNOR U39793 ( .A(n36407), .B(n36041), .Z(n36043) );
  XNOR U39794 ( .A(n36408), .B(n36409), .Z(n36041) );
  ANDN U39795 ( .B(n36410), .A(n36411), .Z(n36408) );
  AND U39796 ( .A(a[1]), .B(b[61]), .Z(n36407) );
  XOR U39797 ( .A(n36413), .B(n36414), .Z(n36046) );
  ANDN U39798 ( .B(n36415), .A(n36416), .Z(n36413) );
  AND U39799 ( .A(a[2]), .B(b[60]), .Z(n36412) );
  XOR U39800 ( .A(n36418), .B(n36419), .Z(n36051) );
  ANDN U39801 ( .B(n36420), .A(n36421), .Z(n36418) );
  AND U39802 ( .A(a[3]), .B(b[59]), .Z(n36417) );
  XOR U39803 ( .A(n36423), .B(n36424), .Z(n36056) );
  ANDN U39804 ( .B(n36425), .A(n36426), .Z(n36423) );
  AND U39805 ( .A(a[4]), .B(b[58]), .Z(n36422) );
  XOR U39806 ( .A(n36428), .B(n36429), .Z(n36061) );
  ANDN U39807 ( .B(n36430), .A(n36431), .Z(n36428) );
  AND U39808 ( .A(a[5]), .B(b[57]), .Z(n36427) );
  XOR U39809 ( .A(n36433), .B(n36434), .Z(n36066) );
  ANDN U39810 ( .B(n36435), .A(n36436), .Z(n36433) );
  AND U39811 ( .A(a[6]), .B(b[56]), .Z(n36432) );
  XOR U39812 ( .A(n36438), .B(n36439), .Z(n36071) );
  ANDN U39813 ( .B(n36440), .A(n36441), .Z(n36438) );
  AND U39814 ( .A(a[7]), .B(b[55]), .Z(n36437) );
  XOR U39815 ( .A(n36443), .B(n36444), .Z(n36076) );
  ANDN U39816 ( .B(n36445), .A(n36446), .Z(n36443) );
  AND U39817 ( .A(a[8]), .B(b[54]), .Z(n36442) );
  XOR U39818 ( .A(n36448), .B(n36449), .Z(n36081) );
  ANDN U39819 ( .B(n36450), .A(n36451), .Z(n36448) );
  AND U39820 ( .A(a[9]), .B(b[53]), .Z(n36447) );
  XOR U39821 ( .A(n36453), .B(n36454), .Z(n36086) );
  ANDN U39822 ( .B(n36455), .A(n36456), .Z(n36453) );
  AND U39823 ( .A(a[10]), .B(b[52]), .Z(n36452) );
  XOR U39824 ( .A(n36458), .B(n36459), .Z(n36091) );
  ANDN U39825 ( .B(n36460), .A(n36461), .Z(n36458) );
  AND U39826 ( .A(a[11]), .B(b[51]), .Z(n36457) );
  XOR U39827 ( .A(n36463), .B(n36464), .Z(n36096) );
  ANDN U39828 ( .B(n36465), .A(n36466), .Z(n36463) );
  AND U39829 ( .A(a[12]), .B(b[50]), .Z(n36462) );
  XOR U39830 ( .A(n36468), .B(n36469), .Z(n36101) );
  ANDN U39831 ( .B(n36470), .A(n36471), .Z(n36468) );
  AND U39832 ( .A(a[13]), .B(b[49]), .Z(n36467) );
  XOR U39833 ( .A(n36473), .B(n36474), .Z(n36106) );
  ANDN U39834 ( .B(n36475), .A(n36476), .Z(n36473) );
  AND U39835 ( .A(a[14]), .B(b[48]), .Z(n36472) );
  XOR U39836 ( .A(n36478), .B(n36479), .Z(n36111) );
  ANDN U39837 ( .B(n36480), .A(n36481), .Z(n36478) );
  AND U39838 ( .A(a[15]), .B(b[47]), .Z(n36477) );
  XOR U39839 ( .A(n36483), .B(n36484), .Z(n36116) );
  ANDN U39840 ( .B(n36485), .A(n36486), .Z(n36483) );
  AND U39841 ( .A(a[16]), .B(b[46]), .Z(n36482) );
  XOR U39842 ( .A(n36488), .B(n36489), .Z(n36121) );
  ANDN U39843 ( .B(n36490), .A(n36491), .Z(n36488) );
  AND U39844 ( .A(a[17]), .B(b[45]), .Z(n36487) );
  XOR U39845 ( .A(n36493), .B(n36494), .Z(n36126) );
  ANDN U39846 ( .B(n36495), .A(n36496), .Z(n36493) );
  AND U39847 ( .A(a[18]), .B(b[44]), .Z(n36492) );
  XOR U39848 ( .A(n36498), .B(n36499), .Z(n36131) );
  ANDN U39849 ( .B(n36500), .A(n36501), .Z(n36498) );
  AND U39850 ( .A(a[19]), .B(b[43]), .Z(n36497) );
  XOR U39851 ( .A(n36503), .B(n36504), .Z(n36136) );
  ANDN U39852 ( .B(n36505), .A(n36506), .Z(n36503) );
  AND U39853 ( .A(a[20]), .B(b[42]), .Z(n36502) );
  XOR U39854 ( .A(n36508), .B(n36509), .Z(n36141) );
  ANDN U39855 ( .B(n36510), .A(n36511), .Z(n36508) );
  AND U39856 ( .A(a[21]), .B(b[41]), .Z(n36507) );
  XOR U39857 ( .A(n36513), .B(n36514), .Z(n36146) );
  ANDN U39858 ( .B(n36515), .A(n36516), .Z(n36513) );
  AND U39859 ( .A(a[22]), .B(b[40]), .Z(n36512) );
  XOR U39860 ( .A(n36518), .B(n36519), .Z(n36151) );
  ANDN U39861 ( .B(n36520), .A(n36521), .Z(n36518) );
  AND U39862 ( .A(a[23]), .B(b[39]), .Z(n36517) );
  XOR U39863 ( .A(n36523), .B(n36524), .Z(n36156) );
  ANDN U39864 ( .B(n36525), .A(n36526), .Z(n36523) );
  AND U39865 ( .A(a[24]), .B(b[38]), .Z(n36522) );
  XOR U39866 ( .A(n36528), .B(n36529), .Z(n36161) );
  ANDN U39867 ( .B(n36530), .A(n36531), .Z(n36528) );
  AND U39868 ( .A(a[25]), .B(b[37]), .Z(n36527) );
  XOR U39869 ( .A(n36533), .B(n36534), .Z(n36166) );
  ANDN U39870 ( .B(n36535), .A(n36536), .Z(n36533) );
  AND U39871 ( .A(a[26]), .B(b[36]), .Z(n36532) );
  XOR U39872 ( .A(n36538), .B(n36539), .Z(n36171) );
  ANDN U39873 ( .B(n36540), .A(n36541), .Z(n36538) );
  AND U39874 ( .A(a[27]), .B(b[35]), .Z(n36537) );
  XOR U39875 ( .A(n36543), .B(n36544), .Z(n36176) );
  ANDN U39876 ( .B(n36545), .A(n36546), .Z(n36543) );
  AND U39877 ( .A(a[28]), .B(b[34]), .Z(n36542) );
  XOR U39878 ( .A(n36548), .B(n36549), .Z(n36181) );
  ANDN U39879 ( .B(n36550), .A(n36551), .Z(n36548) );
  AND U39880 ( .A(a[29]), .B(b[33]), .Z(n36547) );
  XOR U39881 ( .A(n36553), .B(n36554), .Z(n36186) );
  ANDN U39882 ( .B(n36555), .A(n36556), .Z(n36553) );
  AND U39883 ( .A(a[30]), .B(b[32]), .Z(n36552) );
  XOR U39884 ( .A(n36558), .B(n36559), .Z(n36191) );
  ANDN U39885 ( .B(n36560), .A(n36561), .Z(n36558) );
  AND U39886 ( .A(a[31]), .B(b[31]), .Z(n36557) );
  XOR U39887 ( .A(n36563), .B(n36564), .Z(n36196) );
  ANDN U39888 ( .B(n36565), .A(n36566), .Z(n36563) );
  AND U39889 ( .A(a[32]), .B(b[30]), .Z(n36562) );
  XOR U39890 ( .A(n36568), .B(n36569), .Z(n36201) );
  ANDN U39891 ( .B(n36570), .A(n36571), .Z(n36568) );
  AND U39892 ( .A(a[33]), .B(b[29]), .Z(n36567) );
  XOR U39893 ( .A(n36573), .B(n36574), .Z(n36206) );
  ANDN U39894 ( .B(n36575), .A(n36576), .Z(n36573) );
  AND U39895 ( .A(a[34]), .B(b[28]), .Z(n36572) );
  XOR U39896 ( .A(n36578), .B(n36579), .Z(n36211) );
  ANDN U39897 ( .B(n36580), .A(n36581), .Z(n36578) );
  AND U39898 ( .A(a[35]), .B(b[27]), .Z(n36577) );
  XOR U39899 ( .A(n36583), .B(n36584), .Z(n36216) );
  ANDN U39900 ( .B(n36585), .A(n36586), .Z(n36583) );
  AND U39901 ( .A(a[36]), .B(b[26]), .Z(n36582) );
  XOR U39902 ( .A(n36588), .B(n36589), .Z(n36221) );
  ANDN U39903 ( .B(n36590), .A(n36591), .Z(n36588) );
  AND U39904 ( .A(a[37]), .B(b[25]), .Z(n36587) );
  XOR U39905 ( .A(n36593), .B(n36594), .Z(n36226) );
  ANDN U39906 ( .B(n36595), .A(n36596), .Z(n36593) );
  AND U39907 ( .A(a[38]), .B(b[24]), .Z(n36592) );
  XOR U39908 ( .A(n36598), .B(n36599), .Z(n36231) );
  ANDN U39909 ( .B(n36600), .A(n36601), .Z(n36598) );
  AND U39910 ( .A(a[39]), .B(b[23]), .Z(n36597) );
  XOR U39911 ( .A(n36603), .B(n36604), .Z(n36236) );
  ANDN U39912 ( .B(n36605), .A(n36606), .Z(n36603) );
  AND U39913 ( .A(a[40]), .B(b[22]), .Z(n36602) );
  XOR U39914 ( .A(n36608), .B(n36609), .Z(n36241) );
  ANDN U39915 ( .B(n36610), .A(n36611), .Z(n36608) );
  AND U39916 ( .A(a[41]), .B(b[21]), .Z(n36607) );
  XOR U39917 ( .A(n36613), .B(n36614), .Z(n36246) );
  ANDN U39918 ( .B(n36615), .A(n36616), .Z(n36613) );
  AND U39919 ( .A(a[42]), .B(b[20]), .Z(n36612) );
  XOR U39920 ( .A(n36618), .B(n36619), .Z(n36251) );
  ANDN U39921 ( .B(n36620), .A(n36621), .Z(n36618) );
  AND U39922 ( .A(a[43]), .B(b[19]), .Z(n36617) );
  XOR U39923 ( .A(n36623), .B(n36624), .Z(n36256) );
  ANDN U39924 ( .B(n36625), .A(n36626), .Z(n36623) );
  AND U39925 ( .A(a[44]), .B(b[18]), .Z(n36622) );
  XOR U39926 ( .A(n36628), .B(n36629), .Z(n36261) );
  ANDN U39927 ( .B(n36630), .A(n36631), .Z(n36628) );
  AND U39928 ( .A(a[45]), .B(b[17]), .Z(n36627) );
  XOR U39929 ( .A(n36633), .B(n36634), .Z(n36266) );
  ANDN U39930 ( .B(n36635), .A(n36636), .Z(n36633) );
  AND U39931 ( .A(a[46]), .B(b[16]), .Z(n36632) );
  XOR U39932 ( .A(n36638), .B(n36639), .Z(n36271) );
  ANDN U39933 ( .B(n36640), .A(n36641), .Z(n36638) );
  AND U39934 ( .A(a[47]), .B(b[15]), .Z(n36637) );
  XOR U39935 ( .A(n36643), .B(n36644), .Z(n36276) );
  ANDN U39936 ( .B(n36645), .A(n36646), .Z(n36643) );
  AND U39937 ( .A(a[48]), .B(b[14]), .Z(n36642) );
  XOR U39938 ( .A(n36648), .B(n36649), .Z(n36281) );
  ANDN U39939 ( .B(n36650), .A(n36651), .Z(n36648) );
  AND U39940 ( .A(a[49]), .B(b[13]), .Z(n36647) );
  XOR U39941 ( .A(n36653), .B(n36654), .Z(n36286) );
  ANDN U39942 ( .B(n36655), .A(n36656), .Z(n36653) );
  AND U39943 ( .A(a[50]), .B(b[12]), .Z(n36652) );
  XOR U39944 ( .A(n36658), .B(n36659), .Z(n36291) );
  ANDN U39945 ( .B(n36660), .A(n36661), .Z(n36658) );
  AND U39946 ( .A(a[51]), .B(b[11]), .Z(n36657) );
  XOR U39947 ( .A(n36663), .B(n36664), .Z(n36296) );
  ANDN U39948 ( .B(n36665), .A(n36666), .Z(n36663) );
  AND U39949 ( .A(a[52]), .B(b[10]), .Z(n36662) );
  XOR U39950 ( .A(n36668), .B(n36669), .Z(n36301) );
  ANDN U39951 ( .B(n36670), .A(n36671), .Z(n36668) );
  AND U39952 ( .A(b[9]), .B(a[53]), .Z(n36667) );
  XOR U39953 ( .A(n36673), .B(n36674), .Z(n36306) );
  ANDN U39954 ( .B(n36675), .A(n36676), .Z(n36673) );
  AND U39955 ( .A(b[8]), .B(a[54]), .Z(n36672) );
  XOR U39956 ( .A(n36678), .B(n36679), .Z(n36311) );
  ANDN U39957 ( .B(n36680), .A(n36681), .Z(n36678) );
  AND U39958 ( .A(b[7]), .B(a[55]), .Z(n36677) );
  XOR U39959 ( .A(n36683), .B(n36684), .Z(n36316) );
  ANDN U39960 ( .B(n36685), .A(n36686), .Z(n36683) );
  AND U39961 ( .A(b[6]), .B(a[56]), .Z(n36682) );
  XOR U39962 ( .A(n36688), .B(n36689), .Z(n36321) );
  ANDN U39963 ( .B(n36690), .A(n36691), .Z(n36688) );
  AND U39964 ( .A(b[5]), .B(a[57]), .Z(n36687) );
  XOR U39965 ( .A(n36693), .B(n36694), .Z(n36326) );
  ANDN U39966 ( .B(n36695), .A(n36696), .Z(n36693) );
  AND U39967 ( .A(b[4]), .B(a[58]), .Z(n36692) );
  XOR U39968 ( .A(n36698), .B(n36699), .Z(n36331) );
  ANDN U39969 ( .B(n36343), .A(n36344), .Z(n36698) );
  AND U39970 ( .A(b[2]), .B(a[59]), .Z(n36700) );
  XNOR U39971 ( .A(n36695), .B(n36699), .Z(n36701) );
  XOR U39972 ( .A(n36702), .B(n36703), .Z(n36699) );
  OR U39973 ( .A(n36346), .B(n36347), .Z(n36703) );
  XNOR U39974 ( .A(n36705), .B(n36706), .Z(n36704) );
  XOR U39975 ( .A(n36705), .B(n36708), .Z(n36346) );
  NAND U39976 ( .A(b[1]), .B(a[59]), .Z(n36708) );
  IV U39977 ( .A(n36702), .Z(n36705) );
  NANDN U39978 ( .A(n91), .B(n92), .Z(n36702) );
  XOR U39979 ( .A(n36709), .B(n36710), .Z(n92) );
  NAND U39980 ( .A(a[59]), .B(b[0]), .Z(n91) );
  XNOR U39981 ( .A(n36690), .B(n36694), .Z(n36711) );
  XNOR U39982 ( .A(n36685), .B(n36689), .Z(n36712) );
  XNOR U39983 ( .A(n36680), .B(n36684), .Z(n36713) );
  XNOR U39984 ( .A(n36675), .B(n36679), .Z(n36714) );
  XNOR U39985 ( .A(n36670), .B(n36674), .Z(n36715) );
  XNOR U39986 ( .A(n36665), .B(n36669), .Z(n36716) );
  XNOR U39987 ( .A(n36660), .B(n36664), .Z(n36717) );
  XNOR U39988 ( .A(n36655), .B(n36659), .Z(n36718) );
  XNOR U39989 ( .A(n36650), .B(n36654), .Z(n36719) );
  XNOR U39990 ( .A(n36645), .B(n36649), .Z(n36720) );
  XNOR U39991 ( .A(n36640), .B(n36644), .Z(n36721) );
  XNOR U39992 ( .A(n36635), .B(n36639), .Z(n36722) );
  XNOR U39993 ( .A(n36630), .B(n36634), .Z(n36723) );
  XNOR U39994 ( .A(n36625), .B(n36629), .Z(n36724) );
  XNOR U39995 ( .A(n36620), .B(n36624), .Z(n36725) );
  XNOR U39996 ( .A(n36615), .B(n36619), .Z(n36726) );
  XNOR U39997 ( .A(n36610), .B(n36614), .Z(n36727) );
  XNOR U39998 ( .A(n36605), .B(n36609), .Z(n36728) );
  XNOR U39999 ( .A(n36600), .B(n36604), .Z(n36729) );
  XNOR U40000 ( .A(n36595), .B(n36599), .Z(n36730) );
  XNOR U40001 ( .A(n36590), .B(n36594), .Z(n36731) );
  XNOR U40002 ( .A(n36585), .B(n36589), .Z(n36732) );
  XNOR U40003 ( .A(n36580), .B(n36584), .Z(n36733) );
  XNOR U40004 ( .A(n36575), .B(n36579), .Z(n36734) );
  XNOR U40005 ( .A(n36570), .B(n36574), .Z(n36735) );
  XNOR U40006 ( .A(n36565), .B(n36569), .Z(n36736) );
  XNOR U40007 ( .A(n36560), .B(n36564), .Z(n36737) );
  XNOR U40008 ( .A(n36555), .B(n36559), .Z(n36738) );
  XNOR U40009 ( .A(n36550), .B(n36554), .Z(n36739) );
  XNOR U40010 ( .A(n36545), .B(n36549), .Z(n36740) );
  XNOR U40011 ( .A(n36540), .B(n36544), .Z(n36741) );
  XNOR U40012 ( .A(n36535), .B(n36539), .Z(n36742) );
  XNOR U40013 ( .A(n36530), .B(n36534), .Z(n36743) );
  XNOR U40014 ( .A(n36525), .B(n36529), .Z(n36744) );
  XNOR U40015 ( .A(n36520), .B(n36524), .Z(n36745) );
  XNOR U40016 ( .A(n36515), .B(n36519), .Z(n36746) );
  XNOR U40017 ( .A(n36510), .B(n36514), .Z(n36747) );
  XNOR U40018 ( .A(n36505), .B(n36509), .Z(n36748) );
  XNOR U40019 ( .A(n36500), .B(n36504), .Z(n36749) );
  XNOR U40020 ( .A(n36495), .B(n36499), .Z(n36750) );
  XNOR U40021 ( .A(n36490), .B(n36494), .Z(n36751) );
  XNOR U40022 ( .A(n36485), .B(n36489), .Z(n36752) );
  XNOR U40023 ( .A(n36480), .B(n36484), .Z(n36753) );
  XNOR U40024 ( .A(n36475), .B(n36479), .Z(n36754) );
  XNOR U40025 ( .A(n36470), .B(n36474), .Z(n36755) );
  XNOR U40026 ( .A(n36465), .B(n36469), .Z(n36756) );
  XNOR U40027 ( .A(n36460), .B(n36464), .Z(n36757) );
  XNOR U40028 ( .A(n36455), .B(n36459), .Z(n36758) );
  XNOR U40029 ( .A(n36450), .B(n36454), .Z(n36759) );
  XNOR U40030 ( .A(n36445), .B(n36449), .Z(n36760) );
  XNOR U40031 ( .A(n36440), .B(n36444), .Z(n36761) );
  XNOR U40032 ( .A(n36435), .B(n36439), .Z(n36762) );
  XNOR U40033 ( .A(n36430), .B(n36434), .Z(n36763) );
  XNOR U40034 ( .A(n36425), .B(n36429), .Z(n36764) );
  XNOR U40035 ( .A(n36420), .B(n36424), .Z(n36765) );
  XNOR U40036 ( .A(n36415), .B(n36419), .Z(n36766) );
  XNOR U40037 ( .A(n36410), .B(n36414), .Z(n36767) );
  XNOR U40038 ( .A(n36768), .B(n36409), .Z(n36410) );
  AND U40039 ( .A(a[0]), .B(b[61]), .Z(n36768) );
  XOR U40040 ( .A(n36769), .B(n36409), .Z(n36411) );
  XNOR U40041 ( .A(n36770), .B(n36771), .Z(n36409) );
  ANDN U40042 ( .B(n36772), .A(n36773), .Z(n36770) );
  AND U40043 ( .A(a[1]), .B(b[60]), .Z(n36769) );
  XOR U40044 ( .A(n36775), .B(n36776), .Z(n36414) );
  ANDN U40045 ( .B(n36777), .A(n36778), .Z(n36775) );
  AND U40046 ( .A(a[2]), .B(b[59]), .Z(n36774) );
  XOR U40047 ( .A(n36780), .B(n36781), .Z(n36419) );
  ANDN U40048 ( .B(n36782), .A(n36783), .Z(n36780) );
  AND U40049 ( .A(a[3]), .B(b[58]), .Z(n36779) );
  XOR U40050 ( .A(n36785), .B(n36786), .Z(n36424) );
  ANDN U40051 ( .B(n36787), .A(n36788), .Z(n36785) );
  AND U40052 ( .A(a[4]), .B(b[57]), .Z(n36784) );
  XOR U40053 ( .A(n36790), .B(n36791), .Z(n36429) );
  ANDN U40054 ( .B(n36792), .A(n36793), .Z(n36790) );
  AND U40055 ( .A(a[5]), .B(b[56]), .Z(n36789) );
  XOR U40056 ( .A(n36795), .B(n36796), .Z(n36434) );
  ANDN U40057 ( .B(n36797), .A(n36798), .Z(n36795) );
  AND U40058 ( .A(a[6]), .B(b[55]), .Z(n36794) );
  XOR U40059 ( .A(n36800), .B(n36801), .Z(n36439) );
  ANDN U40060 ( .B(n36802), .A(n36803), .Z(n36800) );
  AND U40061 ( .A(a[7]), .B(b[54]), .Z(n36799) );
  XOR U40062 ( .A(n36805), .B(n36806), .Z(n36444) );
  ANDN U40063 ( .B(n36807), .A(n36808), .Z(n36805) );
  AND U40064 ( .A(a[8]), .B(b[53]), .Z(n36804) );
  XOR U40065 ( .A(n36810), .B(n36811), .Z(n36449) );
  ANDN U40066 ( .B(n36812), .A(n36813), .Z(n36810) );
  AND U40067 ( .A(a[9]), .B(b[52]), .Z(n36809) );
  XOR U40068 ( .A(n36815), .B(n36816), .Z(n36454) );
  ANDN U40069 ( .B(n36817), .A(n36818), .Z(n36815) );
  AND U40070 ( .A(a[10]), .B(b[51]), .Z(n36814) );
  XOR U40071 ( .A(n36820), .B(n36821), .Z(n36459) );
  ANDN U40072 ( .B(n36822), .A(n36823), .Z(n36820) );
  AND U40073 ( .A(a[11]), .B(b[50]), .Z(n36819) );
  XOR U40074 ( .A(n36825), .B(n36826), .Z(n36464) );
  ANDN U40075 ( .B(n36827), .A(n36828), .Z(n36825) );
  AND U40076 ( .A(a[12]), .B(b[49]), .Z(n36824) );
  XOR U40077 ( .A(n36830), .B(n36831), .Z(n36469) );
  ANDN U40078 ( .B(n36832), .A(n36833), .Z(n36830) );
  AND U40079 ( .A(a[13]), .B(b[48]), .Z(n36829) );
  XOR U40080 ( .A(n36835), .B(n36836), .Z(n36474) );
  ANDN U40081 ( .B(n36837), .A(n36838), .Z(n36835) );
  AND U40082 ( .A(a[14]), .B(b[47]), .Z(n36834) );
  XOR U40083 ( .A(n36840), .B(n36841), .Z(n36479) );
  ANDN U40084 ( .B(n36842), .A(n36843), .Z(n36840) );
  AND U40085 ( .A(a[15]), .B(b[46]), .Z(n36839) );
  XOR U40086 ( .A(n36845), .B(n36846), .Z(n36484) );
  ANDN U40087 ( .B(n36847), .A(n36848), .Z(n36845) );
  AND U40088 ( .A(a[16]), .B(b[45]), .Z(n36844) );
  XOR U40089 ( .A(n36850), .B(n36851), .Z(n36489) );
  ANDN U40090 ( .B(n36852), .A(n36853), .Z(n36850) );
  AND U40091 ( .A(a[17]), .B(b[44]), .Z(n36849) );
  XOR U40092 ( .A(n36855), .B(n36856), .Z(n36494) );
  ANDN U40093 ( .B(n36857), .A(n36858), .Z(n36855) );
  AND U40094 ( .A(a[18]), .B(b[43]), .Z(n36854) );
  XOR U40095 ( .A(n36860), .B(n36861), .Z(n36499) );
  ANDN U40096 ( .B(n36862), .A(n36863), .Z(n36860) );
  AND U40097 ( .A(a[19]), .B(b[42]), .Z(n36859) );
  XOR U40098 ( .A(n36865), .B(n36866), .Z(n36504) );
  ANDN U40099 ( .B(n36867), .A(n36868), .Z(n36865) );
  AND U40100 ( .A(a[20]), .B(b[41]), .Z(n36864) );
  XOR U40101 ( .A(n36870), .B(n36871), .Z(n36509) );
  ANDN U40102 ( .B(n36872), .A(n36873), .Z(n36870) );
  AND U40103 ( .A(a[21]), .B(b[40]), .Z(n36869) );
  XOR U40104 ( .A(n36875), .B(n36876), .Z(n36514) );
  ANDN U40105 ( .B(n36877), .A(n36878), .Z(n36875) );
  AND U40106 ( .A(a[22]), .B(b[39]), .Z(n36874) );
  XOR U40107 ( .A(n36880), .B(n36881), .Z(n36519) );
  ANDN U40108 ( .B(n36882), .A(n36883), .Z(n36880) );
  AND U40109 ( .A(a[23]), .B(b[38]), .Z(n36879) );
  XOR U40110 ( .A(n36885), .B(n36886), .Z(n36524) );
  ANDN U40111 ( .B(n36887), .A(n36888), .Z(n36885) );
  AND U40112 ( .A(a[24]), .B(b[37]), .Z(n36884) );
  XOR U40113 ( .A(n36890), .B(n36891), .Z(n36529) );
  ANDN U40114 ( .B(n36892), .A(n36893), .Z(n36890) );
  AND U40115 ( .A(a[25]), .B(b[36]), .Z(n36889) );
  XOR U40116 ( .A(n36895), .B(n36896), .Z(n36534) );
  ANDN U40117 ( .B(n36897), .A(n36898), .Z(n36895) );
  AND U40118 ( .A(a[26]), .B(b[35]), .Z(n36894) );
  XOR U40119 ( .A(n36900), .B(n36901), .Z(n36539) );
  ANDN U40120 ( .B(n36902), .A(n36903), .Z(n36900) );
  AND U40121 ( .A(a[27]), .B(b[34]), .Z(n36899) );
  XOR U40122 ( .A(n36905), .B(n36906), .Z(n36544) );
  ANDN U40123 ( .B(n36907), .A(n36908), .Z(n36905) );
  AND U40124 ( .A(a[28]), .B(b[33]), .Z(n36904) );
  XOR U40125 ( .A(n36910), .B(n36911), .Z(n36549) );
  ANDN U40126 ( .B(n36912), .A(n36913), .Z(n36910) );
  AND U40127 ( .A(a[29]), .B(b[32]), .Z(n36909) );
  XOR U40128 ( .A(n36915), .B(n36916), .Z(n36554) );
  ANDN U40129 ( .B(n36917), .A(n36918), .Z(n36915) );
  AND U40130 ( .A(a[30]), .B(b[31]), .Z(n36914) );
  XOR U40131 ( .A(n36920), .B(n36921), .Z(n36559) );
  ANDN U40132 ( .B(n36922), .A(n36923), .Z(n36920) );
  AND U40133 ( .A(a[31]), .B(b[30]), .Z(n36919) );
  XOR U40134 ( .A(n36925), .B(n36926), .Z(n36564) );
  ANDN U40135 ( .B(n36927), .A(n36928), .Z(n36925) );
  AND U40136 ( .A(a[32]), .B(b[29]), .Z(n36924) );
  XOR U40137 ( .A(n36930), .B(n36931), .Z(n36569) );
  ANDN U40138 ( .B(n36932), .A(n36933), .Z(n36930) );
  AND U40139 ( .A(a[33]), .B(b[28]), .Z(n36929) );
  XOR U40140 ( .A(n36935), .B(n36936), .Z(n36574) );
  ANDN U40141 ( .B(n36937), .A(n36938), .Z(n36935) );
  AND U40142 ( .A(a[34]), .B(b[27]), .Z(n36934) );
  XOR U40143 ( .A(n36940), .B(n36941), .Z(n36579) );
  ANDN U40144 ( .B(n36942), .A(n36943), .Z(n36940) );
  AND U40145 ( .A(a[35]), .B(b[26]), .Z(n36939) );
  XOR U40146 ( .A(n36945), .B(n36946), .Z(n36584) );
  ANDN U40147 ( .B(n36947), .A(n36948), .Z(n36945) );
  AND U40148 ( .A(a[36]), .B(b[25]), .Z(n36944) );
  XOR U40149 ( .A(n36950), .B(n36951), .Z(n36589) );
  ANDN U40150 ( .B(n36952), .A(n36953), .Z(n36950) );
  AND U40151 ( .A(a[37]), .B(b[24]), .Z(n36949) );
  XOR U40152 ( .A(n36955), .B(n36956), .Z(n36594) );
  ANDN U40153 ( .B(n36957), .A(n36958), .Z(n36955) );
  AND U40154 ( .A(a[38]), .B(b[23]), .Z(n36954) );
  XOR U40155 ( .A(n36960), .B(n36961), .Z(n36599) );
  ANDN U40156 ( .B(n36962), .A(n36963), .Z(n36960) );
  AND U40157 ( .A(a[39]), .B(b[22]), .Z(n36959) );
  XOR U40158 ( .A(n36965), .B(n36966), .Z(n36604) );
  ANDN U40159 ( .B(n36967), .A(n36968), .Z(n36965) );
  AND U40160 ( .A(a[40]), .B(b[21]), .Z(n36964) );
  XOR U40161 ( .A(n36970), .B(n36971), .Z(n36609) );
  ANDN U40162 ( .B(n36972), .A(n36973), .Z(n36970) );
  AND U40163 ( .A(a[41]), .B(b[20]), .Z(n36969) );
  XOR U40164 ( .A(n36975), .B(n36976), .Z(n36614) );
  ANDN U40165 ( .B(n36977), .A(n36978), .Z(n36975) );
  AND U40166 ( .A(a[42]), .B(b[19]), .Z(n36974) );
  XOR U40167 ( .A(n36980), .B(n36981), .Z(n36619) );
  ANDN U40168 ( .B(n36982), .A(n36983), .Z(n36980) );
  AND U40169 ( .A(a[43]), .B(b[18]), .Z(n36979) );
  XOR U40170 ( .A(n36985), .B(n36986), .Z(n36624) );
  ANDN U40171 ( .B(n36987), .A(n36988), .Z(n36985) );
  AND U40172 ( .A(a[44]), .B(b[17]), .Z(n36984) );
  XOR U40173 ( .A(n36990), .B(n36991), .Z(n36629) );
  ANDN U40174 ( .B(n36992), .A(n36993), .Z(n36990) );
  AND U40175 ( .A(a[45]), .B(b[16]), .Z(n36989) );
  XOR U40176 ( .A(n36995), .B(n36996), .Z(n36634) );
  ANDN U40177 ( .B(n36997), .A(n36998), .Z(n36995) );
  AND U40178 ( .A(a[46]), .B(b[15]), .Z(n36994) );
  XOR U40179 ( .A(n37000), .B(n37001), .Z(n36639) );
  ANDN U40180 ( .B(n37002), .A(n37003), .Z(n37000) );
  AND U40181 ( .A(a[47]), .B(b[14]), .Z(n36999) );
  XOR U40182 ( .A(n37005), .B(n37006), .Z(n36644) );
  ANDN U40183 ( .B(n37007), .A(n37008), .Z(n37005) );
  AND U40184 ( .A(a[48]), .B(b[13]), .Z(n37004) );
  XOR U40185 ( .A(n37010), .B(n37011), .Z(n36649) );
  ANDN U40186 ( .B(n37012), .A(n37013), .Z(n37010) );
  AND U40187 ( .A(a[49]), .B(b[12]), .Z(n37009) );
  XOR U40188 ( .A(n37015), .B(n37016), .Z(n36654) );
  ANDN U40189 ( .B(n37017), .A(n37018), .Z(n37015) );
  AND U40190 ( .A(a[50]), .B(b[11]), .Z(n37014) );
  XOR U40191 ( .A(n37020), .B(n37021), .Z(n36659) );
  ANDN U40192 ( .B(n37022), .A(n37023), .Z(n37020) );
  AND U40193 ( .A(a[51]), .B(b[10]), .Z(n37019) );
  XOR U40194 ( .A(n37025), .B(n37026), .Z(n36664) );
  ANDN U40195 ( .B(n37027), .A(n37028), .Z(n37025) );
  AND U40196 ( .A(b[9]), .B(a[52]), .Z(n37024) );
  XOR U40197 ( .A(n37030), .B(n37031), .Z(n36669) );
  ANDN U40198 ( .B(n37032), .A(n37033), .Z(n37030) );
  AND U40199 ( .A(b[8]), .B(a[53]), .Z(n37029) );
  XOR U40200 ( .A(n37035), .B(n37036), .Z(n36674) );
  ANDN U40201 ( .B(n37037), .A(n37038), .Z(n37035) );
  AND U40202 ( .A(b[7]), .B(a[54]), .Z(n37034) );
  XOR U40203 ( .A(n37040), .B(n37041), .Z(n36679) );
  ANDN U40204 ( .B(n37042), .A(n37043), .Z(n37040) );
  AND U40205 ( .A(b[6]), .B(a[55]), .Z(n37039) );
  XOR U40206 ( .A(n37045), .B(n37046), .Z(n36684) );
  ANDN U40207 ( .B(n37047), .A(n37048), .Z(n37045) );
  AND U40208 ( .A(b[5]), .B(a[56]), .Z(n37044) );
  XOR U40209 ( .A(n37050), .B(n37051), .Z(n36689) );
  ANDN U40210 ( .B(n37052), .A(n37053), .Z(n37050) );
  AND U40211 ( .A(b[4]), .B(a[57]), .Z(n37049) );
  XOR U40212 ( .A(n37055), .B(n37056), .Z(n36694) );
  ANDN U40213 ( .B(n36706), .A(n36707), .Z(n37055) );
  AND U40214 ( .A(b[2]), .B(a[58]), .Z(n37057) );
  XNOR U40215 ( .A(n37052), .B(n37056), .Z(n37058) );
  XOR U40216 ( .A(n37059), .B(n37060), .Z(n37056) );
  OR U40217 ( .A(n36709), .B(n36710), .Z(n37060) );
  XNOR U40218 ( .A(n37062), .B(n37063), .Z(n37061) );
  XOR U40219 ( .A(n37062), .B(n37065), .Z(n36709) );
  NAND U40220 ( .A(b[1]), .B(a[58]), .Z(n37065) );
  IV U40221 ( .A(n37059), .Z(n37062) );
  NANDN U40222 ( .A(n93), .B(n94), .Z(n37059) );
  XOR U40223 ( .A(n37066), .B(n37067), .Z(n94) );
  NAND U40224 ( .A(a[58]), .B(b[0]), .Z(n93) );
  XNOR U40225 ( .A(n37047), .B(n37051), .Z(n37068) );
  XNOR U40226 ( .A(n37042), .B(n37046), .Z(n37069) );
  XNOR U40227 ( .A(n37037), .B(n37041), .Z(n37070) );
  XNOR U40228 ( .A(n37032), .B(n37036), .Z(n37071) );
  XNOR U40229 ( .A(n37027), .B(n37031), .Z(n37072) );
  XNOR U40230 ( .A(n37022), .B(n37026), .Z(n37073) );
  XNOR U40231 ( .A(n37017), .B(n37021), .Z(n37074) );
  XNOR U40232 ( .A(n37012), .B(n37016), .Z(n37075) );
  XNOR U40233 ( .A(n37007), .B(n37011), .Z(n37076) );
  XNOR U40234 ( .A(n37002), .B(n37006), .Z(n37077) );
  XNOR U40235 ( .A(n36997), .B(n37001), .Z(n37078) );
  XNOR U40236 ( .A(n36992), .B(n36996), .Z(n37079) );
  XNOR U40237 ( .A(n36987), .B(n36991), .Z(n37080) );
  XNOR U40238 ( .A(n36982), .B(n36986), .Z(n37081) );
  XNOR U40239 ( .A(n36977), .B(n36981), .Z(n37082) );
  XNOR U40240 ( .A(n36972), .B(n36976), .Z(n37083) );
  XNOR U40241 ( .A(n36967), .B(n36971), .Z(n37084) );
  XNOR U40242 ( .A(n36962), .B(n36966), .Z(n37085) );
  XNOR U40243 ( .A(n36957), .B(n36961), .Z(n37086) );
  XNOR U40244 ( .A(n36952), .B(n36956), .Z(n37087) );
  XNOR U40245 ( .A(n36947), .B(n36951), .Z(n37088) );
  XNOR U40246 ( .A(n36942), .B(n36946), .Z(n37089) );
  XNOR U40247 ( .A(n36937), .B(n36941), .Z(n37090) );
  XNOR U40248 ( .A(n36932), .B(n36936), .Z(n37091) );
  XNOR U40249 ( .A(n36927), .B(n36931), .Z(n37092) );
  XNOR U40250 ( .A(n36922), .B(n36926), .Z(n37093) );
  XNOR U40251 ( .A(n36917), .B(n36921), .Z(n37094) );
  XNOR U40252 ( .A(n36912), .B(n36916), .Z(n37095) );
  XNOR U40253 ( .A(n36907), .B(n36911), .Z(n37096) );
  XNOR U40254 ( .A(n36902), .B(n36906), .Z(n37097) );
  XNOR U40255 ( .A(n36897), .B(n36901), .Z(n37098) );
  XNOR U40256 ( .A(n36892), .B(n36896), .Z(n37099) );
  XNOR U40257 ( .A(n36887), .B(n36891), .Z(n37100) );
  XNOR U40258 ( .A(n36882), .B(n36886), .Z(n37101) );
  XNOR U40259 ( .A(n36877), .B(n36881), .Z(n37102) );
  XNOR U40260 ( .A(n36872), .B(n36876), .Z(n37103) );
  XNOR U40261 ( .A(n36867), .B(n36871), .Z(n37104) );
  XNOR U40262 ( .A(n36862), .B(n36866), .Z(n37105) );
  XNOR U40263 ( .A(n36857), .B(n36861), .Z(n37106) );
  XNOR U40264 ( .A(n36852), .B(n36856), .Z(n37107) );
  XNOR U40265 ( .A(n36847), .B(n36851), .Z(n37108) );
  XNOR U40266 ( .A(n36842), .B(n36846), .Z(n37109) );
  XNOR U40267 ( .A(n36837), .B(n36841), .Z(n37110) );
  XNOR U40268 ( .A(n36832), .B(n36836), .Z(n37111) );
  XNOR U40269 ( .A(n36827), .B(n36831), .Z(n37112) );
  XNOR U40270 ( .A(n36822), .B(n36826), .Z(n37113) );
  XNOR U40271 ( .A(n36817), .B(n36821), .Z(n37114) );
  XNOR U40272 ( .A(n36812), .B(n36816), .Z(n37115) );
  XNOR U40273 ( .A(n36807), .B(n36811), .Z(n37116) );
  XNOR U40274 ( .A(n36802), .B(n36806), .Z(n37117) );
  XNOR U40275 ( .A(n36797), .B(n36801), .Z(n37118) );
  XNOR U40276 ( .A(n36792), .B(n36796), .Z(n37119) );
  XNOR U40277 ( .A(n36787), .B(n36791), .Z(n37120) );
  XNOR U40278 ( .A(n36782), .B(n36786), .Z(n37121) );
  XNOR U40279 ( .A(n36777), .B(n36781), .Z(n37122) );
  XNOR U40280 ( .A(n36772), .B(n36776), .Z(n37123) );
  XOR U40281 ( .A(n37124), .B(n36771), .Z(n36772) );
  AND U40282 ( .A(a[0]), .B(b[60]), .Z(n37124) );
  XNOR U40283 ( .A(n37125), .B(n36771), .Z(n36773) );
  XNOR U40284 ( .A(n37126), .B(n37127), .Z(n36771) );
  ANDN U40285 ( .B(n37128), .A(n37129), .Z(n37126) );
  AND U40286 ( .A(a[1]), .B(b[59]), .Z(n37125) );
  XOR U40287 ( .A(n37131), .B(n37132), .Z(n36776) );
  ANDN U40288 ( .B(n37133), .A(n37134), .Z(n37131) );
  AND U40289 ( .A(a[2]), .B(b[58]), .Z(n37130) );
  XOR U40290 ( .A(n37136), .B(n37137), .Z(n36781) );
  ANDN U40291 ( .B(n37138), .A(n37139), .Z(n37136) );
  AND U40292 ( .A(a[3]), .B(b[57]), .Z(n37135) );
  XOR U40293 ( .A(n37141), .B(n37142), .Z(n36786) );
  ANDN U40294 ( .B(n37143), .A(n37144), .Z(n37141) );
  AND U40295 ( .A(a[4]), .B(b[56]), .Z(n37140) );
  XOR U40296 ( .A(n37146), .B(n37147), .Z(n36791) );
  ANDN U40297 ( .B(n37148), .A(n37149), .Z(n37146) );
  AND U40298 ( .A(a[5]), .B(b[55]), .Z(n37145) );
  XOR U40299 ( .A(n37151), .B(n37152), .Z(n36796) );
  ANDN U40300 ( .B(n37153), .A(n37154), .Z(n37151) );
  AND U40301 ( .A(a[6]), .B(b[54]), .Z(n37150) );
  XOR U40302 ( .A(n37156), .B(n37157), .Z(n36801) );
  ANDN U40303 ( .B(n37158), .A(n37159), .Z(n37156) );
  AND U40304 ( .A(a[7]), .B(b[53]), .Z(n37155) );
  XOR U40305 ( .A(n37161), .B(n37162), .Z(n36806) );
  ANDN U40306 ( .B(n37163), .A(n37164), .Z(n37161) );
  AND U40307 ( .A(a[8]), .B(b[52]), .Z(n37160) );
  XOR U40308 ( .A(n37166), .B(n37167), .Z(n36811) );
  ANDN U40309 ( .B(n37168), .A(n37169), .Z(n37166) );
  AND U40310 ( .A(a[9]), .B(b[51]), .Z(n37165) );
  XOR U40311 ( .A(n37171), .B(n37172), .Z(n36816) );
  ANDN U40312 ( .B(n37173), .A(n37174), .Z(n37171) );
  AND U40313 ( .A(a[10]), .B(b[50]), .Z(n37170) );
  XOR U40314 ( .A(n37176), .B(n37177), .Z(n36821) );
  ANDN U40315 ( .B(n37178), .A(n37179), .Z(n37176) );
  AND U40316 ( .A(a[11]), .B(b[49]), .Z(n37175) );
  XOR U40317 ( .A(n37181), .B(n37182), .Z(n36826) );
  ANDN U40318 ( .B(n37183), .A(n37184), .Z(n37181) );
  AND U40319 ( .A(a[12]), .B(b[48]), .Z(n37180) );
  XOR U40320 ( .A(n37186), .B(n37187), .Z(n36831) );
  ANDN U40321 ( .B(n37188), .A(n37189), .Z(n37186) );
  AND U40322 ( .A(a[13]), .B(b[47]), .Z(n37185) );
  XOR U40323 ( .A(n37191), .B(n37192), .Z(n36836) );
  ANDN U40324 ( .B(n37193), .A(n37194), .Z(n37191) );
  AND U40325 ( .A(a[14]), .B(b[46]), .Z(n37190) );
  XOR U40326 ( .A(n37196), .B(n37197), .Z(n36841) );
  ANDN U40327 ( .B(n37198), .A(n37199), .Z(n37196) );
  AND U40328 ( .A(a[15]), .B(b[45]), .Z(n37195) );
  XOR U40329 ( .A(n37201), .B(n37202), .Z(n36846) );
  ANDN U40330 ( .B(n37203), .A(n37204), .Z(n37201) );
  AND U40331 ( .A(a[16]), .B(b[44]), .Z(n37200) );
  XOR U40332 ( .A(n37206), .B(n37207), .Z(n36851) );
  ANDN U40333 ( .B(n37208), .A(n37209), .Z(n37206) );
  AND U40334 ( .A(a[17]), .B(b[43]), .Z(n37205) );
  XOR U40335 ( .A(n37211), .B(n37212), .Z(n36856) );
  ANDN U40336 ( .B(n37213), .A(n37214), .Z(n37211) );
  AND U40337 ( .A(a[18]), .B(b[42]), .Z(n37210) );
  XOR U40338 ( .A(n37216), .B(n37217), .Z(n36861) );
  ANDN U40339 ( .B(n37218), .A(n37219), .Z(n37216) );
  AND U40340 ( .A(a[19]), .B(b[41]), .Z(n37215) );
  XOR U40341 ( .A(n37221), .B(n37222), .Z(n36866) );
  ANDN U40342 ( .B(n37223), .A(n37224), .Z(n37221) );
  AND U40343 ( .A(a[20]), .B(b[40]), .Z(n37220) );
  XOR U40344 ( .A(n37226), .B(n37227), .Z(n36871) );
  ANDN U40345 ( .B(n37228), .A(n37229), .Z(n37226) );
  AND U40346 ( .A(a[21]), .B(b[39]), .Z(n37225) );
  XOR U40347 ( .A(n37231), .B(n37232), .Z(n36876) );
  ANDN U40348 ( .B(n37233), .A(n37234), .Z(n37231) );
  AND U40349 ( .A(a[22]), .B(b[38]), .Z(n37230) );
  XOR U40350 ( .A(n37236), .B(n37237), .Z(n36881) );
  ANDN U40351 ( .B(n37238), .A(n37239), .Z(n37236) );
  AND U40352 ( .A(a[23]), .B(b[37]), .Z(n37235) );
  XOR U40353 ( .A(n37241), .B(n37242), .Z(n36886) );
  ANDN U40354 ( .B(n37243), .A(n37244), .Z(n37241) );
  AND U40355 ( .A(a[24]), .B(b[36]), .Z(n37240) );
  XOR U40356 ( .A(n37246), .B(n37247), .Z(n36891) );
  ANDN U40357 ( .B(n37248), .A(n37249), .Z(n37246) );
  AND U40358 ( .A(a[25]), .B(b[35]), .Z(n37245) );
  XOR U40359 ( .A(n37251), .B(n37252), .Z(n36896) );
  ANDN U40360 ( .B(n37253), .A(n37254), .Z(n37251) );
  AND U40361 ( .A(a[26]), .B(b[34]), .Z(n37250) );
  XOR U40362 ( .A(n37256), .B(n37257), .Z(n36901) );
  ANDN U40363 ( .B(n37258), .A(n37259), .Z(n37256) );
  AND U40364 ( .A(a[27]), .B(b[33]), .Z(n37255) );
  XOR U40365 ( .A(n37261), .B(n37262), .Z(n36906) );
  ANDN U40366 ( .B(n37263), .A(n37264), .Z(n37261) );
  AND U40367 ( .A(a[28]), .B(b[32]), .Z(n37260) );
  XOR U40368 ( .A(n37266), .B(n37267), .Z(n36911) );
  ANDN U40369 ( .B(n37268), .A(n37269), .Z(n37266) );
  AND U40370 ( .A(a[29]), .B(b[31]), .Z(n37265) );
  XOR U40371 ( .A(n37271), .B(n37272), .Z(n36916) );
  ANDN U40372 ( .B(n37273), .A(n37274), .Z(n37271) );
  AND U40373 ( .A(a[30]), .B(b[30]), .Z(n37270) );
  XOR U40374 ( .A(n37276), .B(n37277), .Z(n36921) );
  ANDN U40375 ( .B(n37278), .A(n37279), .Z(n37276) );
  AND U40376 ( .A(a[31]), .B(b[29]), .Z(n37275) );
  XOR U40377 ( .A(n37281), .B(n37282), .Z(n36926) );
  ANDN U40378 ( .B(n37283), .A(n37284), .Z(n37281) );
  AND U40379 ( .A(a[32]), .B(b[28]), .Z(n37280) );
  XOR U40380 ( .A(n37286), .B(n37287), .Z(n36931) );
  ANDN U40381 ( .B(n37288), .A(n37289), .Z(n37286) );
  AND U40382 ( .A(a[33]), .B(b[27]), .Z(n37285) );
  XOR U40383 ( .A(n37291), .B(n37292), .Z(n36936) );
  ANDN U40384 ( .B(n37293), .A(n37294), .Z(n37291) );
  AND U40385 ( .A(a[34]), .B(b[26]), .Z(n37290) );
  XOR U40386 ( .A(n37296), .B(n37297), .Z(n36941) );
  ANDN U40387 ( .B(n37298), .A(n37299), .Z(n37296) );
  AND U40388 ( .A(a[35]), .B(b[25]), .Z(n37295) );
  XOR U40389 ( .A(n37301), .B(n37302), .Z(n36946) );
  ANDN U40390 ( .B(n37303), .A(n37304), .Z(n37301) );
  AND U40391 ( .A(a[36]), .B(b[24]), .Z(n37300) );
  XOR U40392 ( .A(n37306), .B(n37307), .Z(n36951) );
  ANDN U40393 ( .B(n37308), .A(n37309), .Z(n37306) );
  AND U40394 ( .A(a[37]), .B(b[23]), .Z(n37305) );
  XOR U40395 ( .A(n37311), .B(n37312), .Z(n36956) );
  ANDN U40396 ( .B(n37313), .A(n37314), .Z(n37311) );
  AND U40397 ( .A(a[38]), .B(b[22]), .Z(n37310) );
  XOR U40398 ( .A(n37316), .B(n37317), .Z(n36961) );
  ANDN U40399 ( .B(n37318), .A(n37319), .Z(n37316) );
  AND U40400 ( .A(a[39]), .B(b[21]), .Z(n37315) );
  XOR U40401 ( .A(n37321), .B(n37322), .Z(n36966) );
  ANDN U40402 ( .B(n37323), .A(n37324), .Z(n37321) );
  AND U40403 ( .A(a[40]), .B(b[20]), .Z(n37320) );
  XOR U40404 ( .A(n37326), .B(n37327), .Z(n36971) );
  ANDN U40405 ( .B(n37328), .A(n37329), .Z(n37326) );
  AND U40406 ( .A(a[41]), .B(b[19]), .Z(n37325) );
  XOR U40407 ( .A(n37331), .B(n37332), .Z(n36976) );
  ANDN U40408 ( .B(n37333), .A(n37334), .Z(n37331) );
  AND U40409 ( .A(a[42]), .B(b[18]), .Z(n37330) );
  XOR U40410 ( .A(n37336), .B(n37337), .Z(n36981) );
  ANDN U40411 ( .B(n37338), .A(n37339), .Z(n37336) );
  AND U40412 ( .A(a[43]), .B(b[17]), .Z(n37335) );
  XOR U40413 ( .A(n37341), .B(n37342), .Z(n36986) );
  ANDN U40414 ( .B(n37343), .A(n37344), .Z(n37341) );
  AND U40415 ( .A(a[44]), .B(b[16]), .Z(n37340) );
  XOR U40416 ( .A(n37346), .B(n37347), .Z(n36991) );
  ANDN U40417 ( .B(n37348), .A(n37349), .Z(n37346) );
  AND U40418 ( .A(a[45]), .B(b[15]), .Z(n37345) );
  XOR U40419 ( .A(n37351), .B(n37352), .Z(n36996) );
  ANDN U40420 ( .B(n37353), .A(n37354), .Z(n37351) );
  AND U40421 ( .A(a[46]), .B(b[14]), .Z(n37350) );
  XOR U40422 ( .A(n37356), .B(n37357), .Z(n37001) );
  ANDN U40423 ( .B(n37358), .A(n37359), .Z(n37356) );
  AND U40424 ( .A(a[47]), .B(b[13]), .Z(n37355) );
  XOR U40425 ( .A(n37361), .B(n37362), .Z(n37006) );
  ANDN U40426 ( .B(n37363), .A(n37364), .Z(n37361) );
  AND U40427 ( .A(a[48]), .B(b[12]), .Z(n37360) );
  XOR U40428 ( .A(n37366), .B(n37367), .Z(n37011) );
  ANDN U40429 ( .B(n37368), .A(n37369), .Z(n37366) );
  AND U40430 ( .A(a[49]), .B(b[11]), .Z(n37365) );
  XOR U40431 ( .A(n37371), .B(n37372), .Z(n37016) );
  ANDN U40432 ( .B(n37373), .A(n37374), .Z(n37371) );
  AND U40433 ( .A(a[50]), .B(b[10]), .Z(n37370) );
  XOR U40434 ( .A(n37376), .B(n37377), .Z(n37021) );
  ANDN U40435 ( .B(n37378), .A(n37379), .Z(n37376) );
  AND U40436 ( .A(b[9]), .B(a[51]), .Z(n37375) );
  XOR U40437 ( .A(n37381), .B(n37382), .Z(n37026) );
  ANDN U40438 ( .B(n37383), .A(n37384), .Z(n37381) );
  AND U40439 ( .A(b[8]), .B(a[52]), .Z(n37380) );
  XOR U40440 ( .A(n37386), .B(n37387), .Z(n37031) );
  ANDN U40441 ( .B(n37388), .A(n37389), .Z(n37386) );
  AND U40442 ( .A(b[7]), .B(a[53]), .Z(n37385) );
  XOR U40443 ( .A(n37391), .B(n37392), .Z(n37036) );
  ANDN U40444 ( .B(n37393), .A(n37394), .Z(n37391) );
  AND U40445 ( .A(b[6]), .B(a[54]), .Z(n37390) );
  XOR U40446 ( .A(n37396), .B(n37397), .Z(n37041) );
  ANDN U40447 ( .B(n37398), .A(n37399), .Z(n37396) );
  AND U40448 ( .A(b[5]), .B(a[55]), .Z(n37395) );
  XOR U40449 ( .A(n37401), .B(n37402), .Z(n37046) );
  ANDN U40450 ( .B(n37403), .A(n37404), .Z(n37401) );
  AND U40451 ( .A(b[4]), .B(a[56]), .Z(n37400) );
  XOR U40452 ( .A(n37406), .B(n37407), .Z(n37051) );
  ANDN U40453 ( .B(n37063), .A(n37064), .Z(n37406) );
  AND U40454 ( .A(b[2]), .B(a[57]), .Z(n37408) );
  XNOR U40455 ( .A(n37403), .B(n37407), .Z(n37409) );
  XOR U40456 ( .A(n37410), .B(n37411), .Z(n37407) );
  OR U40457 ( .A(n37066), .B(n37067), .Z(n37411) );
  XNOR U40458 ( .A(n37413), .B(n37414), .Z(n37412) );
  XOR U40459 ( .A(n37413), .B(n37416), .Z(n37066) );
  NAND U40460 ( .A(b[1]), .B(a[57]), .Z(n37416) );
  IV U40461 ( .A(n37410), .Z(n37413) );
  NANDN U40462 ( .A(n95), .B(n96), .Z(n37410) );
  XOR U40463 ( .A(n37417), .B(n37418), .Z(n96) );
  NAND U40464 ( .A(a[57]), .B(b[0]), .Z(n95) );
  XNOR U40465 ( .A(n37398), .B(n37402), .Z(n37419) );
  XNOR U40466 ( .A(n37393), .B(n37397), .Z(n37420) );
  XNOR U40467 ( .A(n37388), .B(n37392), .Z(n37421) );
  XNOR U40468 ( .A(n37383), .B(n37387), .Z(n37422) );
  XNOR U40469 ( .A(n37378), .B(n37382), .Z(n37423) );
  XNOR U40470 ( .A(n37373), .B(n37377), .Z(n37424) );
  XNOR U40471 ( .A(n37368), .B(n37372), .Z(n37425) );
  XNOR U40472 ( .A(n37363), .B(n37367), .Z(n37426) );
  XNOR U40473 ( .A(n37358), .B(n37362), .Z(n37427) );
  XNOR U40474 ( .A(n37353), .B(n37357), .Z(n37428) );
  XNOR U40475 ( .A(n37348), .B(n37352), .Z(n37429) );
  XNOR U40476 ( .A(n37343), .B(n37347), .Z(n37430) );
  XNOR U40477 ( .A(n37338), .B(n37342), .Z(n37431) );
  XNOR U40478 ( .A(n37333), .B(n37337), .Z(n37432) );
  XNOR U40479 ( .A(n37328), .B(n37332), .Z(n37433) );
  XNOR U40480 ( .A(n37323), .B(n37327), .Z(n37434) );
  XNOR U40481 ( .A(n37318), .B(n37322), .Z(n37435) );
  XNOR U40482 ( .A(n37313), .B(n37317), .Z(n37436) );
  XNOR U40483 ( .A(n37308), .B(n37312), .Z(n37437) );
  XNOR U40484 ( .A(n37303), .B(n37307), .Z(n37438) );
  XNOR U40485 ( .A(n37298), .B(n37302), .Z(n37439) );
  XNOR U40486 ( .A(n37293), .B(n37297), .Z(n37440) );
  XNOR U40487 ( .A(n37288), .B(n37292), .Z(n37441) );
  XNOR U40488 ( .A(n37283), .B(n37287), .Z(n37442) );
  XNOR U40489 ( .A(n37278), .B(n37282), .Z(n37443) );
  XNOR U40490 ( .A(n37273), .B(n37277), .Z(n37444) );
  XNOR U40491 ( .A(n37268), .B(n37272), .Z(n37445) );
  XNOR U40492 ( .A(n37263), .B(n37267), .Z(n37446) );
  XNOR U40493 ( .A(n37258), .B(n37262), .Z(n37447) );
  XNOR U40494 ( .A(n37253), .B(n37257), .Z(n37448) );
  XNOR U40495 ( .A(n37248), .B(n37252), .Z(n37449) );
  XNOR U40496 ( .A(n37243), .B(n37247), .Z(n37450) );
  XNOR U40497 ( .A(n37238), .B(n37242), .Z(n37451) );
  XNOR U40498 ( .A(n37233), .B(n37237), .Z(n37452) );
  XNOR U40499 ( .A(n37228), .B(n37232), .Z(n37453) );
  XNOR U40500 ( .A(n37223), .B(n37227), .Z(n37454) );
  XNOR U40501 ( .A(n37218), .B(n37222), .Z(n37455) );
  XNOR U40502 ( .A(n37213), .B(n37217), .Z(n37456) );
  XNOR U40503 ( .A(n37208), .B(n37212), .Z(n37457) );
  XNOR U40504 ( .A(n37203), .B(n37207), .Z(n37458) );
  XNOR U40505 ( .A(n37198), .B(n37202), .Z(n37459) );
  XNOR U40506 ( .A(n37193), .B(n37197), .Z(n37460) );
  XNOR U40507 ( .A(n37188), .B(n37192), .Z(n37461) );
  XNOR U40508 ( .A(n37183), .B(n37187), .Z(n37462) );
  XNOR U40509 ( .A(n37178), .B(n37182), .Z(n37463) );
  XNOR U40510 ( .A(n37173), .B(n37177), .Z(n37464) );
  XNOR U40511 ( .A(n37168), .B(n37172), .Z(n37465) );
  XNOR U40512 ( .A(n37163), .B(n37167), .Z(n37466) );
  XNOR U40513 ( .A(n37158), .B(n37162), .Z(n37467) );
  XNOR U40514 ( .A(n37153), .B(n37157), .Z(n37468) );
  XNOR U40515 ( .A(n37148), .B(n37152), .Z(n37469) );
  XNOR U40516 ( .A(n37143), .B(n37147), .Z(n37470) );
  XNOR U40517 ( .A(n37138), .B(n37142), .Z(n37471) );
  XNOR U40518 ( .A(n37133), .B(n37137), .Z(n37472) );
  XNOR U40519 ( .A(n37128), .B(n37132), .Z(n37473) );
  XNOR U40520 ( .A(n37474), .B(n37127), .Z(n37128) );
  AND U40521 ( .A(a[0]), .B(b[59]), .Z(n37474) );
  XOR U40522 ( .A(n37475), .B(n37127), .Z(n37129) );
  XNOR U40523 ( .A(n37476), .B(n37477), .Z(n37127) );
  ANDN U40524 ( .B(n37478), .A(n37479), .Z(n37476) );
  AND U40525 ( .A(a[1]), .B(b[58]), .Z(n37475) );
  XOR U40526 ( .A(n37481), .B(n37482), .Z(n37132) );
  ANDN U40527 ( .B(n37483), .A(n37484), .Z(n37481) );
  AND U40528 ( .A(a[2]), .B(b[57]), .Z(n37480) );
  XOR U40529 ( .A(n37486), .B(n37487), .Z(n37137) );
  ANDN U40530 ( .B(n37488), .A(n37489), .Z(n37486) );
  AND U40531 ( .A(a[3]), .B(b[56]), .Z(n37485) );
  XOR U40532 ( .A(n37491), .B(n37492), .Z(n37142) );
  ANDN U40533 ( .B(n37493), .A(n37494), .Z(n37491) );
  AND U40534 ( .A(a[4]), .B(b[55]), .Z(n37490) );
  XOR U40535 ( .A(n37496), .B(n37497), .Z(n37147) );
  ANDN U40536 ( .B(n37498), .A(n37499), .Z(n37496) );
  AND U40537 ( .A(a[5]), .B(b[54]), .Z(n37495) );
  XOR U40538 ( .A(n37501), .B(n37502), .Z(n37152) );
  ANDN U40539 ( .B(n37503), .A(n37504), .Z(n37501) );
  AND U40540 ( .A(a[6]), .B(b[53]), .Z(n37500) );
  XOR U40541 ( .A(n37506), .B(n37507), .Z(n37157) );
  ANDN U40542 ( .B(n37508), .A(n37509), .Z(n37506) );
  AND U40543 ( .A(a[7]), .B(b[52]), .Z(n37505) );
  XOR U40544 ( .A(n37511), .B(n37512), .Z(n37162) );
  ANDN U40545 ( .B(n37513), .A(n37514), .Z(n37511) );
  AND U40546 ( .A(a[8]), .B(b[51]), .Z(n37510) );
  XOR U40547 ( .A(n37516), .B(n37517), .Z(n37167) );
  ANDN U40548 ( .B(n37518), .A(n37519), .Z(n37516) );
  AND U40549 ( .A(a[9]), .B(b[50]), .Z(n37515) );
  XOR U40550 ( .A(n37521), .B(n37522), .Z(n37172) );
  ANDN U40551 ( .B(n37523), .A(n37524), .Z(n37521) );
  AND U40552 ( .A(a[10]), .B(b[49]), .Z(n37520) );
  XOR U40553 ( .A(n37526), .B(n37527), .Z(n37177) );
  ANDN U40554 ( .B(n37528), .A(n37529), .Z(n37526) );
  AND U40555 ( .A(a[11]), .B(b[48]), .Z(n37525) );
  XOR U40556 ( .A(n37531), .B(n37532), .Z(n37182) );
  ANDN U40557 ( .B(n37533), .A(n37534), .Z(n37531) );
  AND U40558 ( .A(a[12]), .B(b[47]), .Z(n37530) );
  XOR U40559 ( .A(n37536), .B(n37537), .Z(n37187) );
  ANDN U40560 ( .B(n37538), .A(n37539), .Z(n37536) );
  AND U40561 ( .A(a[13]), .B(b[46]), .Z(n37535) );
  XOR U40562 ( .A(n37541), .B(n37542), .Z(n37192) );
  ANDN U40563 ( .B(n37543), .A(n37544), .Z(n37541) );
  AND U40564 ( .A(a[14]), .B(b[45]), .Z(n37540) );
  XOR U40565 ( .A(n37546), .B(n37547), .Z(n37197) );
  ANDN U40566 ( .B(n37548), .A(n37549), .Z(n37546) );
  AND U40567 ( .A(a[15]), .B(b[44]), .Z(n37545) );
  XOR U40568 ( .A(n37551), .B(n37552), .Z(n37202) );
  ANDN U40569 ( .B(n37553), .A(n37554), .Z(n37551) );
  AND U40570 ( .A(a[16]), .B(b[43]), .Z(n37550) );
  XOR U40571 ( .A(n37556), .B(n37557), .Z(n37207) );
  ANDN U40572 ( .B(n37558), .A(n37559), .Z(n37556) );
  AND U40573 ( .A(a[17]), .B(b[42]), .Z(n37555) );
  XOR U40574 ( .A(n37561), .B(n37562), .Z(n37212) );
  ANDN U40575 ( .B(n37563), .A(n37564), .Z(n37561) );
  AND U40576 ( .A(a[18]), .B(b[41]), .Z(n37560) );
  XOR U40577 ( .A(n37566), .B(n37567), .Z(n37217) );
  ANDN U40578 ( .B(n37568), .A(n37569), .Z(n37566) );
  AND U40579 ( .A(a[19]), .B(b[40]), .Z(n37565) );
  XOR U40580 ( .A(n37571), .B(n37572), .Z(n37222) );
  ANDN U40581 ( .B(n37573), .A(n37574), .Z(n37571) );
  AND U40582 ( .A(a[20]), .B(b[39]), .Z(n37570) );
  XOR U40583 ( .A(n37576), .B(n37577), .Z(n37227) );
  ANDN U40584 ( .B(n37578), .A(n37579), .Z(n37576) );
  AND U40585 ( .A(a[21]), .B(b[38]), .Z(n37575) );
  XOR U40586 ( .A(n37581), .B(n37582), .Z(n37232) );
  ANDN U40587 ( .B(n37583), .A(n37584), .Z(n37581) );
  AND U40588 ( .A(a[22]), .B(b[37]), .Z(n37580) );
  XOR U40589 ( .A(n37586), .B(n37587), .Z(n37237) );
  ANDN U40590 ( .B(n37588), .A(n37589), .Z(n37586) );
  AND U40591 ( .A(a[23]), .B(b[36]), .Z(n37585) );
  XOR U40592 ( .A(n37591), .B(n37592), .Z(n37242) );
  ANDN U40593 ( .B(n37593), .A(n37594), .Z(n37591) );
  AND U40594 ( .A(a[24]), .B(b[35]), .Z(n37590) );
  XOR U40595 ( .A(n37596), .B(n37597), .Z(n37247) );
  ANDN U40596 ( .B(n37598), .A(n37599), .Z(n37596) );
  AND U40597 ( .A(a[25]), .B(b[34]), .Z(n37595) );
  XOR U40598 ( .A(n37601), .B(n37602), .Z(n37252) );
  ANDN U40599 ( .B(n37603), .A(n37604), .Z(n37601) );
  AND U40600 ( .A(a[26]), .B(b[33]), .Z(n37600) );
  XOR U40601 ( .A(n37606), .B(n37607), .Z(n37257) );
  ANDN U40602 ( .B(n37608), .A(n37609), .Z(n37606) );
  AND U40603 ( .A(a[27]), .B(b[32]), .Z(n37605) );
  XOR U40604 ( .A(n37611), .B(n37612), .Z(n37262) );
  ANDN U40605 ( .B(n37613), .A(n37614), .Z(n37611) );
  AND U40606 ( .A(a[28]), .B(b[31]), .Z(n37610) );
  XOR U40607 ( .A(n37616), .B(n37617), .Z(n37267) );
  ANDN U40608 ( .B(n37618), .A(n37619), .Z(n37616) );
  AND U40609 ( .A(a[29]), .B(b[30]), .Z(n37615) );
  XOR U40610 ( .A(n37621), .B(n37622), .Z(n37272) );
  ANDN U40611 ( .B(n37623), .A(n37624), .Z(n37621) );
  AND U40612 ( .A(a[30]), .B(b[29]), .Z(n37620) );
  XOR U40613 ( .A(n37626), .B(n37627), .Z(n37277) );
  ANDN U40614 ( .B(n37628), .A(n37629), .Z(n37626) );
  AND U40615 ( .A(a[31]), .B(b[28]), .Z(n37625) );
  XOR U40616 ( .A(n37631), .B(n37632), .Z(n37282) );
  ANDN U40617 ( .B(n37633), .A(n37634), .Z(n37631) );
  AND U40618 ( .A(a[32]), .B(b[27]), .Z(n37630) );
  XOR U40619 ( .A(n37636), .B(n37637), .Z(n37287) );
  ANDN U40620 ( .B(n37638), .A(n37639), .Z(n37636) );
  AND U40621 ( .A(a[33]), .B(b[26]), .Z(n37635) );
  XOR U40622 ( .A(n37641), .B(n37642), .Z(n37292) );
  ANDN U40623 ( .B(n37643), .A(n37644), .Z(n37641) );
  AND U40624 ( .A(a[34]), .B(b[25]), .Z(n37640) );
  XOR U40625 ( .A(n37646), .B(n37647), .Z(n37297) );
  ANDN U40626 ( .B(n37648), .A(n37649), .Z(n37646) );
  AND U40627 ( .A(a[35]), .B(b[24]), .Z(n37645) );
  XOR U40628 ( .A(n37651), .B(n37652), .Z(n37302) );
  ANDN U40629 ( .B(n37653), .A(n37654), .Z(n37651) );
  AND U40630 ( .A(a[36]), .B(b[23]), .Z(n37650) );
  XOR U40631 ( .A(n37656), .B(n37657), .Z(n37307) );
  ANDN U40632 ( .B(n37658), .A(n37659), .Z(n37656) );
  AND U40633 ( .A(a[37]), .B(b[22]), .Z(n37655) );
  XOR U40634 ( .A(n37661), .B(n37662), .Z(n37312) );
  ANDN U40635 ( .B(n37663), .A(n37664), .Z(n37661) );
  AND U40636 ( .A(a[38]), .B(b[21]), .Z(n37660) );
  XOR U40637 ( .A(n37666), .B(n37667), .Z(n37317) );
  ANDN U40638 ( .B(n37668), .A(n37669), .Z(n37666) );
  AND U40639 ( .A(a[39]), .B(b[20]), .Z(n37665) );
  XOR U40640 ( .A(n37671), .B(n37672), .Z(n37322) );
  ANDN U40641 ( .B(n37673), .A(n37674), .Z(n37671) );
  AND U40642 ( .A(a[40]), .B(b[19]), .Z(n37670) );
  XOR U40643 ( .A(n37676), .B(n37677), .Z(n37327) );
  ANDN U40644 ( .B(n37678), .A(n37679), .Z(n37676) );
  AND U40645 ( .A(a[41]), .B(b[18]), .Z(n37675) );
  XOR U40646 ( .A(n37681), .B(n37682), .Z(n37332) );
  ANDN U40647 ( .B(n37683), .A(n37684), .Z(n37681) );
  AND U40648 ( .A(a[42]), .B(b[17]), .Z(n37680) );
  XOR U40649 ( .A(n37686), .B(n37687), .Z(n37337) );
  ANDN U40650 ( .B(n37688), .A(n37689), .Z(n37686) );
  AND U40651 ( .A(a[43]), .B(b[16]), .Z(n37685) );
  XOR U40652 ( .A(n37691), .B(n37692), .Z(n37342) );
  ANDN U40653 ( .B(n37693), .A(n37694), .Z(n37691) );
  AND U40654 ( .A(a[44]), .B(b[15]), .Z(n37690) );
  XOR U40655 ( .A(n37696), .B(n37697), .Z(n37347) );
  ANDN U40656 ( .B(n37698), .A(n37699), .Z(n37696) );
  AND U40657 ( .A(a[45]), .B(b[14]), .Z(n37695) );
  XOR U40658 ( .A(n37701), .B(n37702), .Z(n37352) );
  ANDN U40659 ( .B(n37703), .A(n37704), .Z(n37701) );
  AND U40660 ( .A(a[46]), .B(b[13]), .Z(n37700) );
  XOR U40661 ( .A(n37706), .B(n37707), .Z(n37357) );
  ANDN U40662 ( .B(n37708), .A(n37709), .Z(n37706) );
  AND U40663 ( .A(a[47]), .B(b[12]), .Z(n37705) );
  XOR U40664 ( .A(n37711), .B(n37712), .Z(n37362) );
  ANDN U40665 ( .B(n37713), .A(n37714), .Z(n37711) );
  AND U40666 ( .A(a[48]), .B(b[11]), .Z(n37710) );
  XOR U40667 ( .A(n37716), .B(n37717), .Z(n37367) );
  ANDN U40668 ( .B(n37718), .A(n37719), .Z(n37716) );
  AND U40669 ( .A(a[49]), .B(b[10]), .Z(n37715) );
  XOR U40670 ( .A(n37721), .B(n37722), .Z(n37372) );
  ANDN U40671 ( .B(n37723), .A(n37724), .Z(n37721) );
  AND U40672 ( .A(b[9]), .B(a[50]), .Z(n37720) );
  XOR U40673 ( .A(n37726), .B(n37727), .Z(n37377) );
  ANDN U40674 ( .B(n37728), .A(n37729), .Z(n37726) );
  AND U40675 ( .A(b[8]), .B(a[51]), .Z(n37725) );
  XOR U40676 ( .A(n37731), .B(n37732), .Z(n37382) );
  ANDN U40677 ( .B(n37733), .A(n37734), .Z(n37731) );
  AND U40678 ( .A(b[7]), .B(a[52]), .Z(n37730) );
  XOR U40679 ( .A(n37736), .B(n37737), .Z(n37387) );
  ANDN U40680 ( .B(n37738), .A(n37739), .Z(n37736) );
  AND U40681 ( .A(b[6]), .B(a[53]), .Z(n37735) );
  XOR U40682 ( .A(n37741), .B(n37742), .Z(n37392) );
  ANDN U40683 ( .B(n37743), .A(n37744), .Z(n37741) );
  AND U40684 ( .A(b[5]), .B(a[54]), .Z(n37740) );
  XOR U40685 ( .A(n37746), .B(n37747), .Z(n37397) );
  ANDN U40686 ( .B(n37748), .A(n37749), .Z(n37746) );
  AND U40687 ( .A(b[4]), .B(a[55]), .Z(n37745) );
  XOR U40688 ( .A(n37751), .B(n37752), .Z(n37402) );
  ANDN U40689 ( .B(n37414), .A(n37415), .Z(n37751) );
  AND U40690 ( .A(b[2]), .B(a[56]), .Z(n37753) );
  XNOR U40691 ( .A(n37748), .B(n37752), .Z(n37754) );
  XOR U40692 ( .A(n37755), .B(n37756), .Z(n37752) );
  OR U40693 ( .A(n37417), .B(n37418), .Z(n37756) );
  XNOR U40694 ( .A(n37758), .B(n37759), .Z(n37757) );
  XOR U40695 ( .A(n37758), .B(n37761), .Z(n37417) );
  NAND U40696 ( .A(b[1]), .B(a[56]), .Z(n37761) );
  IV U40697 ( .A(n37755), .Z(n37758) );
  NANDN U40698 ( .A(n97), .B(n98), .Z(n37755) );
  XOR U40699 ( .A(n37762), .B(n37763), .Z(n98) );
  NAND U40700 ( .A(a[56]), .B(b[0]), .Z(n97) );
  XNOR U40701 ( .A(n37743), .B(n37747), .Z(n37764) );
  XNOR U40702 ( .A(n37738), .B(n37742), .Z(n37765) );
  XNOR U40703 ( .A(n37733), .B(n37737), .Z(n37766) );
  XNOR U40704 ( .A(n37728), .B(n37732), .Z(n37767) );
  XNOR U40705 ( .A(n37723), .B(n37727), .Z(n37768) );
  XNOR U40706 ( .A(n37718), .B(n37722), .Z(n37769) );
  XNOR U40707 ( .A(n37713), .B(n37717), .Z(n37770) );
  XNOR U40708 ( .A(n37708), .B(n37712), .Z(n37771) );
  XNOR U40709 ( .A(n37703), .B(n37707), .Z(n37772) );
  XNOR U40710 ( .A(n37698), .B(n37702), .Z(n37773) );
  XNOR U40711 ( .A(n37693), .B(n37697), .Z(n37774) );
  XNOR U40712 ( .A(n37688), .B(n37692), .Z(n37775) );
  XNOR U40713 ( .A(n37683), .B(n37687), .Z(n37776) );
  XNOR U40714 ( .A(n37678), .B(n37682), .Z(n37777) );
  XNOR U40715 ( .A(n37673), .B(n37677), .Z(n37778) );
  XNOR U40716 ( .A(n37668), .B(n37672), .Z(n37779) );
  XNOR U40717 ( .A(n37663), .B(n37667), .Z(n37780) );
  XNOR U40718 ( .A(n37658), .B(n37662), .Z(n37781) );
  XNOR U40719 ( .A(n37653), .B(n37657), .Z(n37782) );
  XNOR U40720 ( .A(n37648), .B(n37652), .Z(n37783) );
  XNOR U40721 ( .A(n37643), .B(n37647), .Z(n37784) );
  XNOR U40722 ( .A(n37638), .B(n37642), .Z(n37785) );
  XNOR U40723 ( .A(n37633), .B(n37637), .Z(n37786) );
  XNOR U40724 ( .A(n37628), .B(n37632), .Z(n37787) );
  XNOR U40725 ( .A(n37623), .B(n37627), .Z(n37788) );
  XNOR U40726 ( .A(n37618), .B(n37622), .Z(n37789) );
  XNOR U40727 ( .A(n37613), .B(n37617), .Z(n37790) );
  XNOR U40728 ( .A(n37608), .B(n37612), .Z(n37791) );
  XNOR U40729 ( .A(n37603), .B(n37607), .Z(n37792) );
  XNOR U40730 ( .A(n37598), .B(n37602), .Z(n37793) );
  XNOR U40731 ( .A(n37593), .B(n37597), .Z(n37794) );
  XNOR U40732 ( .A(n37588), .B(n37592), .Z(n37795) );
  XNOR U40733 ( .A(n37583), .B(n37587), .Z(n37796) );
  XNOR U40734 ( .A(n37578), .B(n37582), .Z(n37797) );
  XNOR U40735 ( .A(n37573), .B(n37577), .Z(n37798) );
  XNOR U40736 ( .A(n37568), .B(n37572), .Z(n37799) );
  XNOR U40737 ( .A(n37563), .B(n37567), .Z(n37800) );
  XNOR U40738 ( .A(n37558), .B(n37562), .Z(n37801) );
  XNOR U40739 ( .A(n37553), .B(n37557), .Z(n37802) );
  XNOR U40740 ( .A(n37548), .B(n37552), .Z(n37803) );
  XNOR U40741 ( .A(n37543), .B(n37547), .Z(n37804) );
  XNOR U40742 ( .A(n37538), .B(n37542), .Z(n37805) );
  XNOR U40743 ( .A(n37533), .B(n37537), .Z(n37806) );
  XNOR U40744 ( .A(n37528), .B(n37532), .Z(n37807) );
  XNOR U40745 ( .A(n37523), .B(n37527), .Z(n37808) );
  XNOR U40746 ( .A(n37518), .B(n37522), .Z(n37809) );
  XNOR U40747 ( .A(n37513), .B(n37517), .Z(n37810) );
  XNOR U40748 ( .A(n37508), .B(n37512), .Z(n37811) );
  XNOR U40749 ( .A(n37503), .B(n37507), .Z(n37812) );
  XNOR U40750 ( .A(n37498), .B(n37502), .Z(n37813) );
  XNOR U40751 ( .A(n37493), .B(n37497), .Z(n37814) );
  XNOR U40752 ( .A(n37488), .B(n37492), .Z(n37815) );
  XNOR U40753 ( .A(n37483), .B(n37487), .Z(n37816) );
  XNOR U40754 ( .A(n37478), .B(n37482), .Z(n37817) );
  XOR U40755 ( .A(n37818), .B(n37477), .Z(n37478) );
  AND U40756 ( .A(a[0]), .B(b[58]), .Z(n37818) );
  XNOR U40757 ( .A(n37819), .B(n37477), .Z(n37479) );
  XNOR U40758 ( .A(n37820), .B(n37821), .Z(n37477) );
  ANDN U40759 ( .B(n37822), .A(n37823), .Z(n37820) );
  AND U40760 ( .A(a[1]), .B(b[57]), .Z(n37819) );
  XOR U40761 ( .A(n37825), .B(n37826), .Z(n37482) );
  ANDN U40762 ( .B(n37827), .A(n37828), .Z(n37825) );
  AND U40763 ( .A(a[2]), .B(b[56]), .Z(n37824) );
  XOR U40764 ( .A(n37830), .B(n37831), .Z(n37487) );
  ANDN U40765 ( .B(n37832), .A(n37833), .Z(n37830) );
  AND U40766 ( .A(a[3]), .B(b[55]), .Z(n37829) );
  XOR U40767 ( .A(n37835), .B(n37836), .Z(n37492) );
  ANDN U40768 ( .B(n37837), .A(n37838), .Z(n37835) );
  AND U40769 ( .A(a[4]), .B(b[54]), .Z(n37834) );
  XOR U40770 ( .A(n37840), .B(n37841), .Z(n37497) );
  ANDN U40771 ( .B(n37842), .A(n37843), .Z(n37840) );
  AND U40772 ( .A(a[5]), .B(b[53]), .Z(n37839) );
  XOR U40773 ( .A(n37845), .B(n37846), .Z(n37502) );
  ANDN U40774 ( .B(n37847), .A(n37848), .Z(n37845) );
  AND U40775 ( .A(a[6]), .B(b[52]), .Z(n37844) );
  XOR U40776 ( .A(n37850), .B(n37851), .Z(n37507) );
  ANDN U40777 ( .B(n37852), .A(n37853), .Z(n37850) );
  AND U40778 ( .A(a[7]), .B(b[51]), .Z(n37849) );
  XOR U40779 ( .A(n37855), .B(n37856), .Z(n37512) );
  ANDN U40780 ( .B(n37857), .A(n37858), .Z(n37855) );
  AND U40781 ( .A(a[8]), .B(b[50]), .Z(n37854) );
  XOR U40782 ( .A(n37860), .B(n37861), .Z(n37517) );
  ANDN U40783 ( .B(n37862), .A(n37863), .Z(n37860) );
  AND U40784 ( .A(a[9]), .B(b[49]), .Z(n37859) );
  XOR U40785 ( .A(n37865), .B(n37866), .Z(n37522) );
  ANDN U40786 ( .B(n37867), .A(n37868), .Z(n37865) );
  AND U40787 ( .A(a[10]), .B(b[48]), .Z(n37864) );
  XOR U40788 ( .A(n37870), .B(n37871), .Z(n37527) );
  ANDN U40789 ( .B(n37872), .A(n37873), .Z(n37870) );
  AND U40790 ( .A(a[11]), .B(b[47]), .Z(n37869) );
  XOR U40791 ( .A(n37875), .B(n37876), .Z(n37532) );
  ANDN U40792 ( .B(n37877), .A(n37878), .Z(n37875) );
  AND U40793 ( .A(a[12]), .B(b[46]), .Z(n37874) );
  XOR U40794 ( .A(n37880), .B(n37881), .Z(n37537) );
  ANDN U40795 ( .B(n37882), .A(n37883), .Z(n37880) );
  AND U40796 ( .A(a[13]), .B(b[45]), .Z(n37879) );
  XOR U40797 ( .A(n37885), .B(n37886), .Z(n37542) );
  ANDN U40798 ( .B(n37887), .A(n37888), .Z(n37885) );
  AND U40799 ( .A(a[14]), .B(b[44]), .Z(n37884) );
  XOR U40800 ( .A(n37890), .B(n37891), .Z(n37547) );
  ANDN U40801 ( .B(n37892), .A(n37893), .Z(n37890) );
  AND U40802 ( .A(a[15]), .B(b[43]), .Z(n37889) );
  XOR U40803 ( .A(n37895), .B(n37896), .Z(n37552) );
  ANDN U40804 ( .B(n37897), .A(n37898), .Z(n37895) );
  AND U40805 ( .A(a[16]), .B(b[42]), .Z(n37894) );
  XOR U40806 ( .A(n37900), .B(n37901), .Z(n37557) );
  ANDN U40807 ( .B(n37902), .A(n37903), .Z(n37900) );
  AND U40808 ( .A(a[17]), .B(b[41]), .Z(n37899) );
  XOR U40809 ( .A(n37905), .B(n37906), .Z(n37562) );
  ANDN U40810 ( .B(n37907), .A(n37908), .Z(n37905) );
  AND U40811 ( .A(a[18]), .B(b[40]), .Z(n37904) );
  XOR U40812 ( .A(n37910), .B(n37911), .Z(n37567) );
  ANDN U40813 ( .B(n37912), .A(n37913), .Z(n37910) );
  AND U40814 ( .A(a[19]), .B(b[39]), .Z(n37909) );
  XOR U40815 ( .A(n37915), .B(n37916), .Z(n37572) );
  ANDN U40816 ( .B(n37917), .A(n37918), .Z(n37915) );
  AND U40817 ( .A(a[20]), .B(b[38]), .Z(n37914) );
  XOR U40818 ( .A(n37920), .B(n37921), .Z(n37577) );
  ANDN U40819 ( .B(n37922), .A(n37923), .Z(n37920) );
  AND U40820 ( .A(a[21]), .B(b[37]), .Z(n37919) );
  XOR U40821 ( .A(n37925), .B(n37926), .Z(n37582) );
  ANDN U40822 ( .B(n37927), .A(n37928), .Z(n37925) );
  AND U40823 ( .A(a[22]), .B(b[36]), .Z(n37924) );
  XOR U40824 ( .A(n37930), .B(n37931), .Z(n37587) );
  ANDN U40825 ( .B(n37932), .A(n37933), .Z(n37930) );
  AND U40826 ( .A(a[23]), .B(b[35]), .Z(n37929) );
  XOR U40827 ( .A(n37935), .B(n37936), .Z(n37592) );
  ANDN U40828 ( .B(n37937), .A(n37938), .Z(n37935) );
  AND U40829 ( .A(a[24]), .B(b[34]), .Z(n37934) );
  XOR U40830 ( .A(n37940), .B(n37941), .Z(n37597) );
  ANDN U40831 ( .B(n37942), .A(n37943), .Z(n37940) );
  AND U40832 ( .A(a[25]), .B(b[33]), .Z(n37939) );
  XOR U40833 ( .A(n37945), .B(n37946), .Z(n37602) );
  ANDN U40834 ( .B(n37947), .A(n37948), .Z(n37945) );
  AND U40835 ( .A(a[26]), .B(b[32]), .Z(n37944) );
  XOR U40836 ( .A(n37950), .B(n37951), .Z(n37607) );
  ANDN U40837 ( .B(n37952), .A(n37953), .Z(n37950) );
  AND U40838 ( .A(a[27]), .B(b[31]), .Z(n37949) );
  XOR U40839 ( .A(n37955), .B(n37956), .Z(n37612) );
  ANDN U40840 ( .B(n37957), .A(n37958), .Z(n37955) );
  AND U40841 ( .A(a[28]), .B(b[30]), .Z(n37954) );
  XOR U40842 ( .A(n37960), .B(n37961), .Z(n37617) );
  ANDN U40843 ( .B(n37962), .A(n37963), .Z(n37960) );
  AND U40844 ( .A(a[29]), .B(b[29]), .Z(n37959) );
  XOR U40845 ( .A(n37965), .B(n37966), .Z(n37622) );
  ANDN U40846 ( .B(n37967), .A(n37968), .Z(n37965) );
  AND U40847 ( .A(a[30]), .B(b[28]), .Z(n37964) );
  XOR U40848 ( .A(n37970), .B(n37971), .Z(n37627) );
  ANDN U40849 ( .B(n37972), .A(n37973), .Z(n37970) );
  AND U40850 ( .A(a[31]), .B(b[27]), .Z(n37969) );
  XOR U40851 ( .A(n37975), .B(n37976), .Z(n37632) );
  ANDN U40852 ( .B(n37977), .A(n37978), .Z(n37975) );
  AND U40853 ( .A(a[32]), .B(b[26]), .Z(n37974) );
  XOR U40854 ( .A(n37980), .B(n37981), .Z(n37637) );
  ANDN U40855 ( .B(n37982), .A(n37983), .Z(n37980) );
  AND U40856 ( .A(a[33]), .B(b[25]), .Z(n37979) );
  XOR U40857 ( .A(n37985), .B(n37986), .Z(n37642) );
  ANDN U40858 ( .B(n37987), .A(n37988), .Z(n37985) );
  AND U40859 ( .A(a[34]), .B(b[24]), .Z(n37984) );
  XOR U40860 ( .A(n37990), .B(n37991), .Z(n37647) );
  ANDN U40861 ( .B(n37992), .A(n37993), .Z(n37990) );
  AND U40862 ( .A(a[35]), .B(b[23]), .Z(n37989) );
  XOR U40863 ( .A(n37995), .B(n37996), .Z(n37652) );
  ANDN U40864 ( .B(n37997), .A(n37998), .Z(n37995) );
  AND U40865 ( .A(a[36]), .B(b[22]), .Z(n37994) );
  XOR U40866 ( .A(n38000), .B(n38001), .Z(n37657) );
  ANDN U40867 ( .B(n38002), .A(n38003), .Z(n38000) );
  AND U40868 ( .A(a[37]), .B(b[21]), .Z(n37999) );
  XOR U40869 ( .A(n38005), .B(n38006), .Z(n37662) );
  ANDN U40870 ( .B(n38007), .A(n38008), .Z(n38005) );
  AND U40871 ( .A(a[38]), .B(b[20]), .Z(n38004) );
  XOR U40872 ( .A(n38010), .B(n38011), .Z(n37667) );
  ANDN U40873 ( .B(n38012), .A(n38013), .Z(n38010) );
  AND U40874 ( .A(a[39]), .B(b[19]), .Z(n38009) );
  XOR U40875 ( .A(n38015), .B(n38016), .Z(n37672) );
  ANDN U40876 ( .B(n38017), .A(n38018), .Z(n38015) );
  AND U40877 ( .A(a[40]), .B(b[18]), .Z(n38014) );
  XOR U40878 ( .A(n38020), .B(n38021), .Z(n37677) );
  ANDN U40879 ( .B(n38022), .A(n38023), .Z(n38020) );
  AND U40880 ( .A(a[41]), .B(b[17]), .Z(n38019) );
  XOR U40881 ( .A(n38025), .B(n38026), .Z(n37682) );
  ANDN U40882 ( .B(n38027), .A(n38028), .Z(n38025) );
  AND U40883 ( .A(a[42]), .B(b[16]), .Z(n38024) );
  XOR U40884 ( .A(n38030), .B(n38031), .Z(n37687) );
  ANDN U40885 ( .B(n38032), .A(n38033), .Z(n38030) );
  AND U40886 ( .A(a[43]), .B(b[15]), .Z(n38029) );
  XOR U40887 ( .A(n38035), .B(n38036), .Z(n37692) );
  ANDN U40888 ( .B(n38037), .A(n38038), .Z(n38035) );
  AND U40889 ( .A(a[44]), .B(b[14]), .Z(n38034) );
  XOR U40890 ( .A(n38040), .B(n38041), .Z(n37697) );
  ANDN U40891 ( .B(n38042), .A(n38043), .Z(n38040) );
  AND U40892 ( .A(a[45]), .B(b[13]), .Z(n38039) );
  XOR U40893 ( .A(n38045), .B(n38046), .Z(n37702) );
  ANDN U40894 ( .B(n38047), .A(n38048), .Z(n38045) );
  AND U40895 ( .A(a[46]), .B(b[12]), .Z(n38044) );
  XOR U40896 ( .A(n38050), .B(n38051), .Z(n37707) );
  ANDN U40897 ( .B(n38052), .A(n38053), .Z(n38050) );
  AND U40898 ( .A(a[47]), .B(b[11]), .Z(n38049) );
  XOR U40899 ( .A(n38055), .B(n38056), .Z(n37712) );
  ANDN U40900 ( .B(n38057), .A(n38058), .Z(n38055) );
  AND U40901 ( .A(a[48]), .B(b[10]), .Z(n38054) );
  XOR U40902 ( .A(n38060), .B(n38061), .Z(n37717) );
  ANDN U40903 ( .B(n38062), .A(n38063), .Z(n38060) );
  AND U40904 ( .A(b[9]), .B(a[49]), .Z(n38059) );
  XOR U40905 ( .A(n38065), .B(n38066), .Z(n37722) );
  ANDN U40906 ( .B(n38067), .A(n38068), .Z(n38065) );
  AND U40907 ( .A(b[8]), .B(a[50]), .Z(n38064) );
  XOR U40908 ( .A(n38070), .B(n38071), .Z(n37727) );
  ANDN U40909 ( .B(n38072), .A(n38073), .Z(n38070) );
  AND U40910 ( .A(b[7]), .B(a[51]), .Z(n38069) );
  XOR U40911 ( .A(n38075), .B(n38076), .Z(n37732) );
  ANDN U40912 ( .B(n38077), .A(n38078), .Z(n38075) );
  AND U40913 ( .A(b[6]), .B(a[52]), .Z(n38074) );
  XOR U40914 ( .A(n38080), .B(n38081), .Z(n37737) );
  ANDN U40915 ( .B(n38082), .A(n38083), .Z(n38080) );
  AND U40916 ( .A(b[5]), .B(a[53]), .Z(n38079) );
  XOR U40917 ( .A(n38085), .B(n38086), .Z(n37742) );
  ANDN U40918 ( .B(n38087), .A(n38088), .Z(n38085) );
  AND U40919 ( .A(b[4]), .B(a[54]), .Z(n38084) );
  XOR U40920 ( .A(n38090), .B(n38091), .Z(n37747) );
  ANDN U40921 ( .B(n37759), .A(n37760), .Z(n38090) );
  AND U40922 ( .A(b[2]), .B(a[55]), .Z(n38092) );
  XNOR U40923 ( .A(n38087), .B(n38091), .Z(n38093) );
  XOR U40924 ( .A(n38094), .B(n38095), .Z(n38091) );
  OR U40925 ( .A(n37762), .B(n37763), .Z(n38095) );
  XNOR U40926 ( .A(n38097), .B(n38098), .Z(n38096) );
  XOR U40927 ( .A(n38097), .B(n38100), .Z(n37762) );
  NAND U40928 ( .A(b[1]), .B(a[55]), .Z(n38100) );
  IV U40929 ( .A(n38094), .Z(n38097) );
  NANDN U40930 ( .A(n99), .B(n100), .Z(n38094) );
  XOR U40931 ( .A(n38101), .B(n38102), .Z(n100) );
  NAND U40932 ( .A(a[55]), .B(b[0]), .Z(n99) );
  XNOR U40933 ( .A(n38082), .B(n38086), .Z(n38103) );
  XNOR U40934 ( .A(n38077), .B(n38081), .Z(n38104) );
  XNOR U40935 ( .A(n38072), .B(n38076), .Z(n38105) );
  XNOR U40936 ( .A(n38067), .B(n38071), .Z(n38106) );
  XNOR U40937 ( .A(n38062), .B(n38066), .Z(n38107) );
  XNOR U40938 ( .A(n38057), .B(n38061), .Z(n38108) );
  XNOR U40939 ( .A(n38052), .B(n38056), .Z(n38109) );
  XNOR U40940 ( .A(n38047), .B(n38051), .Z(n38110) );
  XNOR U40941 ( .A(n38042), .B(n38046), .Z(n38111) );
  XNOR U40942 ( .A(n38037), .B(n38041), .Z(n38112) );
  XNOR U40943 ( .A(n38032), .B(n38036), .Z(n38113) );
  XNOR U40944 ( .A(n38027), .B(n38031), .Z(n38114) );
  XNOR U40945 ( .A(n38022), .B(n38026), .Z(n38115) );
  XNOR U40946 ( .A(n38017), .B(n38021), .Z(n38116) );
  XNOR U40947 ( .A(n38012), .B(n38016), .Z(n38117) );
  XNOR U40948 ( .A(n38007), .B(n38011), .Z(n38118) );
  XNOR U40949 ( .A(n38002), .B(n38006), .Z(n38119) );
  XNOR U40950 ( .A(n37997), .B(n38001), .Z(n38120) );
  XNOR U40951 ( .A(n37992), .B(n37996), .Z(n38121) );
  XNOR U40952 ( .A(n37987), .B(n37991), .Z(n38122) );
  XNOR U40953 ( .A(n37982), .B(n37986), .Z(n38123) );
  XNOR U40954 ( .A(n37977), .B(n37981), .Z(n38124) );
  XNOR U40955 ( .A(n37972), .B(n37976), .Z(n38125) );
  XNOR U40956 ( .A(n37967), .B(n37971), .Z(n38126) );
  XNOR U40957 ( .A(n37962), .B(n37966), .Z(n38127) );
  XNOR U40958 ( .A(n37957), .B(n37961), .Z(n38128) );
  XNOR U40959 ( .A(n37952), .B(n37956), .Z(n38129) );
  XNOR U40960 ( .A(n37947), .B(n37951), .Z(n38130) );
  XNOR U40961 ( .A(n37942), .B(n37946), .Z(n38131) );
  XNOR U40962 ( .A(n37937), .B(n37941), .Z(n38132) );
  XNOR U40963 ( .A(n37932), .B(n37936), .Z(n38133) );
  XNOR U40964 ( .A(n37927), .B(n37931), .Z(n38134) );
  XNOR U40965 ( .A(n37922), .B(n37926), .Z(n38135) );
  XNOR U40966 ( .A(n37917), .B(n37921), .Z(n38136) );
  XNOR U40967 ( .A(n37912), .B(n37916), .Z(n38137) );
  XNOR U40968 ( .A(n37907), .B(n37911), .Z(n38138) );
  XNOR U40969 ( .A(n37902), .B(n37906), .Z(n38139) );
  XNOR U40970 ( .A(n37897), .B(n37901), .Z(n38140) );
  XNOR U40971 ( .A(n37892), .B(n37896), .Z(n38141) );
  XNOR U40972 ( .A(n37887), .B(n37891), .Z(n38142) );
  XNOR U40973 ( .A(n37882), .B(n37886), .Z(n38143) );
  XNOR U40974 ( .A(n37877), .B(n37881), .Z(n38144) );
  XNOR U40975 ( .A(n37872), .B(n37876), .Z(n38145) );
  XNOR U40976 ( .A(n37867), .B(n37871), .Z(n38146) );
  XNOR U40977 ( .A(n37862), .B(n37866), .Z(n38147) );
  XNOR U40978 ( .A(n37857), .B(n37861), .Z(n38148) );
  XNOR U40979 ( .A(n37852), .B(n37856), .Z(n38149) );
  XNOR U40980 ( .A(n37847), .B(n37851), .Z(n38150) );
  XNOR U40981 ( .A(n37842), .B(n37846), .Z(n38151) );
  XNOR U40982 ( .A(n37837), .B(n37841), .Z(n38152) );
  XNOR U40983 ( .A(n37832), .B(n37836), .Z(n38153) );
  XNOR U40984 ( .A(n37827), .B(n37831), .Z(n38154) );
  XNOR U40985 ( .A(n37822), .B(n37826), .Z(n38155) );
  XNOR U40986 ( .A(n38156), .B(n37821), .Z(n37822) );
  AND U40987 ( .A(a[0]), .B(b[57]), .Z(n38156) );
  XOR U40988 ( .A(n38157), .B(n37821), .Z(n37823) );
  XNOR U40989 ( .A(n38158), .B(n38159), .Z(n37821) );
  ANDN U40990 ( .B(n38160), .A(n38161), .Z(n38158) );
  AND U40991 ( .A(a[1]), .B(b[56]), .Z(n38157) );
  XOR U40992 ( .A(n38163), .B(n38164), .Z(n37826) );
  ANDN U40993 ( .B(n38165), .A(n38166), .Z(n38163) );
  AND U40994 ( .A(a[2]), .B(b[55]), .Z(n38162) );
  XOR U40995 ( .A(n38168), .B(n38169), .Z(n37831) );
  ANDN U40996 ( .B(n38170), .A(n38171), .Z(n38168) );
  AND U40997 ( .A(a[3]), .B(b[54]), .Z(n38167) );
  XOR U40998 ( .A(n38173), .B(n38174), .Z(n37836) );
  ANDN U40999 ( .B(n38175), .A(n38176), .Z(n38173) );
  AND U41000 ( .A(a[4]), .B(b[53]), .Z(n38172) );
  XOR U41001 ( .A(n38178), .B(n38179), .Z(n37841) );
  ANDN U41002 ( .B(n38180), .A(n38181), .Z(n38178) );
  AND U41003 ( .A(a[5]), .B(b[52]), .Z(n38177) );
  XOR U41004 ( .A(n38183), .B(n38184), .Z(n37846) );
  ANDN U41005 ( .B(n38185), .A(n38186), .Z(n38183) );
  AND U41006 ( .A(a[6]), .B(b[51]), .Z(n38182) );
  XOR U41007 ( .A(n38188), .B(n38189), .Z(n37851) );
  ANDN U41008 ( .B(n38190), .A(n38191), .Z(n38188) );
  AND U41009 ( .A(a[7]), .B(b[50]), .Z(n38187) );
  XOR U41010 ( .A(n38193), .B(n38194), .Z(n37856) );
  ANDN U41011 ( .B(n38195), .A(n38196), .Z(n38193) );
  AND U41012 ( .A(a[8]), .B(b[49]), .Z(n38192) );
  XOR U41013 ( .A(n38198), .B(n38199), .Z(n37861) );
  ANDN U41014 ( .B(n38200), .A(n38201), .Z(n38198) );
  AND U41015 ( .A(a[9]), .B(b[48]), .Z(n38197) );
  XOR U41016 ( .A(n38203), .B(n38204), .Z(n37866) );
  ANDN U41017 ( .B(n38205), .A(n38206), .Z(n38203) );
  AND U41018 ( .A(a[10]), .B(b[47]), .Z(n38202) );
  XOR U41019 ( .A(n38208), .B(n38209), .Z(n37871) );
  ANDN U41020 ( .B(n38210), .A(n38211), .Z(n38208) );
  AND U41021 ( .A(a[11]), .B(b[46]), .Z(n38207) );
  XOR U41022 ( .A(n38213), .B(n38214), .Z(n37876) );
  ANDN U41023 ( .B(n38215), .A(n38216), .Z(n38213) );
  AND U41024 ( .A(a[12]), .B(b[45]), .Z(n38212) );
  XOR U41025 ( .A(n38218), .B(n38219), .Z(n37881) );
  ANDN U41026 ( .B(n38220), .A(n38221), .Z(n38218) );
  AND U41027 ( .A(a[13]), .B(b[44]), .Z(n38217) );
  XOR U41028 ( .A(n38223), .B(n38224), .Z(n37886) );
  ANDN U41029 ( .B(n38225), .A(n38226), .Z(n38223) );
  AND U41030 ( .A(a[14]), .B(b[43]), .Z(n38222) );
  XOR U41031 ( .A(n38228), .B(n38229), .Z(n37891) );
  ANDN U41032 ( .B(n38230), .A(n38231), .Z(n38228) );
  AND U41033 ( .A(a[15]), .B(b[42]), .Z(n38227) );
  XOR U41034 ( .A(n38233), .B(n38234), .Z(n37896) );
  ANDN U41035 ( .B(n38235), .A(n38236), .Z(n38233) );
  AND U41036 ( .A(a[16]), .B(b[41]), .Z(n38232) );
  XOR U41037 ( .A(n38238), .B(n38239), .Z(n37901) );
  ANDN U41038 ( .B(n38240), .A(n38241), .Z(n38238) );
  AND U41039 ( .A(a[17]), .B(b[40]), .Z(n38237) );
  XOR U41040 ( .A(n38243), .B(n38244), .Z(n37906) );
  ANDN U41041 ( .B(n38245), .A(n38246), .Z(n38243) );
  AND U41042 ( .A(a[18]), .B(b[39]), .Z(n38242) );
  XOR U41043 ( .A(n38248), .B(n38249), .Z(n37911) );
  ANDN U41044 ( .B(n38250), .A(n38251), .Z(n38248) );
  AND U41045 ( .A(a[19]), .B(b[38]), .Z(n38247) );
  XOR U41046 ( .A(n38253), .B(n38254), .Z(n37916) );
  ANDN U41047 ( .B(n38255), .A(n38256), .Z(n38253) );
  AND U41048 ( .A(a[20]), .B(b[37]), .Z(n38252) );
  XOR U41049 ( .A(n38258), .B(n38259), .Z(n37921) );
  ANDN U41050 ( .B(n38260), .A(n38261), .Z(n38258) );
  AND U41051 ( .A(a[21]), .B(b[36]), .Z(n38257) );
  XOR U41052 ( .A(n38263), .B(n38264), .Z(n37926) );
  ANDN U41053 ( .B(n38265), .A(n38266), .Z(n38263) );
  AND U41054 ( .A(a[22]), .B(b[35]), .Z(n38262) );
  XOR U41055 ( .A(n38268), .B(n38269), .Z(n37931) );
  ANDN U41056 ( .B(n38270), .A(n38271), .Z(n38268) );
  AND U41057 ( .A(a[23]), .B(b[34]), .Z(n38267) );
  XOR U41058 ( .A(n38273), .B(n38274), .Z(n37936) );
  ANDN U41059 ( .B(n38275), .A(n38276), .Z(n38273) );
  AND U41060 ( .A(a[24]), .B(b[33]), .Z(n38272) );
  XOR U41061 ( .A(n38278), .B(n38279), .Z(n37941) );
  ANDN U41062 ( .B(n38280), .A(n38281), .Z(n38278) );
  AND U41063 ( .A(a[25]), .B(b[32]), .Z(n38277) );
  XOR U41064 ( .A(n38283), .B(n38284), .Z(n37946) );
  ANDN U41065 ( .B(n38285), .A(n38286), .Z(n38283) );
  AND U41066 ( .A(a[26]), .B(b[31]), .Z(n38282) );
  XOR U41067 ( .A(n38288), .B(n38289), .Z(n37951) );
  ANDN U41068 ( .B(n38290), .A(n38291), .Z(n38288) );
  AND U41069 ( .A(a[27]), .B(b[30]), .Z(n38287) );
  XOR U41070 ( .A(n38293), .B(n38294), .Z(n37956) );
  ANDN U41071 ( .B(n38295), .A(n38296), .Z(n38293) );
  AND U41072 ( .A(a[28]), .B(b[29]), .Z(n38292) );
  XOR U41073 ( .A(n38298), .B(n38299), .Z(n37961) );
  ANDN U41074 ( .B(n38300), .A(n38301), .Z(n38298) );
  AND U41075 ( .A(a[29]), .B(b[28]), .Z(n38297) );
  XOR U41076 ( .A(n38303), .B(n38304), .Z(n37966) );
  ANDN U41077 ( .B(n38305), .A(n38306), .Z(n38303) );
  AND U41078 ( .A(a[30]), .B(b[27]), .Z(n38302) );
  XOR U41079 ( .A(n38308), .B(n38309), .Z(n37971) );
  ANDN U41080 ( .B(n38310), .A(n38311), .Z(n38308) );
  AND U41081 ( .A(a[31]), .B(b[26]), .Z(n38307) );
  XOR U41082 ( .A(n38313), .B(n38314), .Z(n37976) );
  ANDN U41083 ( .B(n38315), .A(n38316), .Z(n38313) );
  AND U41084 ( .A(a[32]), .B(b[25]), .Z(n38312) );
  XOR U41085 ( .A(n38318), .B(n38319), .Z(n37981) );
  ANDN U41086 ( .B(n38320), .A(n38321), .Z(n38318) );
  AND U41087 ( .A(a[33]), .B(b[24]), .Z(n38317) );
  XOR U41088 ( .A(n38323), .B(n38324), .Z(n37986) );
  ANDN U41089 ( .B(n38325), .A(n38326), .Z(n38323) );
  AND U41090 ( .A(a[34]), .B(b[23]), .Z(n38322) );
  XOR U41091 ( .A(n38328), .B(n38329), .Z(n37991) );
  ANDN U41092 ( .B(n38330), .A(n38331), .Z(n38328) );
  AND U41093 ( .A(a[35]), .B(b[22]), .Z(n38327) );
  XOR U41094 ( .A(n38333), .B(n38334), .Z(n37996) );
  ANDN U41095 ( .B(n38335), .A(n38336), .Z(n38333) );
  AND U41096 ( .A(a[36]), .B(b[21]), .Z(n38332) );
  XOR U41097 ( .A(n38338), .B(n38339), .Z(n38001) );
  ANDN U41098 ( .B(n38340), .A(n38341), .Z(n38338) );
  AND U41099 ( .A(a[37]), .B(b[20]), .Z(n38337) );
  XOR U41100 ( .A(n38343), .B(n38344), .Z(n38006) );
  ANDN U41101 ( .B(n38345), .A(n38346), .Z(n38343) );
  AND U41102 ( .A(a[38]), .B(b[19]), .Z(n38342) );
  XOR U41103 ( .A(n38348), .B(n38349), .Z(n38011) );
  ANDN U41104 ( .B(n38350), .A(n38351), .Z(n38348) );
  AND U41105 ( .A(a[39]), .B(b[18]), .Z(n38347) );
  XOR U41106 ( .A(n38353), .B(n38354), .Z(n38016) );
  ANDN U41107 ( .B(n38355), .A(n38356), .Z(n38353) );
  AND U41108 ( .A(a[40]), .B(b[17]), .Z(n38352) );
  XOR U41109 ( .A(n38358), .B(n38359), .Z(n38021) );
  ANDN U41110 ( .B(n38360), .A(n38361), .Z(n38358) );
  AND U41111 ( .A(a[41]), .B(b[16]), .Z(n38357) );
  XOR U41112 ( .A(n38363), .B(n38364), .Z(n38026) );
  ANDN U41113 ( .B(n38365), .A(n38366), .Z(n38363) );
  AND U41114 ( .A(a[42]), .B(b[15]), .Z(n38362) );
  XOR U41115 ( .A(n38368), .B(n38369), .Z(n38031) );
  ANDN U41116 ( .B(n38370), .A(n38371), .Z(n38368) );
  AND U41117 ( .A(a[43]), .B(b[14]), .Z(n38367) );
  XOR U41118 ( .A(n38373), .B(n38374), .Z(n38036) );
  ANDN U41119 ( .B(n38375), .A(n38376), .Z(n38373) );
  AND U41120 ( .A(a[44]), .B(b[13]), .Z(n38372) );
  XOR U41121 ( .A(n38378), .B(n38379), .Z(n38041) );
  ANDN U41122 ( .B(n38380), .A(n38381), .Z(n38378) );
  AND U41123 ( .A(a[45]), .B(b[12]), .Z(n38377) );
  XOR U41124 ( .A(n38383), .B(n38384), .Z(n38046) );
  ANDN U41125 ( .B(n38385), .A(n38386), .Z(n38383) );
  AND U41126 ( .A(a[46]), .B(b[11]), .Z(n38382) );
  XOR U41127 ( .A(n38388), .B(n38389), .Z(n38051) );
  ANDN U41128 ( .B(n38390), .A(n38391), .Z(n38388) );
  AND U41129 ( .A(a[47]), .B(b[10]), .Z(n38387) );
  XOR U41130 ( .A(n38393), .B(n38394), .Z(n38056) );
  ANDN U41131 ( .B(n38395), .A(n38396), .Z(n38393) );
  AND U41132 ( .A(b[9]), .B(a[48]), .Z(n38392) );
  XOR U41133 ( .A(n38398), .B(n38399), .Z(n38061) );
  ANDN U41134 ( .B(n38400), .A(n38401), .Z(n38398) );
  AND U41135 ( .A(b[8]), .B(a[49]), .Z(n38397) );
  XOR U41136 ( .A(n38403), .B(n38404), .Z(n38066) );
  ANDN U41137 ( .B(n38405), .A(n38406), .Z(n38403) );
  AND U41138 ( .A(b[7]), .B(a[50]), .Z(n38402) );
  XOR U41139 ( .A(n38408), .B(n38409), .Z(n38071) );
  ANDN U41140 ( .B(n38410), .A(n38411), .Z(n38408) );
  AND U41141 ( .A(b[6]), .B(a[51]), .Z(n38407) );
  XOR U41142 ( .A(n38413), .B(n38414), .Z(n38076) );
  ANDN U41143 ( .B(n38415), .A(n38416), .Z(n38413) );
  AND U41144 ( .A(b[5]), .B(a[52]), .Z(n38412) );
  XOR U41145 ( .A(n38418), .B(n38419), .Z(n38081) );
  ANDN U41146 ( .B(n38420), .A(n38421), .Z(n38418) );
  AND U41147 ( .A(b[4]), .B(a[53]), .Z(n38417) );
  XOR U41148 ( .A(n38423), .B(n38424), .Z(n38086) );
  ANDN U41149 ( .B(n38098), .A(n38099), .Z(n38423) );
  AND U41150 ( .A(b[2]), .B(a[54]), .Z(n38425) );
  XNOR U41151 ( .A(n38420), .B(n38424), .Z(n38426) );
  XOR U41152 ( .A(n38427), .B(n38428), .Z(n38424) );
  OR U41153 ( .A(n38101), .B(n38102), .Z(n38428) );
  XNOR U41154 ( .A(n38430), .B(n38431), .Z(n38429) );
  XOR U41155 ( .A(n38430), .B(n38433), .Z(n38101) );
  NAND U41156 ( .A(b[1]), .B(a[54]), .Z(n38433) );
  IV U41157 ( .A(n38427), .Z(n38430) );
  NANDN U41158 ( .A(n101), .B(n102), .Z(n38427) );
  XOR U41159 ( .A(n38434), .B(n38435), .Z(n102) );
  NAND U41160 ( .A(a[54]), .B(b[0]), .Z(n101) );
  XNOR U41161 ( .A(n38415), .B(n38419), .Z(n38436) );
  XNOR U41162 ( .A(n38410), .B(n38414), .Z(n38437) );
  XNOR U41163 ( .A(n38405), .B(n38409), .Z(n38438) );
  XNOR U41164 ( .A(n38400), .B(n38404), .Z(n38439) );
  XNOR U41165 ( .A(n38395), .B(n38399), .Z(n38440) );
  XNOR U41166 ( .A(n38390), .B(n38394), .Z(n38441) );
  XNOR U41167 ( .A(n38385), .B(n38389), .Z(n38442) );
  XNOR U41168 ( .A(n38380), .B(n38384), .Z(n38443) );
  XNOR U41169 ( .A(n38375), .B(n38379), .Z(n38444) );
  XNOR U41170 ( .A(n38370), .B(n38374), .Z(n38445) );
  XNOR U41171 ( .A(n38365), .B(n38369), .Z(n38446) );
  XNOR U41172 ( .A(n38360), .B(n38364), .Z(n38447) );
  XNOR U41173 ( .A(n38355), .B(n38359), .Z(n38448) );
  XNOR U41174 ( .A(n38350), .B(n38354), .Z(n38449) );
  XNOR U41175 ( .A(n38345), .B(n38349), .Z(n38450) );
  XNOR U41176 ( .A(n38340), .B(n38344), .Z(n38451) );
  XNOR U41177 ( .A(n38335), .B(n38339), .Z(n38452) );
  XNOR U41178 ( .A(n38330), .B(n38334), .Z(n38453) );
  XNOR U41179 ( .A(n38325), .B(n38329), .Z(n38454) );
  XNOR U41180 ( .A(n38320), .B(n38324), .Z(n38455) );
  XNOR U41181 ( .A(n38315), .B(n38319), .Z(n38456) );
  XNOR U41182 ( .A(n38310), .B(n38314), .Z(n38457) );
  XNOR U41183 ( .A(n38305), .B(n38309), .Z(n38458) );
  XNOR U41184 ( .A(n38300), .B(n38304), .Z(n38459) );
  XNOR U41185 ( .A(n38295), .B(n38299), .Z(n38460) );
  XNOR U41186 ( .A(n38290), .B(n38294), .Z(n38461) );
  XNOR U41187 ( .A(n38285), .B(n38289), .Z(n38462) );
  XNOR U41188 ( .A(n38280), .B(n38284), .Z(n38463) );
  XNOR U41189 ( .A(n38275), .B(n38279), .Z(n38464) );
  XNOR U41190 ( .A(n38270), .B(n38274), .Z(n38465) );
  XNOR U41191 ( .A(n38265), .B(n38269), .Z(n38466) );
  XNOR U41192 ( .A(n38260), .B(n38264), .Z(n38467) );
  XNOR U41193 ( .A(n38255), .B(n38259), .Z(n38468) );
  XNOR U41194 ( .A(n38250), .B(n38254), .Z(n38469) );
  XNOR U41195 ( .A(n38245), .B(n38249), .Z(n38470) );
  XNOR U41196 ( .A(n38240), .B(n38244), .Z(n38471) );
  XNOR U41197 ( .A(n38235), .B(n38239), .Z(n38472) );
  XNOR U41198 ( .A(n38230), .B(n38234), .Z(n38473) );
  XNOR U41199 ( .A(n38225), .B(n38229), .Z(n38474) );
  XNOR U41200 ( .A(n38220), .B(n38224), .Z(n38475) );
  XNOR U41201 ( .A(n38215), .B(n38219), .Z(n38476) );
  XNOR U41202 ( .A(n38210), .B(n38214), .Z(n38477) );
  XNOR U41203 ( .A(n38205), .B(n38209), .Z(n38478) );
  XNOR U41204 ( .A(n38200), .B(n38204), .Z(n38479) );
  XNOR U41205 ( .A(n38195), .B(n38199), .Z(n38480) );
  XNOR U41206 ( .A(n38190), .B(n38194), .Z(n38481) );
  XNOR U41207 ( .A(n38185), .B(n38189), .Z(n38482) );
  XNOR U41208 ( .A(n38180), .B(n38184), .Z(n38483) );
  XNOR U41209 ( .A(n38175), .B(n38179), .Z(n38484) );
  XNOR U41210 ( .A(n38170), .B(n38174), .Z(n38485) );
  XNOR U41211 ( .A(n38165), .B(n38169), .Z(n38486) );
  XNOR U41212 ( .A(n38160), .B(n38164), .Z(n38487) );
  XOR U41213 ( .A(n38488), .B(n38159), .Z(n38160) );
  AND U41214 ( .A(a[0]), .B(b[56]), .Z(n38488) );
  XNOR U41215 ( .A(n38489), .B(n38159), .Z(n38161) );
  XNOR U41216 ( .A(n38490), .B(n38491), .Z(n38159) );
  ANDN U41217 ( .B(n38492), .A(n38493), .Z(n38490) );
  AND U41218 ( .A(a[1]), .B(b[55]), .Z(n38489) );
  XOR U41219 ( .A(n38495), .B(n38496), .Z(n38164) );
  ANDN U41220 ( .B(n38497), .A(n38498), .Z(n38495) );
  AND U41221 ( .A(a[2]), .B(b[54]), .Z(n38494) );
  XOR U41222 ( .A(n38500), .B(n38501), .Z(n38169) );
  ANDN U41223 ( .B(n38502), .A(n38503), .Z(n38500) );
  AND U41224 ( .A(a[3]), .B(b[53]), .Z(n38499) );
  XOR U41225 ( .A(n38505), .B(n38506), .Z(n38174) );
  ANDN U41226 ( .B(n38507), .A(n38508), .Z(n38505) );
  AND U41227 ( .A(a[4]), .B(b[52]), .Z(n38504) );
  XOR U41228 ( .A(n38510), .B(n38511), .Z(n38179) );
  ANDN U41229 ( .B(n38512), .A(n38513), .Z(n38510) );
  AND U41230 ( .A(a[5]), .B(b[51]), .Z(n38509) );
  XOR U41231 ( .A(n38515), .B(n38516), .Z(n38184) );
  ANDN U41232 ( .B(n38517), .A(n38518), .Z(n38515) );
  AND U41233 ( .A(a[6]), .B(b[50]), .Z(n38514) );
  XOR U41234 ( .A(n38520), .B(n38521), .Z(n38189) );
  ANDN U41235 ( .B(n38522), .A(n38523), .Z(n38520) );
  AND U41236 ( .A(a[7]), .B(b[49]), .Z(n38519) );
  XOR U41237 ( .A(n38525), .B(n38526), .Z(n38194) );
  ANDN U41238 ( .B(n38527), .A(n38528), .Z(n38525) );
  AND U41239 ( .A(a[8]), .B(b[48]), .Z(n38524) );
  XOR U41240 ( .A(n38530), .B(n38531), .Z(n38199) );
  ANDN U41241 ( .B(n38532), .A(n38533), .Z(n38530) );
  AND U41242 ( .A(a[9]), .B(b[47]), .Z(n38529) );
  XOR U41243 ( .A(n38535), .B(n38536), .Z(n38204) );
  ANDN U41244 ( .B(n38537), .A(n38538), .Z(n38535) );
  AND U41245 ( .A(a[10]), .B(b[46]), .Z(n38534) );
  XOR U41246 ( .A(n38540), .B(n38541), .Z(n38209) );
  ANDN U41247 ( .B(n38542), .A(n38543), .Z(n38540) );
  AND U41248 ( .A(a[11]), .B(b[45]), .Z(n38539) );
  XOR U41249 ( .A(n38545), .B(n38546), .Z(n38214) );
  ANDN U41250 ( .B(n38547), .A(n38548), .Z(n38545) );
  AND U41251 ( .A(a[12]), .B(b[44]), .Z(n38544) );
  XOR U41252 ( .A(n38550), .B(n38551), .Z(n38219) );
  ANDN U41253 ( .B(n38552), .A(n38553), .Z(n38550) );
  AND U41254 ( .A(a[13]), .B(b[43]), .Z(n38549) );
  XOR U41255 ( .A(n38555), .B(n38556), .Z(n38224) );
  ANDN U41256 ( .B(n38557), .A(n38558), .Z(n38555) );
  AND U41257 ( .A(a[14]), .B(b[42]), .Z(n38554) );
  XOR U41258 ( .A(n38560), .B(n38561), .Z(n38229) );
  ANDN U41259 ( .B(n38562), .A(n38563), .Z(n38560) );
  AND U41260 ( .A(a[15]), .B(b[41]), .Z(n38559) );
  XOR U41261 ( .A(n38565), .B(n38566), .Z(n38234) );
  ANDN U41262 ( .B(n38567), .A(n38568), .Z(n38565) );
  AND U41263 ( .A(a[16]), .B(b[40]), .Z(n38564) );
  XOR U41264 ( .A(n38570), .B(n38571), .Z(n38239) );
  ANDN U41265 ( .B(n38572), .A(n38573), .Z(n38570) );
  AND U41266 ( .A(a[17]), .B(b[39]), .Z(n38569) );
  XOR U41267 ( .A(n38575), .B(n38576), .Z(n38244) );
  ANDN U41268 ( .B(n38577), .A(n38578), .Z(n38575) );
  AND U41269 ( .A(a[18]), .B(b[38]), .Z(n38574) );
  XOR U41270 ( .A(n38580), .B(n38581), .Z(n38249) );
  ANDN U41271 ( .B(n38582), .A(n38583), .Z(n38580) );
  AND U41272 ( .A(a[19]), .B(b[37]), .Z(n38579) );
  XOR U41273 ( .A(n38585), .B(n38586), .Z(n38254) );
  ANDN U41274 ( .B(n38587), .A(n38588), .Z(n38585) );
  AND U41275 ( .A(a[20]), .B(b[36]), .Z(n38584) );
  XOR U41276 ( .A(n38590), .B(n38591), .Z(n38259) );
  ANDN U41277 ( .B(n38592), .A(n38593), .Z(n38590) );
  AND U41278 ( .A(a[21]), .B(b[35]), .Z(n38589) );
  XOR U41279 ( .A(n38595), .B(n38596), .Z(n38264) );
  ANDN U41280 ( .B(n38597), .A(n38598), .Z(n38595) );
  AND U41281 ( .A(a[22]), .B(b[34]), .Z(n38594) );
  XOR U41282 ( .A(n38600), .B(n38601), .Z(n38269) );
  ANDN U41283 ( .B(n38602), .A(n38603), .Z(n38600) );
  AND U41284 ( .A(a[23]), .B(b[33]), .Z(n38599) );
  XOR U41285 ( .A(n38605), .B(n38606), .Z(n38274) );
  ANDN U41286 ( .B(n38607), .A(n38608), .Z(n38605) );
  AND U41287 ( .A(a[24]), .B(b[32]), .Z(n38604) );
  XOR U41288 ( .A(n38610), .B(n38611), .Z(n38279) );
  ANDN U41289 ( .B(n38612), .A(n38613), .Z(n38610) );
  AND U41290 ( .A(a[25]), .B(b[31]), .Z(n38609) );
  XOR U41291 ( .A(n38615), .B(n38616), .Z(n38284) );
  ANDN U41292 ( .B(n38617), .A(n38618), .Z(n38615) );
  AND U41293 ( .A(a[26]), .B(b[30]), .Z(n38614) );
  XOR U41294 ( .A(n38620), .B(n38621), .Z(n38289) );
  ANDN U41295 ( .B(n38622), .A(n38623), .Z(n38620) );
  AND U41296 ( .A(a[27]), .B(b[29]), .Z(n38619) );
  XOR U41297 ( .A(n38625), .B(n38626), .Z(n38294) );
  ANDN U41298 ( .B(n38627), .A(n38628), .Z(n38625) );
  AND U41299 ( .A(a[28]), .B(b[28]), .Z(n38624) );
  XOR U41300 ( .A(n38630), .B(n38631), .Z(n38299) );
  ANDN U41301 ( .B(n38632), .A(n38633), .Z(n38630) );
  AND U41302 ( .A(a[29]), .B(b[27]), .Z(n38629) );
  XOR U41303 ( .A(n38635), .B(n38636), .Z(n38304) );
  ANDN U41304 ( .B(n38637), .A(n38638), .Z(n38635) );
  AND U41305 ( .A(a[30]), .B(b[26]), .Z(n38634) );
  XOR U41306 ( .A(n38640), .B(n38641), .Z(n38309) );
  ANDN U41307 ( .B(n38642), .A(n38643), .Z(n38640) );
  AND U41308 ( .A(a[31]), .B(b[25]), .Z(n38639) );
  XOR U41309 ( .A(n38645), .B(n38646), .Z(n38314) );
  ANDN U41310 ( .B(n38647), .A(n38648), .Z(n38645) );
  AND U41311 ( .A(a[32]), .B(b[24]), .Z(n38644) );
  XOR U41312 ( .A(n38650), .B(n38651), .Z(n38319) );
  ANDN U41313 ( .B(n38652), .A(n38653), .Z(n38650) );
  AND U41314 ( .A(a[33]), .B(b[23]), .Z(n38649) );
  XOR U41315 ( .A(n38655), .B(n38656), .Z(n38324) );
  ANDN U41316 ( .B(n38657), .A(n38658), .Z(n38655) );
  AND U41317 ( .A(a[34]), .B(b[22]), .Z(n38654) );
  XOR U41318 ( .A(n38660), .B(n38661), .Z(n38329) );
  ANDN U41319 ( .B(n38662), .A(n38663), .Z(n38660) );
  AND U41320 ( .A(a[35]), .B(b[21]), .Z(n38659) );
  XOR U41321 ( .A(n38665), .B(n38666), .Z(n38334) );
  ANDN U41322 ( .B(n38667), .A(n38668), .Z(n38665) );
  AND U41323 ( .A(a[36]), .B(b[20]), .Z(n38664) );
  XOR U41324 ( .A(n38670), .B(n38671), .Z(n38339) );
  ANDN U41325 ( .B(n38672), .A(n38673), .Z(n38670) );
  AND U41326 ( .A(a[37]), .B(b[19]), .Z(n38669) );
  XOR U41327 ( .A(n38675), .B(n38676), .Z(n38344) );
  ANDN U41328 ( .B(n38677), .A(n38678), .Z(n38675) );
  AND U41329 ( .A(a[38]), .B(b[18]), .Z(n38674) );
  XOR U41330 ( .A(n38680), .B(n38681), .Z(n38349) );
  ANDN U41331 ( .B(n38682), .A(n38683), .Z(n38680) );
  AND U41332 ( .A(a[39]), .B(b[17]), .Z(n38679) );
  XOR U41333 ( .A(n38685), .B(n38686), .Z(n38354) );
  ANDN U41334 ( .B(n38687), .A(n38688), .Z(n38685) );
  AND U41335 ( .A(a[40]), .B(b[16]), .Z(n38684) );
  XOR U41336 ( .A(n38690), .B(n38691), .Z(n38359) );
  ANDN U41337 ( .B(n38692), .A(n38693), .Z(n38690) );
  AND U41338 ( .A(a[41]), .B(b[15]), .Z(n38689) );
  XOR U41339 ( .A(n38695), .B(n38696), .Z(n38364) );
  ANDN U41340 ( .B(n38697), .A(n38698), .Z(n38695) );
  AND U41341 ( .A(a[42]), .B(b[14]), .Z(n38694) );
  XOR U41342 ( .A(n38700), .B(n38701), .Z(n38369) );
  ANDN U41343 ( .B(n38702), .A(n38703), .Z(n38700) );
  AND U41344 ( .A(a[43]), .B(b[13]), .Z(n38699) );
  XOR U41345 ( .A(n38705), .B(n38706), .Z(n38374) );
  ANDN U41346 ( .B(n38707), .A(n38708), .Z(n38705) );
  AND U41347 ( .A(a[44]), .B(b[12]), .Z(n38704) );
  XOR U41348 ( .A(n38710), .B(n38711), .Z(n38379) );
  ANDN U41349 ( .B(n38712), .A(n38713), .Z(n38710) );
  AND U41350 ( .A(a[45]), .B(b[11]), .Z(n38709) );
  XOR U41351 ( .A(n38715), .B(n38716), .Z(n38384) );
  ANDN U41352 ( .B(n38717), .A(n38718), .Z(n38715) );
  AND U41353 ( .A(a[46]), .B(b[10]), .Z(n38714) );
  XOR U41354 ( .A(n38720), .B(n38721), .Z(n38389) );
  ANDN U41355 ( .B(n38722), .A(n38723), .Z(n38720) );
  AND U41356 ( .A(b[9]), .B(a[47]), .Z(n38719) );
  XOR U41357 ( .A(n38725), .B(n38726), .Z(n38394) );
  ANDN U41358 ( .B(n38727), .A(n38728), .Z(n38725) );
  AND U41359 ( .A(b[8]), .B(a[48]), .Z(n38724) );
  XOR U41360 ( .A(n38730), .B(n38731), .Z(n38399) );
  ANDN U41361 ( .B(n38732), .A(n38733), .Z(n38730) );
  AND U41362 ( .A(b[7]), .B(a[49]), .Z(n38729) );
  XOR U41363 ( .A(n38735), .B(n38736), .Z(n38404) );
  ANDN U41364 ( .B(n38737), .A(n38738), .Z(n38735) );
  AND U41365 ( .A(b[6]), .B(a[50]), .Z(n38734) );
  XOR U41366 ( .A(n38740), .B(n38741), .Z(n38409) );
  ANDN U41367 ( .B(n38742), .A(n38743), .Z(n38740) );
  AND U41368 ( .A(b[5]), .B(a[51]), .Z(n38739) );
  XOR U41369 ( .A(n38745), .B(n38746), .Z(n38414) );
  ANDN U41370 ( .B(n38747), .A(n38748), .Z(n38745) );
  AND U41371 ( .A(b[4]), .B(a[52]), .Z(n38744) );
  XOR U41372 ( .A(n38750), .B(n38751), .Z(n38419) );
  ANDN U41373 ( .B(n38431), .A(n38432), .Z(n38750) );
  AND U41374 ( .A(b[2]), .B(a[53]), .Z(n38752) );
  XNOR U41375 ( .A(n38747), .B(n38751), .Z(n38753) );
  XOR U41376 ( .A(n38754), .B(n38755), .Z(n38751) );
  OR U41377 ( .A(n38434), .B(n38435), .Z(n38755) );
  XNOR U41378 ( .A(n38757), .B(n38758), .Z(n38756) );
  XOR U41379 ( .A(n38757), .B(n38760), .Z(n38434) );
  NAND U41380 ( .A(b[1]), .B(a[53]), .Z(n38760) );
  IV U41381 ( .A(n38754), .Z(n38757) );
  NANDN U41382 ( .A(n103), .B(n104), .Z(n38754) );
  XOR U41383 ( .A(n38761), .B(n38762), .Z(n104) );
  NAND U41384 ( .A(a[53]), .B(b[0]), .Z(n103) );
  XNOR U41385 ( .A(n38742), .B(n38746), .Z(n38763) );
  XNOR U41386 ( .A(n38737), .B(n38741), .Z(n38764) );
  XNOR U41387 ( .A(n38732), .B(n38736), .Z(n38765) );
  XNOR U41388 ( .A(n38727), .B(n38731), .Z(n38766) );
  XNOR U41389 ( .A(n38722), .B(n38726), .Z(n38767) );
  XNOR U41390 ( .A(n38717), .B(n38721), .Z(n38768) );
  XNOR U41391 ( .A(n38712), .B(n38716), .Z(n38769) );
  XNOR U41392 ( .A(n38707), .B(n38711), .Z(n38770) );
  XNOR U41393 ( .A(n38702), .B(n38706), .Z(n38771) );
  XNOR U41394 ( .A(n38697), .B(n38701), .Z(n38772) );
  XNOR U41395 ( .A(n38692), .B(n38696), .Z(n38773) );
  XNOR U41396 ( .A(n38687), .B(n38691), .Z(n38774) );
  XNOR U41397 ( .A(n38682), .B(n38686), .Z(n38775) );
  XNOR U41398 ( .A(n38677), .B(n38681), .Z(n38776) );
  XNOR U41399 ( .A(n38672), .B(n38676), .Z(n38777) );
  XNOR U41400 ( .A(n38667), .B(n38671), .Z(n38778) );
  XNOR U41401 ( .A(n38662), .B(n38666), .Z(n38779) );
  XNOR U41402 ( .A(n38657), .B(n38661), .Z(n38780) );
  XNOR U41403 ( .A(n38652), .B(n38656), .Z(n38781) );
  XNOR U41404 ( .A(n38647), .B(n38651), .Z(n38782) );
  XNOR U41405 ( .A(n38642), .B(n38646), .Z(n38783) );
  XNOR U41406 ( .A(n38637), .B(n38641), .Z(n38784) );
  XNOR U41407 ( .A(n38632), .B(n38636), .Z(n38785) );
  XNOR U41408 ( .A(n38627), .B(n38631), .Z(n38786) );
  XNOR U41409 ( .A(n38622), .B(n38626), .Z(n38787) );
  XNOR U41410 ( .A(n38617), .B(n38621), .Z(n38788) );
  XNOR U41411 ( .A(n38612), .B(n38616), .Z(n38789) );
  XNOR U41412 ( .A(n38607), .B(n38611), .Z(n38790) );
  XNOR U41413 ( .A(n38602), .B(n38606), .Z(n38791) );
  XNOR U41414 ( .A(n38597), .B(n38601), .Z(n38792) );
  XNOR U41415 ( .A(n38592), .B(n38596), .Z(n38793) );
  XNOR U41416 ( .A(n38587), .B(n38591), .Z(n38794) );
  XNOR U41417 ( .A(n38582), .B(n38586), .Z(n38795) );
  XNOR U41418 ( .A(n38577), .B(n38581), .Z(n38796) );
  XNOR U41419 ( .A(n38572), .B(n38576), .Z(n38797) );
  XNOR U41420 ( .A(n38567), .B(n38571), .Z(n38798) );
  XNOR U41421 ( .A(n38562), .B(n38566), .Z(n38799) );
  XNOR U41422 ( .A(n38557), .B(n38561), .Z(n38800) );
  XNOR U41423 ( .A(n38552), .B(n38556), .Z(n38801) );
  XNOR U41424 ( .A(n38547), .B(n38551), .Z(n38802) );
  XNOR U41425 ( .A(n38542), .B(n38546), .Z(n38803) );
  XNOR U41426 ( .A(n38537), .B(n38541), .Z(n38804) );
  XNOR U41427 ( .A(n38532), .B(n38536), .Z(n38805) );
  XNOR U41428 ( .A(n38527), .B(n38531), .Z(n38806) );
  XNOR U41429 ( .A(n38522), .B(n38526), .Z(n38807) );
  XNOR U41430 ( .A(n38517), .B(n38521), .Z(n38808) );
  XNOR U41431 ( .A(n38512), .B(n38516), .Z(n38809) );
  XNOR U41432 ( .A(n38507), .B(n38511), .Z(n38810) );
  XNOR U41433 ( .A(n38502), .B(n38506), .Z(n38811) );
  XNOR U41434 ( .A(n38497), .B(n38501), .Z(n38812) );
  XNOR U41435 ( .A(n38492), .B(n38496), .Z(n38813) );
  XNOR U41436 ( .A(n38814), .B(n38491), .Z(n38492) );
  AND U41437 ( .A(a[0]), .B(b[55]), .Z(n38814) );
  XOR U41438 ( .A(n38815), .B(n38491), .Z(n38493) );
  XNOR U41439 ( .A(n38816), .B(n38817), .Z(n38491) );
  ANDN U41440 ( .B(n38818), .A(n38819), .Z(n38816) );
  AND U41441 ( .A(a[1]), .B(b[54]), .Z(n38815) );
  XOR U41442 ( .A(n38821), .B(n38822), .Z(n38496) );
  ANDN U41443 ( .B(n38823), .A(n38824), .Z(n38821) );
  AND U41444 ( .A(a[2]), .B(b[53]), .Z(n38820) );
  XOR U41445 ( .A(n38826), .B(n38827), .Z(n38501) );
  ANDN U41446 ( .B(n38828), .A(n38829), .Z(n38826) );
  AND U41447 ( .A(a[3]), .B(b[52]), .Z(n38825) );
  XOR U41448 ( .A(n38831), .B(n38832), .Z(n38506) );
  ANDN U41449 ( .B(n38833), .A(n38834), .Z(n38831) );
  AND U41450 ( .A(a[4]), .B(b[51]), .Z(n38830) );
  XOR U41451 ( .A(n38836), .B(n38837), .Z(n38511) );
  ANDN U41452 ( .B(n38838), .A(n38839), .Z(n38836) );
  AND U41453 ( .A(a[5]), .B(b[50]), .Z(n38835) );
  XOR U41454 ( .A(n38841), .B(n38842), .Z(n38516) );
  ANDN U41455 ( .B(n38843), .A(n38844), .Z(n38841) );
  AND U41456 ( .A(a[6]), .B(b[49]), .Z(n38840) );
  XOR U41457 ( .A(n38846), .B(n38847), .Z(n38521) );
  ANDN U41458 ( .B(n38848), .A(n38849), .Z(n38846) );
  AND U41459 ( .A(a[7]), .B(b[48]), .Z(n38845) );
  XOR U41460 ( .A(n38851), .B(n38852), .Z(n38526) );
  ANDN U41461 ( .B(n38853), .A(n38854), .Z(n38851) );
  AND U41462 ( .A(a[8]), .B(b[47]), .Z(n38850) );
  XOR U41463 ( .A(n38856), .B(n38857), .Z(n38531) );
  ANDN U41464 ( .B(n38858), .A(n38859), .Z(n38856) );
  AND U41465 ( .A(a[9]), .B(b[46]), .Z(n38855) );
  XOR U41466 ( .A(n38861), .B(n38862), .Z(n38536) );
  ANDN U41467 ( .B(n38863), .A(n38864), .Z(n38861) );
  AND U41468 ( .A(a[10]), .B(b[45]), .Z(n38860) );
  XOR U41469 ( .A(n38866), .B(n38867), .Z(n38541) );
  ANDN U41470 ( .B(n38868), .A(n38869), .Z(n38866) );
  AND U41471 ( .A(a[11]), .B(b[44]), .Z(n38865) );
  XOR U41472 ( .A(n38871), .B(n38872), .Z(n38546) );
  ANDN U41473 ( .B(n38873), .A(n38874), .Z(n38871) );
  AND U41474 ( .A(a[12]), .B(b[43]), .Z(n38870) );
  XOR U41475 ( .A(n38876), .B(n38877), .Z(n38551) );
  ANDN U41476 ( .B(n38878), .A(n38879), .Z(n38876) );
  AND U41477 ( .A(a[13]), .B(b[42]), .Z(n38875) );
  XOR U41478 ( .A(n38881), .B(n38882), .Z(n38556) );
  ANDN U41479 ( .B(n38883), .A(n38884), .Z(n38881) );
  AND U41480 ( .A(a[14]), .B(b[41]), .Z(n38880) );
  XOR U41481 ( .A(n38886), .B(n38887), .Z(n38561) );
  ANDN U41482 ( .B(n38888), .A(n38889), .Z(n38886) );
  AND U41483 ( .A(a[15]), .B(b[40]), .Z(n38885) );
  XOR U41484 ( .A(n38891), .B(n38892), .Z(n38566) );
  ANDN U41485 ( .B(n38893), .A(n38894), .Z(n38891) );
  AND U41486 ( .A(a[16]), .B(b[39]), .Z(n38890) );
  XOR U41487 ( .A(n38896), .B(n38897), .Z(n38571) );
  ANDN U41488 ( .B(n38898), .A(n38899), .Z(n38896) );
  AND U41489 ( .A(a[17]), .B(b[38]), .Z(n38895) );
  XOR U41490 ( .A(n38901), .B(n38902), .Z(n38576) );
  ANDN U41491 ( .B(n38903), .A(n38904), .Z(n38901) );
  AND U41492 ( .A(a[18]), .B(b[37]), .Z(n38900) );
  XOR U41493 ( .A(n38906), .B(n38907), .Z(n38581) );
  ANDN U41494 ( .B(n38908), .A(n38909), .Z(n38906) );
  AND U41495 ( .A(a[19]), .B(b[36]), .Z(n38905) );
  XOR U41496 ( .A(n38911), .B(n38912), .Z(n38586) );
  ANDN U41497 ( .B(n38913), .A(n38914), .Z(n38911) );
  AND U41498 ( .A(a[20]), .B(b[35]), .Z(n38910) );
  XOR U41499 ( .A(n38916), .B(n38917), .Z(n38591) );
  ANDN U41500 ( .B(n38918), .A(n38919), .Z(n38916) );
  AND U41501 ( .A(a[21]), .B(b[34]), .Z(n38915) );
  XOR U41502 ( .A(n38921), .B(n38922), .Z(n38596) );
  ANDN U41503 ( .B(n38923), .A(n38924), .Z(n38921) );
  AND U41504 ( .A(a[22]), .B(b[33]), .Z(n38920) );
  XOR U41505 ( .A(n38926), .B(n38927), .Z(n38601) );
  ANDN U41506 ( .B(n38928), .A(n38929), .Z(n38926) );
  AND U41507 ( .A(a[23]), .B(b[32]), .Z(n38925) );
  XOR U41508 ( .A(n38931), .B(n38932), .Z(n38606) );
  ANDN U41509 ( .B(n38933), .A(n38934), .Z(n38931) );
  AND U41510 ( .A(a[24]), .B(b[31]), .Z(n38930) );
  XOR U41511 ( .A(n38936), .B(n38937), .Z(n38611) );
  ANDN U41512 ( .B(n38938), .A(n38939), .Z(n38936) );
  AND U41513 ( .A(a[25]), .B(b[30]), .Z(n38935) );
  XOR U41514 ( .A(n38941), .B(n38942), .Z(n38616) );
  ANDN U41515 ( .B(n38943), .A(n38944), .Z(n38941) );
  AND U41516 ( .A(a[26]), .B(b[29]), .Z(n38940) );
  XOR U41517 ( .A(n38946), .B(n38947), .Z(n38621) );
  ANDN U41518 ( .B(n38948), .A(n38949), .Z(n38946) );
  AND U41519 ( .A(a[27]), .B(b[28]), .Z(n38945) );
  XOR U41520 ( .A(n38951), .B(n38952), .Z(n38626) );
  ANDN U41521 ( .B(n38953), .A(n38954), .Z(n38951) );
  AND U41522 ( .A(a[28]), .B(b[27]), .Z(n38950) );
  XOR U41523 ( .A(n38956), .B(n38957), .Z(n38631) );
  ANDN U41524 ( .B(n38958), .A(n38959), .Z(n38956) );
  AND U41525 ( .A(a[29]), .B(b[26]), .Z(n38955) );
  XOR U41526 ( .A(n38961), .B(n38962), .Z(n38636) );
  ANDN U41527 ( .B(n38963), .A(n38964), .Z(n38961) );
  AND U41528 ( .A(a[30]), .B(b[25]), .Z(n38960) );
  XOR U41529 ( .A(n38966), .B(n38967), .Z(n38641) );
  ANDN U41530 ( .B(n38968), .A(n38969), .Z(n38966) );
  AND U41531 ( .A(a[31]), .B(b[24]), .Z(n38965) );
  XOR U41532 ( .A(n38971), .B(n38972), .Z(n38646) );
  ANDN U41533 ( .B(n38973), .A(n38974), .Z(n38971) );
  AND U41534 ( .A(a[32]), .B(b[23]), .Z(n38970) );
  XOR U41535 ( .A(n38976), .B(n38977), .Z(n38651) );
  ANDN U41536 ( .B(n38978), .A(n38979), .Z(n38976) );
  AND U41537 ( .A(a[33]), .B(b[22]), .Z(n38975) );
  XOR U41538 ( .A(n38981), .B(n38982), .Z(n38656) );
  ANDN U41539 ( .B(n38983), .A(n38984), .Z(n38981) );
  AND U41540 ( .A(a[34]), .B(b[21]), .Z(n38980) );
  XOR U41541 ( .A(n38986), .B(n38987), .Z(n38661) );
  ANDN U41542 ( .B(n38988), .A(n38989), .Z(n38986) );
  AND U41543 ( .A(a[35]), .B(b[20]), .Z(n38985) );
  XOR U41544 ( .A(n38991), .B(n38992), .Z(n38666) );
  ANDN U41545 ( .B(n38993), .A(n38994), .Z(n38991) );
  AND U41546 ( .A(a[36]), .B(b[19]), .Z(n38990) );
  XOR U41547 ( .A(n38996), .B(n38997), .Z(n38671) );
  ANDN U41548 ( .B(n38998), .A(n38999), .Z(n38996) );
  AND U41549 ( .A(a[37]), .B(b[18]), .Z(n38995) );
  XOR U41550 ( .A(n39001), .B(n39002), .Z(n38676) );
  ANDN U41551 ( .B(n39003), .A(n39004), .Z(n39001) );
  AND U41552 ( .A(a[38]), .B(b[17]), .Z(n39000) );
  XOR U41553 ( .A(n39006), .B(n39007), .Z(n38681) );
  ANDN U41554 ( .B(n39008), .A(n39009), .Z(n39006) );
  AND U41555 ( .A(a[39]), .B(b[16]), .Z(n39005) );
  XOR U41556 ( .A(n39011), .B(n39012), .Z(n38686) );
  ANDN U41557 ( .B(n39013), .A(n39014), .Z(n39011) );
  AND U41558 ( .A(a[40]), .B(b[15]), .Z(n39010) );
  XOR U41559 ( .A(n39016), .B(n39017), .Z(n38691) );
  ANDN U41560 ( .B(n39018), .A(n39019), .Z(n39016) );
  AND U41561 ( .A(a[41]), .B(b[14]), .Z(n39015) );
  XOR U41562 ( .A(n39021), .B(n39022), .Z(n38696) );
  ANDN U41563 ( .B(n39023), .A(n39024), .Z(n39021) );
  AND U41564 ( .A(a[42]), .B(b[13]), .Z(n39020) );
  XOR U41565 ( .A(n39026), .B(n39027), .Z(n38701) );
  ANDN U41566 ( .B(n39028), .A(n39029), .Z(n39026) );
  AND U41567 ( .A(a[43]), .B(b[12]), .Z(n39025) );
  XOR U41568 ( .A(n39031), .B(n39032), .Z(n38706) );
  ANDN U41569 ( .B(n39033), .A(n39034), .Z(n39031) );
  AND U41570 ( .A(a[44]), .B(b[11]), .Z(n39030) );
  XOR U41571 ( .A(n39036), .B(n39037), .Z(n38711) );
  ANDN U41572 ( .B(n39038), .A(n39039), .Z(n39036) );
  AND U41573 ( .A(a[45]), .B(b[10]), .Z(n39035) );
  XOR U41574 ( .A(n39041), .B(n39042), .Z(n38716) );
  ANDN U41575 ( .B(n39043), .A(n39044), .Z(n39041) );
  AND U41576 ( .A(b[9]), .B(a[46]), .Z(n39040) );
  XOR U41577 ( .A(n39046), .B(n39047), .Z(n38721) );
  ANDN U41578 ( .B(n39048), .A(n39049), .Z(n39046) );
  AND U41579 ( .A(b[8]), .B(a[47]), .Z(n39045) );
  XOR U41580 ( .A(n39051), .B(n39052), .Z(n38726) );
  ANDN U41581 ( .B(n39053), .A(n39054), .Z(n39051) );
  AND U41582 ( .A(b[7]), .B(a[48]), .Z(n39050) );
  XOR U41583 ( .A(n39056), .B(n39057), .Z(n38731) );
  ANDN U41584 ( .B(n39058), .A(n39059), .Z(n39056) );
  AND U41585 ( .A(b[6]), .B(a[49]), .Z(n39055) );
  XOR U41586 ( .A(n39061), .B(n39062), .Z(n38736) );
  ANDN U41587 ( .B(n39063), .A(n39064), .Z(n39061) );
  AND U41588 ( .A(b[5]), .B(a[50]), .Z(n39060) );
  XOR U41589 ( .A(n39066), .B(n39067), .Z(n38741) );
  ANDN U41590 ( .B(n39068), .A(n39069), .Z(n39066) );
  AND U41591 ( .A(b[4]), .B(a[51]), .Z(n39065) );
  XOR U41592 ( .A(n39071), .B(n39072), .Z(n38746) );
  ANDN U41593 ( .B(n38758), .A(n38759), .Z(n39071) );
  AND U41594 ( .A(b[2]), .B(a[52]), .Z(n39073) );
  XNOR U41595 ( .A(n39068), .B(n39072), .Z(n39074) );
  XOR U41596 ( .A(n39075), .B(n39076), .Z(n39072) );
  OR U41597 ( .A(n38761), .B(n38762), .Z(n39076) );
  XNOR U41598 ( .A(n39078), .B(n39079), .Z(n39077) );
  XOR U41599 ( .A(n39078), .B(n39081), .Z(n38761) );
  NAND U41600 ( .A(b[1]), .B(a[52]), .Z(n39081) );
  IV U41601 ( .A(n39075), .Z(n39078) );
  NANDN U41602 ( .A(n105), .B(n106), .Z(n39075) );
  XOR U41603 ( .A(n39082), .B(n39083), .Z(n106) );
  NAND U41604 ( .A(a[52]), .B(b[0]), .Z(n105) );
  XNOR U41605 ( .A(n39063), .B(n39067), .Z(n39084) );
  XNOR U41606 ( .A(n39058), .B(n39062), .Z(n39085) );
  XNOR U41607 ( .A(n39053), .B(n39057), .Z(n39086) );
  XNOR U41608 ( .A(n39048), .B(n39052), .Z(n39087) );
  XNOR U41609 ( .A(n39043), .B(n39047), .Z(n39088) );
  XNOR U41610 ( .A(n39038), .B(n39042), .Z(n39089) );
  XNOR U41611 ( .A(n39033), .B(n39037), .Z(n39090) );
  XNOR U41612 ( .A(n39028), .B(n39032), .Z(n39091) );
  XNOR U41613 ( .A(n39023), .B(n39027), .Z(n39092) );
  XNOR U41614 ( .A(n39018), .B(n39022), .Z(n39093) );
  XNOR U41615 ( .A(n39013), .B(n39017), .Z(n39094) );
  XNOR U41616 ( .A(n39008), .B(n39012), .Z(n39095) );
  XNOR U41617 ( .A(n39003), .B(n39007), .Z(n39096) );
  XNOR U41618 ( .A(n38998), .B(n39002), .Z(n39097) );
  XNOR U41619 ( .A(n38993), .B(n38997), .Z(n39098) );
  XNOR U41620 ( .A(n38988), .B(n38992), .Z(n39099) );
  XNOR U41621 ( .A(n38983), .B(n38987), .Z(n39100) );
  XNOR U41622 ( .A(n38978), .B(n38982), .Z(n39101) );
  XNOR U41623 ( .A(n38973), .B(n38977), .Z(n39102) );
  XNOR U41624 ( .A(n38968), .B(n38972), .Z(n39103) );
  XNOR U41625 ( .A(n38963), .B(n38967), .Z(n39104) );
  XNOR U41626 ( .A(n38958), .B(n38962), .Z(n39105) );
  XNOR U41627 ( .A(n38953), .B(n38957), .Z(n39106) );
  XNOR U41628 ( .A(n38948), .B(n38952), .Z(n39107) );
  XNOR U41629 ( .A(n38943), .B(n38947), .Z(n39108) );
  XNOR U41630 ( .A(n38938), .B(n38942), .Z(n39109) );
  XNOR U41631 ( .A(n38933), .B(n38937), .Z(n39110) );
  XNOR U41632 ( .A(n38928), .B(n38932), .Z(n39111) );
  XNOR U41633 ( .A(n38923), .B(n38927), .Z(n39112) );
  XNOR U41634 ( .A(n38918), .B(n38922), .Z(n39113) );
  XNOR U41635 ( .A(n38913), .B(n38917), .Z(n39114) );
  XNOR U41636 ( .A(n38908), .B(n38912), .Z(n39115) );
  XNOR U41637 ( .A(n38903), .B(n38907), .Z(n39116) );
  XNOR U41638 ( .A(n38898), .B(n38902), .Z(n39117) );
  XNOR U41639 ( .A(n38893), .B(n38897), .Z(n39118) );
  XNOR U41640 ( .A(n38888), .B(n38892), .Z(n39119) );
  XNOR U41641 ( .A(n38883), .B(n38887), .Z(n39120) );
  XNOR U41642 ( .A(n38878), .B(n38882), .Z(n39121) );
  XNOR U41643 ( .A(n38873), .B(n38877), .Z(n39122) );
  XNOR U41644 ( .A(n38868), .B(n38872), .Z(n39123) );
  XNOR U41645 ( .A(n38863), .B(n38867), .Z(n39124) );
  XNOR U41646 ( .A(n38858), .B(n38862), .Z(n39125) );
  XNOR U41647 ( .A(n38853), .B(n38857), .Z(n39126) );
  XNOR U41648 ( .A(n38848), .B(n38852), .Z(n39127) );
  XNOR U41649 ( .A(n38843), .B(n38847), .Z(n39128) );
  XNOR U41650 ( .A(n38838), .B(n38842), .Z(n39129) );
  XNOR U41651 ( .A(n38833), .B(n38837), .Z(n39130) );
  XNOR U41652 ( .A(n38828), .B(n38832), .Z(n39131) );
  XNOR U41653 ( .A(n38823), .B(n38827), .Z(n39132) );
  XNOR U41654 ( .A(n38818), .B(n38822), .Z(n39133) );
  XOR U41655 ( .A(n39134), .B(n38817), .Z(n38818) );
  AND U41656 ( .A(a[0]), .B(b[54]), .Z(n39134) );
  XNOR U41657 ( .A(n39135), .B(n38817), .Z(n38819) );
  XNOR U41658 ( .A(n39136), .B(n39137), .Z(n38817) );
  ANDN U41659 ( .B(n39138), .A(n39139), .Z(n39136) );
  AND U41660 ( .A(a[1]), .B(b[53]), .Z(n39135) );
  XOR U41661 ( .A(n39141), .B(n39142), .Z(n38822) );
  ANDN U41662 ( .B(n39143), .A(n39144), .Z(n39141) );
  AND U41663 ( .A(a[2]), .B(b[52]), .Z(n39140) );
  XOR U41664 ( .A(n39146), .B(n39147), .Z(n38827) );
  ANDN U41665 ( .B(n39148), .A(n39149), .Z(n39146) );
  AND U41666 ( .A(a[3]), .B(b[51]), .Z(n39145) );
  XOR U41667 ( .A(n39151), .B(n39152), .Z(n38832) );
  ANDN U41668 ( .B(n39153), .A(n39154), .Z(n39151) );
  AND U41669 ( .A(a[4]), .B(b[50]), .Z(n39150) );
  XOR U41670 ( .A(n39156), .B(n39157), .Z(n38837) );
  ANDN U41671 ( .B(n39158), .A(n39159), .Z(n39156) );
  AND U41672 ( .A(a[5]), .B(b[49]), .Z(n39155) );
  XOR U41673 ( .A(n39161), .B(n39162), .Z(n38842) );
  ANDN U41674 ( .B(n39163), .A(n39164), .Z(n39161) );
  AND U41675 ( .A(a[6]), .B(b[48]), .Z(n39160) );
  XOR U41676 ( .A(n39166), .B(n39167), .Z(n38847) );
  ANDN U41677 ( .B(n39168), .A(n39169), .Z(n39166) );
  AND U41678 ( .A(a[7]), .B(b[47]), .Z(n39165) );
  XOR U41679 ( .A(n39171), .B(n39172), .Z(n38852) );
  ANDN U41680 ( .B(n39173), .A(n39174), .Z(n39171) );
  AND U41681 ( .A(a[8]), .B(b[46]), .Z(n39170) );
  XOR U41682 ( .A(n39176), .B(n39177), .Z(n38857) );
  ANDN U41683 ( .B(n39178), .A(n39179), .Z(n39176) );
  AND U41684 ( .A(a[9]), .B(b[45]), .Z(n39175) );
  XOR U41685 ( .A(n39181), .B(n39182), .Z(n38862) );
  ANDN U41686 ( .B(n39183), .A(n39184), .Z(n39181) );
  AND U41687 ( .A(a[10]), .B(b[44]), .Z(n39180) );
  XOR U41688 ( .A(n39186), .B(n39187), .Z(n38867) );
  ANDN U41689 ( .B(n39188), .A(n39189), .Z(n39186) );
  AND U41690 ( .A(a[11]), .B(b[43]), .Z(n39185) );
  XOR U41691 ( .A(n39191), .B(n39192), .Z(n38872) );
  ANDN U41692 ( .B(n39193), .A(n39194), .Z(n39191) );
  AND U41693 ( .A(a[12]), .B(b[42]), .Z(n39190) );
  XOR U41694 ( .A(n39196), .B(n39197), .Z(n38877) );
  ANDN U41695 ( .B(n39198), .A(n39199), .Z(n39196) );
  AND U41696 ( .A(a[13]), .B(b[41]), .Z(n39195) );
  XOR U41697 ( .A(n39201), .B(n39202), .Z(n38882) );
  ANDN U41698 ( .B(n39203), .A(n39204), .Z(n39201) );
  AND U41699 ( .A(a[14]), .B(b[40]), .Z(n39200) );
  XOR U41700 ( .A(n39206), .B(n39207), .Z(n38887) );
  ANDN U41701 ( .B(n39208), .A(n39209), .Z(n39206) );
  AND U41702 ( .A(a[15]), .B(b[39]), .Z(n39205) );
  XOR U41703 ( .A(n39211), .B(n39212), .Z(n38892) );
  ANDN U41704 ( .B(n39213), .A(n39214), .Z(n39211) );
  AND U41705 ( .A(a[16]), .B(b[38]), .Z(n39210) );
  XOR U41706 ( .A(n39216), .B(n39217), .Z(n38897) );
  ANDN U41707 ( .B(n39218), .A(n39219), .Z(n39216) );
  AND U41708 ( .A(a[17]), .B(b[37]), .Z(n39215) );
  XOR U41709 ( .A(n39221), .B(n39222), .Z(n38902) );
  ANDN U41710 ( .B(n39223), .A(n39224), .Z(n39221) );
  AND U41711 ( .A(a[18]), .B(b[36]), .Z(n39220) );
  XOR U41712 ( .A(n39226), .B(n39227), .Z(n38907) );
  ANDN U41713 ( .B(n39228), .A(n39229), .Z(n39226) );
  AND U41714 ( .A(a[19]), .B(b[35]), .Z(n39225) );
  XOR U41715 ( .A(n39231), .B(n39232), .Z(n38912) );
  ANDN U41716 ( .B(n39233), .A(n39234), .Z(n39231) );
  AND U41717 ( .A(a[20]), .B(b[34]), .Z(n39230) );
  XOR U41718 ( .A(n39236), .B(n39237), .Z(n38917) );
  ANDN U41719 ( .B(n39238), .A(n39239), .Z(n39236) );
  AND U41720 ( .A(a[21]), .B(b[33]), .Z(n39235) );
  XOR U41721 ( .A(n39241), .B(n39242), .Z(n38922) );
  ANDN U41722 ( .B(n39243), .A(n39244), .Z(n39241) );
  AND U41723 ( .A(a[22]), .B(b[32]), .Z(n39240) );
  XOR U41724 ( .A(n39246), .B(n39247), .Z(n38927) );
  ANDN U41725 ( .B(n39248), .A(n39249), .Z(n39246) );
  AND U41726 ( .A(a[23]), .B(b[31]), .Z(n39245) );
  XOR U41727 ( .A(n39251), .B(n39252), .Z(n38932) );
  ANDN U41728 ( .B(n39253), .A(n39254), .Z(n39251) );
  AND U41729 ( .A(a[24]), .B(b[30]), .Z(n39250) );
  XOR U41730 ( .A(n39256), .B(n39257), .Z(n38937) );
  ANDN U41731 ( .B(n39258), .A(n39259), .Z(n39256) );
  AND U41732 ( .A(a[25]), .B(b[29]), .Z(n39255) );
  XOR U41733 ( .A(n39261), .B(n39262), .Z(n38942) );
  ANDN U41734 ( .B(n39263), .A(n39264), .Z(n39261) );
  AND U41735 ( .A(a[26]), .B(b[28]), .Z(n39260) );
  XOR U41736 ( .A(n39266), .B(n39267), .Z(n38947) );
  ANDN U41737 ( .B(n39268), .A(n39269), .Z(n39266) );
  AND U41738 ( .A(a[27]), .B(b[27]), .Z(n39265) );
  XOR U41739 ( .A(n39271), .B(n39272), .Z(n38952) );
  ANDN U41740 ( .B(n39273), .A(n39274), .Z(n39271) );
  AND U41741 ( .A(a[28]), .B(b[26]), .Z(n39270) );
  XOR U41742 ( .A(n39276), .B(n39277), .Z(n38957) );
  ANDN U41743 ( .B(n39278), .A(n39279), .Z(n39276) );
  AND U41744 ( .A(a[29]), .B(b[25]), .Z(n39275) );
  XOR U41745 ( .A(n39281), .B(n39282), .Z(n38962) );
  ANDN U41746 ( .B(n39283), .A(n39284), .Z(n39281) );
  AND U41747 ( .A(a[30]), .B(b[24]), .Z(n39280) );
  XOR U41748 ( .A(n39286), .B(n39287), .Z(n38967) );
  ANDN U41749 ( .B(n39288), .A(n39289), .Z(n39286) );
  AND U41750 ( .A(a[31]), .B(b[23]), .Z(n39285) );
  XOR U41751 ( .A(n39291), .B(n39292), .Z(n38972) );
  ANDN U41752 ( .B(n39293), .A(n39294), .Z(n39291) );
  AND U41753 ( .A(a[32]), .B(b[22]), .Z(n39290) );
  XOR U41754 ( .A(n39296), .B(n39297), .Z(n38977) );
  ANDN U41755 ( .B(n39298), .A(n39299), .Z(n39296) );
  AND U41756 ( .A(a[33]), .B(b[21]), .Z(n39295) );
  XOR U41757 ( .A(n39301), .B(n39302), .Z(n38982) );
  ANDN U41758 ( .B(n39303), .A(n39304), .Z(n39301) );
  AND U41759 ( .A(a[34]), .B(b[20]), .Z(n39300) );
  XOR U41760 ( .A(n39306), .B(n39307), .Z(n38987) );
  ANDN U41761 ( .B(n39308), .A(n39309), .Z(n39306) );
  AND U41762 ( .A(a[35]), .B(b[19]), .Z(n39305) );
  XOR U41763 ( .A(n39311), .B(n39312), .Z(n38992) );
  ANDN U41764 ( .B(n39313), .A(n39314), .Z(n39311) );
  AND U41765 ( .A(a[36]), .B(b[18]), .Z(n39310) );
  XOR U41766 ( .A(n39316), .B(n39317), .Z(n38997) );
  ANDN U41767 ( .B(n39318), .A(n39319), .Z(n39316) );
  AND U41768 ( .A(a[37]), .B(b[17]), .Z(n39315) );
  XOR U41769 ( .A(n39321), .B(n39322), .Z(n39002) );
  ANDN U41770 ( .B(n39323), .A(n39324), .Z(n39321) );
  AND U41771 ( .A(a[38]), .B(b[16]), .Z(n39320) );
  XOR U41772 ( .A(n39326), .B(n39327), .Z(n39007) );
  ANDN U41773 ( .B(n39328), .A(n39329), .Z(n39326) );
  AND U41774 ( .A(a[39]), .B(b[15]), .Z(n39325) );
  XOR U41775 ( .A(n39331), .B(n39332), .Z(n39012) );
  ANDN U41776 ( .B(n39333), .A(n39334), .Z(n39331) );
  AND U41777 ( .A(a[40]), .B(b[14]), .Z(n39330) );
  XOR U41778 ( .A(n39336), .B(n39337), .Z(n39017) );
  ANDN U41779 ( .B(n39338), .A(n39339), .Z(n39336) );
  AND U41780 ( .A(a[41]), .B(b[13]), .Z(n39335) );
  XOR U41781 ( .A(n39341), .B(n39342), .Z(n39022) );
  ANDN U41782 ( .B(n39343), .A(n39344), .Z(n39341) );
  AND U41783 ( .A(a[42]), .B(b[12]), .Z(n39340) );
  XOR U41784 ( .A(n39346), .B(n39347), .Z(n39027) );
  ANDN U41785 ( .B(n39348), .A(n39349), .Z(n39346) );
  AND U41786 ( .A(a[43]), .B(b[11]), .Z(n39345) );
  XOR U41787 ( .A(n39351), .B(n39352), .Z(n39032) );
  ANDN U41788 ( .B(n39353), .A(n39354), .Z(n39351) );
  AND U41789 ( .A(a[44]), .B(b[10]), .Z(n39350) );
  XOR U41790 ( .A(n39356), .B(n39357), .Z(n39037) );
  ANDN U41791 ( .B(n39358), .A(n39359), .Z(n39356) );
  AND U41792 ( .A(b[9]), .B(a[45]), .Z(n39355) );
  XOR U41793 ( .A(n39361), .B(n39362), .Z(n39042) );
  ANDN U41794 ( .B(n39363), .A(n39364), .Z(n39361) );
  AND U41795 ( .A(b[8]), .B(a[46]), .Z(n39360) );
  XOR U41796 ( .A(n39366), .B(n39367), .Z(n39047) );
  ANDN U41797 ( .B(n39368), .A(n39369), .Z(n39366) );
  AND U41798 ( .A(b[7]), .B(a[47]), .Z(n39365) );
  XOR U41799 ( .A(n39371), .B(n39372), .Z(n39052) );
  ANDN U41800 ( .B(n39373), .A(n39374), .Z(n39371) );
  AND U41801 ( .A(b[6]), .B(a[48]), .Z(n39370) );
  XOR U41802 ( .A(n39376), .B(n39377), .Z(n39057) );
  ANDN U41803 ( .B(n39378), .A(n39379), .Z(n39376) );
  AND U41804 ( .A(b[5]), .B(a[49]), .Z(n39375) );
  XOR U41805 ( .A(n39381), .B(n39382), .Z(n39062) );
  ANDN U41806 ( .B(n39383), .A(n39384), .Z(n39381) );
  AND U41807 ( .A(b[4]), .B(a[50]), .Z(n39380) );
  XOR U41808 ( .A(n39386), .B(n39387), .Z(n39067) );
  ANDN U41809 ( .B(n39079), .A(n39080), .Z(n39386) );
  AND U41810 ( .A(b[2]), .B(a[51]), .Z(n39388) );
  XNOR U41811 ( .A(n39383), .B(n39387), .Z(n39389) );
  XOR U41812 ( .A(n39390), .B(n39391), .Z(n39387) );
  OR U41813 ( .A(n39082), .B(n39083), .Z(n39391) );
  XNOR U41814 ( .A(n39393), .B(n39394), .Z(n39392) );
  XOR U41815 ( .A(n39393), .B(n39396), .Z(n39082) );
  NAND U41816 ( .A(b[1]), .B(a[51]), .Z(n39396) );
  IV U41817 ( .A(n39390), .Z(n39393) );
  NANDN U41818 ( .A(n107), .B(n108), .Z(n39390) );
  XOR U41819 ( .A(n39397), .B(n39398), .Z(n108) );
  NAND U41820 ( .A(a[51]), .B(b[0]), .Z(n107) );
  XNOR U41821 ( .A(n39378), .B(n39382), .Z(n39399) );
  XNOR U41822 ( .A(n39373), .B(n39377), .Z(n39400) );
  XNOR U41823 ( .A(n39368), .B(n39372), .Z(n39401) );
  XNOR U41824 ( .A(n39363), .B(n39367), .Z(n39402) );
  XNOR U41825 ( .A(n39358), .B(n39362), .Z(n39403) );
  XNOR U41826 ( .A(n39353), .B(n39357), .Z(n39404) );
  XNOR U41827 ( .A(n39348), .B(n39352), .Z(n39405) );
  XNOR U41828 ( .A(n39343), .B(n39347), .Z(n39406) );
  XNOR U41829 ( .A(n39338), .B(n39342), .Z(n39407) );
  XNOR U41830 ( .A(n39333), .B(n39337), .Z(n39408) );
  XNOR U41831 ( .A(n39328), .B(n39332), .Z(n39409) );
  XNOR U41832 ( .A(n39323), .B(n39327), .Z(n39410) );
  XNOR U41833 ( .A(n39318), .B(n39322), .Z(n39411) );
  XNOR U41834 ( .A(n39313), .B(n39317), .Z(n39412) );
  XNOR U41835 ( .A(n39308), .B(n39312), .Z(n39413) );
  XNOR U41836 ( .A(n39303), .B(n39307), .Z(n39414) );
  XNOR U41837 ( .A(n39298), .B(n39302), .Z(n39415) );
  XNOR U41838 ( .A(n39293), .B(n39297), .Z(n39416) );
  XNOR U41839 ( .A(n39288), .B(n39292), .Z(n39417) );
  XNOR U41840 ( .A(n39283), .B(n39287), .Z(n39418) );
  XNOR U41841 ( .A(n39278), .B(n39282), .Z(n39419) );
  XNOR U41842 ( .A(n39273), .B(n39277), .Z(n39420) );
  XNOR U41843 ( .A(n39268), .B(n39272), .Z(n39421) );
  XNOR U41844 ( .A(n39263), .B(n39267), .Z(n39422) );
  XNOR U41845 ( .A(n39258), .B(n39262), .Z(n39423) );
  XNOR U41846 ( .A(n39253), .B(n39257), .Z(n39424) );
  XNOR U41847 ( .A(n39248), .B(n39252), .Z(n39425) );
  XNOR U41848 ( .A(n39243), .B(n39247), .Z(n39426) );
  XNOR U41849 ( .A(n39238), .B(n39242), .Z(n39427) );
  XNOR U41850 ( .A(n39233), .B(n39237), .Z(n39428) );
  XNOR U41851 ( .A(n39228), .B(n39232), .Z(n39429) );
  XNOR U41852 ( .A(n39223), .B(n39227), .Z(n39430) );
  XNOR U41853 ( .A(n39218), .B(n39222), .Z(n39431) );
  XNOR U41854 ( .A(n39213), .B(n39217), .Z(n39432) );
  XNOR U41855 ( .A(n39208), .B(n39212), .Z(n39433) );
  XNOR U41856 ( .A(n39203), .B(n39207), .Z(n39434) );
  XNOR U41857 ( .A(n39198), .B(n39202), .Z(n39435) );
  XNOR U41858 ( .A(n39193), .B(n39197), .Z(n39436) );
  XNOR U41859 ( .A(n39188), .B(n39192), .Z(n39437) );
  XNOR U41860 ( .A(n39183), .B(n39187), .Z(n39438) );
  XNOR U41861 ( .A(n39178), .B(n39182), .Z(n39439) );
  XNOR U41862 ( .A(n39173), .B(n39177), .Z(n39440) );
  XNOR U41863 ( .A(n39168), .B(n39172), .Z(n39441) );
  XNOR U41864 ( .A(n39163), .B(n39167), .Z(n39442) );
  XNOR U41865 ( .A(n39158), .B(n39162), .Z(n39443) );
  XNOR U41866 ( .A(n39153), .B(n39157), .Z(n39444) );
  XNOR U41867 ( .A(n39148), .B(n39152), .Z(n39445) );
  XNOR U41868 ( .A(n39143), .B(n39147), .Z(n39446) );
  XNOR U41869 ( .A(n39138), .B(n39142), .Z(n39447) );
  XNOR U41870 ( .A(n39448), .B(n39137), .Z(n39138) );
  AND U41871 ( .A(a[0]), .B(b[53]), .Z(n39448) );
  XOR U41872 ( .A(n39449), .B(n39137), .Z(n39139) );
  XNOR U41873 ( .A(n39450), .B(n39451), .Z(n39137) );
  ANDN U41874 ( .B(n39452), .A(n39453), .Z(n39450) );
  AND U41875 ( .A(a[1]), .B(b[52]), .Z(n39449) );
  XOR U41876 ( .A(n39455), .B(n39456), .Z(n39142) );
  ANDN U41877 ( .B(n39457), .A(n39458), .Z(n39455) );
  AND U41878 ( .A(a[2]), .B(b[51]), .Z(n39454) );
  XOR U41879 ( .A(n39460), .B(n39461), .Z(n39147) );
  ANDN U41880 ( .B(n39462), .A(n39463), .Z(n39460) );
  AND U41881 ( .A(a[3]), .B(b[50]), .Z(n39459) );
  XOR U41882 ( .A(n39465), .B(n39466), .Z(n39152) );
  ANDN U41883 ( .B(n39467), .A(n39468), .Z(n39465) );
  AND U41884 ( .A(a[4]), .B(b[49]), .Z(n39464) );
  XOR U41885 ( .A(n39470), .B(n39471), .Z(n39157) );
  ANDN U41886 ( .B(n39472), .A(n39473), .Z(n39470) );
  AND U41887 ( .A(a[5]), .B(b[48]), .Z(n39469) );
  XOR U41888 ( .A(n39475), .B(n39476), .Z(n39162) );
  ANDN U41889 ( .B(n39477), .A(n39478), .Z(n39475) );
  AND U41890 ( .A(a[6]), .B(b[47]), .Z(n39474) );
  XOR U41891 ( .A(n39480), .B(n39481), .Z(n39167) );
  ANDN U41892 ( .B(n39482), .A(n39483), .Z(n39480) );
  AND U41893 ( .A(a[7]), .B(b[46]), .Z(n39479) );
  XOR U41894 ( .A(n39485), .B(n39486), .Z(n39172) );
  ANDN U41895 ( .B(n39487), .A(n39488), .Z(n39485) );
  AND U41896 ( .A(a[8]), .B(b[45]), .Z(n39484) );
  XOR U41897 ( .A(n39490), .B(n39491), .Z(n39177) );
  ANDN U41898 ( .B(n39492), .A(n39493), .Z(n39490) );
  AND U41899 ( .A(a[9]), .B(b[44]), .Z(n39489) );
  XOR U41900 ( .A(n39495), .B(n39496), .Z(n39182) );
  ANDN U41901 ( .B(n39497), .A(n39498), .Z(n39495) );
  AND U41902 ( .A(a[10]), .B(b[43]), .Z(n39494) );
  XOR U41903 ( .A(n39500), .B(n39501), .Z(n39187) );
  ANDN U41904 ( .B(n39502), .A(n39503), .Z(n39500) );
  AND U41905 ( .A(a[11]), .B(b[42]), .Z(n39499) );
  XOR U41906 ( .A(n39505), .B(n39506), .Z(n39192) );
  ANDN U41907 ( .B(n39507), .A(n39508), .Z(n39505) );
  AND U41908 ( .A(a[12]), .B(b[41]), .Z(n39504) );
  XOR U41909 ( .A(n39510), .B(n39511), .Z(n39197) );
  ANDN U41910 ( .B(n39512), .A(n39513), .Z(n39510) );
  AND U41911 ( .A(a[13]), .B(b[40]), .Z(n39509) );
  XOR U41912 ( .A(n39515), .B(n39516), .Z(n39202) );
  ANDN U41913 ( .B(n39517), .A(n39518), .Z(n39515) );
  AND U41914 ( .A(a[14]), .B(b[39]), .Z(n39514) );
  XOR U41915 ( .A(n39520), .B(n39521), .Z(n39207) );
  ANDN U41916 ( .B(n39522), .A(n39523), .Z(n39520) );
  AND U41917 ( .A(a[15]), .B(b[38]), .Z(n39519) );
  XOR U41918 ( .A(n39525), .B(n39526), .Z(n39212) );
  ANDN U41919 ( .B(n39527), .A(n39528), .Z(n39525) );
  AND U41920 ( .A(a[16]), .B(b[37]), .Z(n39524) );
  XOR U41921 ( .A(n39530), .B(n39531), .Z(n39217) );
  ANDN U41922 ( .B(n39532), .A(n39533), .Z(n39530) );
  AND U41923 ( .A(a[17]), .B(b[36]), .Z(n39529) );
  XOR U41924 ( .A(n39535), .B(n39536), .Z(n39222) );
  ANDN U41925 ( .B(n39537), .A(n39538), .Z(n39535) );
  AND U41926 ( .A(a[18]), .B(b[35]), .Z(n39534) );
  XOR U41927 ( .A(n39540), .B(n39541), .Z(n39227) );
  ANDN U41928 ( .B(n39542), .A(n39543), .Z(n39540) );
  AND U41929 ( .A(a[19]), .B(b[34]), .Z(n39539) );
  XOR U41930 ( .A(n39545), .B(n39546), .Z(n39232) );
  ANDN U41931 ( .B(n39547), .A(n39548), .Z(n39545) );
  AND U41932 ( .A(a[20]), .B(b[33]), .Z(n39544) );
  XOR U41933 ( .A(n39550), .B(n39551), .Z(n39237) );
  ANDN U41934 ( .B(n39552), .A(n39553), .Z(n39550) );
  AND U41935 ( .A(a[21]), .B(b[32]), .Z(n39549) );
  XOR U41936 ( .A(n39555), .B(n39556), .Z(n39242) );
  ANDN U41937 ( .B(n39557), .A(n39558), .Z(n39555) );
  AND U41938 ( .A(a[22]), .B(b[31]), .Z(n39554) );
  XOR U41939 ( .A(n39560), .B(n39561), .Z(n39247) );
  ANDN U41940 ( .B(n39562), .A(n39563), .Z(n39560) );
  AND U41941 ( .A(a[23]), .B(b[30]), .Z(n39559) );
  XOR U41942 ( .A(n39565), .B(n39566), .Z(n39252) );
  ANDN U41943 ( .B(n39567), .A(n39568), .Z(n39565) );
  AND U41944 ( .A(a[24]), .B(b[29]), .Z(n39564) );
  XOR U41945 ( .A(n39570), .B(n39571), .Z(n39257) );
  ANDN U41946 ( .B(n39572), .A(n39573), .Z(n39570) );
  AND U41947 ( .A(a[25]), .B(b[28]), .Z(n39569) );
  XOR U41948 ( .A(n39575), .B(n39576), .Z(n39262) );
  ANDN U41949 ( .B(n39577), .A(n39578), .Z(n39575) );
  AND U41950 ( .A(a[26]), .B(b[27]), .Z(n39574) );
  XOR U41951 ( .A(n39580), .B(n39581), .Z(n39267) );
  ANDN U41952 ( .B(n39582), .A(n39583), .Z(n39580) );
  AND U41953 ( .A(a[27]), .B(b[26]), .Z(n39579) );
  XOR U41954 ( .A(n39585), .B(n39586), .Z(n39272) );
  ANDN U41955 ( .B(n39587), .A(n39588), .Z(n39585) );
  AND U41956 ( .A(a[28]), .B(b[25]), .Z(n39584) );
  XOR U41957 ( .A(n39590), .B(n39591), .Z(n39277) );
  ANDN U41958 ( .B(n39592), .A(n39593), .Z(n39590) );
  AND U41959 ( .A(a[29]), .B(b[24]), .Z(n39589) );
  XOR U41960 ( .A(n39595), .B(n39596), .Z(n39282) );
  ANDN U41961 ( .B(n39597), .A(n39598), .Z(n39595) );
  AND U41962 ( .A(a[30]), .B(b[23]), .Z(n39594) );
  XOR U41963 ( .A(n39600), .B(n39601), .Z(n39287) );
  ANDN U41964 ( .B(n39602), .A(n39603), .Z(n39600) );
  AND U41965 ( .A(a[31]), .B(b[22]), .Z(n39599) );
  XOR U41966 ( .A(n39605), .B(n39606), .Z(n39292) );
  ANDN U41967 ( .B(n39607), .A(n39608), .Z(n39605) );
  AND U41968 ( .A(a[32]), .B(b[21]), .Z(n39604) );
  XOR U41969 ( .A(n39610), .B(n39611), .Z(n39297) );
  ANDN U41970 ( .B(n39612), .A(n39613), .Z(n39610) );
  AND U41971 ( .A(a[33]), .B(b[20]), .Z(n39609) );
  XOR U41972 ( .A(n39615), .B(n39616), .Z(n39302) );
  ANDN U41973 ( .B(n39617), .A(n39618), .Z(n39615) );
  AND U41974 ( .A(a[34]), .B(b[19]), .Z(n39614) );
  XOR U41975 ( .A(n39620), .B(n39621), .Z(n39307) );
  ANDN U41976 ( .B(n39622), .A(n39623), .Z(n39620) );
  AND U41977 ( .A(a[35]), .B(b[18]), .Z(n39619) );
  XOR U41978 ( .A(n39625), .B(n39626), .Z(n39312) );
  ANDN U41979 ( .B(n39627), .A(n39628), .Z(n39625) );
  AND U41980 ( .A(a[36]), .B(b[17]), .Z(n39624) );
  XOR U41981 ( .A(n39630), .B(n39631), .Z(n39317) );
  ANDN U41982 ( .B(n39632), .A(n39633), .Z(n39630) );
  AND U41983 ( .A(a[37]), .B(b[16]), .Z(n39629) );
  XOR U41984 ( .A(n39635), .B(n39636), .Z(n39322) );
  ANDN U41985 ( .B(n39637), .A(n39638), .Z(n39635) );
  AND U41986 ( .A(a[38]), .B(b[15]), .Z(n39634) );
  XOR U41987 ( .A(n39640), .B(n39641), .Z(n39327) );
  ANDN U41988 ( .B(n39642), .A(n39643), .Z(n39640) );
  AND U41989 ( .A(a[39]), .B(b[14]), .Z(n39639) );
  XOR U41990 ( .A(n39645), .B(n39646), .Z(n39332) );
  ANDN U41991 ( .B(n39647), .A(n39648), .Z(n39645) );
  AND U41992 ( .A(a[40]), .B(b[13]), .Z(n39644) );
  XOR U41993 ( .A(n39650), .B(n39651), .Z(n39337) );
  ANDN U41994 ( .B(n39652), .A(n39653), .Z(n39650) );
  AND U41995 ( .A(a[41]), .B(b[12]), .Z(n39649) );
  XOR U41996 ( .A(n39655), .B(n39656), .Z(n39342) );
  ANDN U41997 ( .B(n39657), .A(n39658), .Z(n39655) );
  AND U41998 ( .A(a[42]), .B(b[11]), .Z(n39654) );
  XOR U41999 ( .A(n39660), .B(n39661), .Z(n39347) );
  ANDN U42000 ( .B(n39662), .A(n39663), .Z(n39660) );
  AND U42001 ( .A(a[43]), .B(b[10]), .Z(n39659) );
  XOR U42002 ( .A(n39665), .B(n39666), .Z(n39352) );
  ANDN U42003 ( .B(n39667), .A(n39668), .Z(n39665) );
  AND U42004 ( .A(b[9]), .B(a[44]), .Z(n39664) );
  XOR U42005 ( .A(n39670), .B(n39671), .Z(n39357) );
  ANDN U42006 ( .B(n39672), .A(n39673), .Z(n39670) );
  AND U42007 ( .A(b[8]), .B(a[45]), .Z(n39669) );
  XOR U42008 ( .A(n39675), .B(n39676), .Z(n39362) );
  ANDN U42009 ( .B(n39677), .A(n39678), .Z(n39675) );
  AND U42010 ( .A(b[7]), .B(a[46]), .Z(n39674) );
  XOR U42011 ( .A(n39680), .B(n39681), .Z(n39367) );
  ANDN U42012 ( .B(n39682), .A(n39683), .Z(n39680) );
  AND U42013 ( .A(b[6]), .B(a[47]), .Z(n39679) );
  XOR U42014 ( .A(n39685), .B(n39686), .Z(n39372) );
  ANDN U42015 ( .B(n39687), .A(n39688), .Z(n39685) );
  AND U42016 ( .A(b[5]), .B(a[48]), .Z(n39684) );
  XOR U42017 ( .A(n39690), .B(n39691), .Z(n39377) );
  ANDN U42018 ( .B(n39692), .A(n39693), .Z(n39690) );
  AND U42019 ( .A(b[4]), .B(a[49]), .Z(n39689) );
  XOR U42020 ( .A(n39695), .B(n39696), .Z(n39382) );
  ANDN U42021 ( .B(n39394), .A(n39395), .Z(n39695) );
  AND U42022 ( .A(b[2]), .B(a[50]), .Z(n39697) );
  XNOR U42023 ( .A(n39692), .B(n39696), .Z(n39698) );
  XOR U42024 ( .A(n39699), .B(n39700), .Z(n39696) );
  OR U42025 ( .A(n39397), .B(n39398), .Z(n39700) );
  XNOR U42026 ( .A(n39702), .B(n39703), .Z(n39701) );
  XOR U42027 ( .A(n39702), .B(n39705), .Z(n39397) );
  NAND U42028 ( .A(b[1]), .B(a[50]), .Z(n39705) );
  IV U42029 ( .A(n39699), .Z(n39702) );
  NANDN U42030 ( .A(n109), .B(n110), .Z(n39699) );
  XOR U42031 ( .A(n39706), .B(n39707), .Z(n110) );
  NAND U42032 ( .A(a[50]), .B(b[0]), .Z(n109) );
  XNOR U42033 ( .A(n39687), .B(n39691), .Z(n39708) );
  XNOR U42034 ( .A(n39682), .B(n39686), .Z(n39709) );
  XNOR U42035 ( .A(n39677), .B(n39681), .Z(n39710) );
  XNOR U42036 ( .A(n39672), .B(n39676), .Z(n39711) );
  XNOR U42037 ( .A(n39667), .B(n39671), .Z(n39712) );
  XNOR U42038 ( .A(n39662), .B(n39666), .Z(n39713) );
  XNOR U42039 ( .A(n39657), .B(n39661), .Z(n39714) );
  XNOR U42040 ( .A(n39652), .B(n39656), .Z(n39715) );
  XNOR U42041 ( .A(n39647), .B(n39651), .Z(n39716) );
  XNOR U42042 ( .A(n39642), .B(n39646), .Z(n39717) );
  XNOR U42043 ( .A(n39637), .B(n39641), .Z(n39718) );
  XNOR U42044 ( .A(n39632), .B(n39636), .Z(n39719) );
  XNOR U42045 ( .A(n39627), .B(n39631), .Z(n39720) );
  XNOR U42046 ( .A(n39622), .B(n39626), .Z(n39721) );
  XNOR U42047 ( .A(n39617), .B(n39621), .Z(n39722) );
  XNOR U42048 ( .A(n39612), .B(n39616), .Z(n39723) );
  XNOR U42049 ( .A(n39607), .B(n39611), .Z(n39724) );
  XNOR U42050 ( .A(n39602), .B(n39606), .Z(n39725) );
  XNOR U42051 ( .A(n39597), .B(n39601), .Z(n39726) );
  XNOR U42052 ( .A(n39592), .B(n39596), .Z(n39727) );
  XNOR U42053 ( .A(n39587), .B(n39591), .Z(n39728) );
  XNOR U42054 ( .A(n39582), .B(n39586), .Z(n39729) );
  XNOR U42055 ( .A(n39577), .B(n39581), .Z(n39730) );
  XNOR U42056 ( .A(n39572), .B(n39576), .Z(n39731) );
  XNOR U42057 ( .A(n39567), .B(n39571), .Z(n39732) );
  XNOR U42058 ( .A(n39562), .B(n39566), .Z(n39733) );
  XNOR U42059 ( .A(n39557), .B(n39561), .Z(n39734) );
  XNOR U42060 ( .A(n39552), .B(n39556), .Z(n39735) );
  XNOR U42061 ( .A(n39547), .B(n39551), .Z(n39736) );
  XNOR U42062 ( .A(n39542), .B(n39546), .Z(n39737) );
  XNOR U42063 ( .A(n39537), .B(n39541), .Z(n39738) );
  XNOR U42064 ( .A(n39532), .B(n39536), .Z(n39739) );
  XNOR U42065 ( .A(n39527), .B(n39531), .Z(n39740) );
  XNOR U42066 ( .A(n39522), .B(n39526), .Z(n39741) );
  XNOR U42067 ( .A(n39517), .B(n39521), .Z(n39742) );
  XNOR U42068 ( .A(n39512), .B(n39516), .Z(n39743) );
  XNOR U42069 ( .A(n39507), .B(n39511), .Z(n39744) );
  XNOR U42070 ( .A(n39502), .B(n39506), .Z(n39745) );
  XNOR U42071 ( .A(n39497), .B(n39501), .Z(n39746) );
  XNOR U42072 ( .A(n39492), .B(n39496), .Z(n39747) );
  XNOR U42073 ( .A(n39487), .B(n39491), .Z(n39748) );
  XNOR U42074 ( .A(n39482), .B(n39486), .Z(n39749) );
  XNOR U42075 ( .A(n39477), .B(n39481), .Z(n39750) );
  XNOR U42076 ( .A(n39472), .B(n39476), .Z(n39751) );
  XNOR U42077 ( .A(n39467), .B(n39471), .Z(n39752) );
  XNOR U42078 ( .A(n39462), .B(n39466), .Z(n39753) );
  XNOR U42079 ( .A(n39457), .B(n39461), .Z(n39754) );
  XNOR U42080 ( .A(n39452), .B(n39456), .Z(n39755) );
  XOR U42081 ( .A(n39756), .B(n39451), .Z(n39452) );
  AND U42082 ( .A(a[0]), .B(b[52]), .Z(n39756) );
  XNOR U42083 ( .A(n39757), .B(n39451), .Z(n39453) );
  XNOR U42084 ( .A(n39758), .B(n39759), .Z(n39451) );
  ANDN U42085 ( .B(n39760), .A(n39761), .Z(n39758) );
  AND U42086 ( .A(a[1]), .B(b[51]), .Z(n39757) );
  XOR U42087 ( .A(n39763), .B(n39764), .Z(n39456) );
  ANDN U42088 ( .B(n39765), .A(n39766), .Z(n39763) );
  AND U42089 ( .A(a[2]), .B(b[50]), .Z(n39762) );
  XOR U42090 ( .A(n39768), .B(n39769), .Z(n39461) );
  ANDN U42091 ( .B(n39770), .A(n39771), .Z(n39768) );
  AND U42092 ( .A(a[3]), .B(b[49]), .Z(n39767) );
  XOR U42093 ( .A(n39773), .B(n39774), .Z(n39466) );
  ANDN U42094 ( .B(n39775), .A(n39776), .Z(n39773) );
  AND U42095 ( .A(a[4]), .B(b[48]), .Z(n39772) );
  XOR U42096 ( .A(n39778), .B(n39779), .Z(n39471) );
  ANDN U42097 ( .B(n39780), .A(n39781), .Z(n39778) );
  AND U42098 ( .A(a[5]), .B(b[47]), .Z(n39777) );
  XOR U42099 ( .A(n39783), .B(n39784), .Z(n39476) );
  ANDN U42100 ( .B(n39785), .A(n39786), .Z(n39783) );
  AND U42101 ( .A(a[6]), .B(b[46]), .Z(n39782) );
  XOR U42102 ( .A(n39788), .B(n39789), .Z(n39481) );
  ANDN U42103 ( .B(n39790), .A(n39791), .Z(n39788) );
  AND U42104 ( .A(a[7]), .B(b[45]), .Z(n39787) );
  XOR U42105 ( .A(n39793), .B(n39794), .Z(n39486) );
  ANDN U42106 ( .B(n39795), .A(n39796), .Z(n39793) );
  AND U42107 ( .A(a[8]), .B(b[44]), .Z(n39792) );
  XOR U42108 ( .A(n39798), .B(n39799), .Z(n39491) );
  ANDN U42109 ( .B(n39800), .A(n39801), .Z(n39798) );
  AND U42110 ( .A(a[9]), .B(b[43]), .Z(n39797) );
  XOR U42111 ( .A(n39803), .B(n39804), .Z(n39496) );
  ANDN U42112 ( .B(n39805), .A(n39806), .Z(n39803) );
  AND U42113 ( .A(a[10]), .B(b[42]), .Z(n39802) );
  XOR U42114 ( .A(n39808), .B(n39809), .Z(n39501) );
  ANDN U42115 ( .B(n39810), .A(n39811), .Z(n39808) );
  AND U42116 ( .A(a[11]), .B(b[41]), .Z(n39807) );
  XOR U42117 ( .A(n39813), .B(n39814), .Z(n39506) );
  ANDN U42118 ( .B(n39815), .A(n39816), .Z(n39813) );
  AND U42119 ( .A(a[12]), .B(b[40]), .Z(n39812) );
  XOR U42120 ( .A(n39818), .B(n39819), .Z(n39511) );
  ANDN U42121 ( .B(n39820), .A(n39821), .Z(n39818) );
  AND U42122 ( .A(a[13]), .B(b[39]), .Z(n39817) );
  XOR U42123 ( .A(n39823), .B(n39824), .Z(n39516) );
  ANDN U42124 ( .B(n39825), .A(n39826), .Z(n39823) );
  AND U42125 ( .A(a[14]), .B(b[38]), .Z(n39822) );
  XOR U42126 ( .A(n39828), .B(n39829), .Z(n39521) );
  ANDN U42127 ( .B(n39830), .A(n39831), .Z(n39828) );
  AND U42128 ( .A(a[15]), .B(b[37]), .Z(n39827) );
  XOR U42129 ( .A(n39833), .B(n39834), .Z(n39526) );
  ANDN U42130 ( .B(n39835), .A(n39836), .Z(n39833) );
  AND U42131 ( .A(a[16]), .B(b[36]), .Z(n39832) );
  XOR U42132 ( .A(n39838), .B(n39839), .Z(n39531) );
  ANDN U42133 ( .B(n39840), .A(n39841), .Z(n39838) );
  AND U42134 ( .A(a[17]), .B(b[35]), .Z(n39837) );
  XOR U42135 ( .A(n39843), .B(n39844), .Z(n39536) );
  ANDN U42136 ( .B(n39845), .A(n39846), .Z(n39843) );
  AND U42137 ( .A(a[18]), .B(b[34]), .Z(n39842) );
  XOR U42138 ( .A(n39848), .B(n39849), .Z(n39541) );
  ANDN U42139 ( .B(n39850), .A(n39851), .Z(n39848) );
  AND U42140 ( .A(a[19]), .B(b[33]), .Z(n39847) );
  XOR U42141 ( .A(n39853), .B(n39854), .Z(n39546) );
  ANDN U42142 ( .B(n39855), .A(n39856), .Z(n39853) );
  AND U42143 ( .A(a[20]), .B(b[32]), .Z(n39852) );
  XOR U42144 ( .A(n39858), .B(n39859), .Z(n39551) );
  ANDN U42145 ( .B(n39860), .A(n39861), .Z(n39858) );
  AND U42146 ( .A(a[21]), .B(b[31]), .Z(n39857) );
  XOR U42147 ( .A(n39863), .B(n39864), .Z(n39556) );
  ANDN U42148 ( .B(n39865), .A(n39866), .Z(n39863) );
  AND U42149 ( .A(a[22]), .B(b[30]), .Z(n39862) );
  XOR U42150 ( .A(n39868), .B(n39869), .Z(n39561) );
  ANDN U42151 ( .B(n39870), .A(n39871), .Z(n39868) );
  AND U42152 ( .A(a[23]), .B(b[29]), .Z(n39867) );
  XOR U42153 ( .A(n39873), .B(n39874), .Z(n39566) );
  ANDN U42154 ( .B(n39875), .A(n39876), .Z(n39873) );
  AND U42155 ( .A(a[24]), .B(b[28]), .Z(n39872) );
  XOR U42156 ( .A(n39878), .B(n39879), .Z(n39571) );
  ANDN U42157 ( .B(n39880), .A(n39881), .Z(n39878) );
  AND U42158 ( .A(a[25]), .B(b[27]), .Z(n39877) );
  XOR U42159 ( .A(n39883), .B(n39884), .Z(n39576) );
  ANDN U42160 ( .B(n39885), .A(n39886), .Z(n39883) );
  AND U42161 ( .A(a[26]), .B(b[26]), .Z(n39882) );
  XOR U42162 ( .A(n39888), .B(n39889), .Z(n39581) );
  ANDN U42163 ( .B(n39890), .A(n39891), .Z(n39888) );
  AND U42164 ( .A(a[27]), .B(b[25]), .Z(n39887) );
  XOR U42165 ( .A(n39893), .B(n39894), .Z(n39586) );
  ANDN U42166 ( .B(n39895), .A(n39896), .Z(n39893) );
  AND U42167 ( .A(a[28]), .B(b[24]), .Z(n39892) );
  XOR U42168 ( .A(n39898), .B(n39899), .Z(n39591) );
  ANDN U42169 ( .B(n39900), .A(n39901), .Z(n39898) );
  AND U42170 ( .A(a[29]), .B(b[23]), .Z(n39897) );
  XOR U42171 ( .A(n39903), .B(n39904), .Z(n39596) );
  ANDN U42172 ( .B(n39905), .A(n39906), .Z(n39903) );
  AND U42173 ( .A(a[30]), .B(b[22]), .Z(n39902) );
  XOR U42174 ( .A(n39908), .B(n39909), .Z(n39601) );
  ANDN U42175 ( .B(n39910), .A(n39911), .Z(n39908) );
  AND U42176 ( .A(a[31]), .B(b[21]), .Z(n39907) );
  XOR U42177 ( .A(n39913), .B(n39914), .Z(n39606) );
  ANDN U42178 ( .B(n39915), .A(n39916), .Z(n39913) );
  AND U42179 ( .A(a[32]), .B(b[20]), .Z(n39912) );
  XOR U42180 ( .A(n39918), .B(n39919), .Z(n39611) );
  ANDN U42181 ( .B(n39920), .A(n39921), .Z(n39918) );
  AND U42182 ( .A(a[33]), .B(b[19]), .Z(n39917) );
  XOR U42183 ( .A(n39923), .B(n39924), .Z(n39616) );
  ANDN U42184 ( .B(n39925), .A(n39926), .Z(n39923) );
  AND U42185 ( .A(a[34]), .B(b[18]), .Z(n39922) );
  XOR U42186 ( .A(n39928), .B(n39929), .Z(n39621) );
  ANDN U42187 ( .B(n39930), .A(n39931), .Z(n39928) );
  AND U42188 ( .A(a[35]), .B(b[17]), .Z(n39927) );
  XOR U42189 ( .A(n39933), .B(n39934), .Z(n39626) );
  ANDN U42190 ( .B(n39935), .A(n39936), .Z(n39933) );
  AND U42191 ( .A(a[36]), .B(b[16]), .Z(n39932) );
  XOR U42192 ( .A(n39938), .B(n39939), .Z(n39631) );
  ANDN U42193 ( .B(n39940), .A(n39941), .Z(n39938) );
  AND U42194 ( .A(a[37]), .B(b[15]), .Z(n39937) );
  XOR U42195 ( .A(n39943), .B(n39944), .Z(n39636) );
  ANDN U42196 ( .B(n39945), .A(n39946), .Z(n39943) );
  AND U42197 ( .A(a[38]), .B(b[14]), .Z(n39942) );
  XOR U42198 ( .A(n39948), .B(n39949), .Z(n39641) );
  ANDN U42199 ( .B(n39950), .A(n39951), .Z(n39948) );
  AND U42200 ( .A(a[39]), .B(b[13]), .Z(n39947) );
  XOR U42201 ( .A(n39953), .B(n39954), .Z(n39646) );
  ANDN U42202 ( .B(n39955), .A(n39956), .Z(n39953) );
  AND U42203 ( .A(a[40]), .B(b[12]), .Z(n39952) );
  XOR U42204 ( .A(n39958), .B(n39959), .Z(n39651) );
  ANDN U42205 ( .B(n39960), .A(n39961), .Z(n39958) );
  AND U42206 ( .A(a[41]), .B(b[11]), .Z(n39957) );
  XOR U42207 ( .A(n39963), .B(n39964), .Z(n39656) );
  ANDN U42208 ( .B(n39965), .A(n39966), .Z(n39963) );
  AND U42209 ( .A(a[42]), .B(b[10]), .Z(n39962) );
  XOR U42210 ( .A(n39968), .B(n39969), .Z(n39661) );
  ANDN U42211 ( .B(n39970), .A(n39971), .Z(n39968) );
  AND U42212 ( .A(b[9]), .B(a[43]), .Z(n39967) );
  XOR U42213 ( .A(n39973), .B(n39974), .Z(n39666) );
  ANDN U42214 ( .B(n39975), .A(n39976), .Z(n39973) );
  AND U42215 ( .A(b[8]), .B(a[44]), .Z(n39972) );
  XOR U42216 ( .A(n39978), .B(n39979), .Z(n39671) );
  ANDN U42217 ( .B(n39980), .A(n39981), .Z(n39978) );
  AND U42218 ( .A(b[7]), .B(a[45]), .Z(n39977) );
  XOR U42219 ( .A(n39983), .B(n39984), .Z(n39676) );
  ANDN U42220 ( .B(n39985), .A(n39986), .Z(n39983) );
  AND U42221 ( .A(b[6]), .B(a[46]), .Z(n39982) );
  XOR U42222 ( .A(n39988), .B(n39989), .Z(n39681) );
  ANDN U42223 ( .B(n39990), .A(n39991), .Z(n39988) );
  AND U42224 ( .A(b[5]), .B(a[47]), .Z(n39987) );
  XOR U42225 ( .A(n39993), .B(n39994), .Z(n39686) );
  ANDN U42226 ( .B(n39995), .A(n39996), .Z(n39993) );
  AND U42227 ( .A(b[4]), .B(a[48]), .Z(n39992) );
  XOR U42228 ( .A(n39998), .B(n39999), .Z(n39691) );
  ANDN U42229 ( .B(n39703), .A(n39704), .Z(n39998) );
  AND U42230 ( .A(b[2]), .B(a[49]), .Z(n40000) );
  XNOR U42231 ( .A(n39995), .B(n39999), .Z(n40001) );
  XOR U42232 ( .A(n40002), .B(n40003), .Z(n39999) );
  OR U42233 ( .A(n39706), .B(n39707), .Z(n40003) );
  XNOR U42234 ( .A(n40005), .B(n40006), .Z(n40004) );
  XOR U42235 ( .A(n40005), .B(n40008), .Z(n39706) );
  NAND U42236 ( .A(b[1]), .B(a[49]), .Z(n40008) );
  IV U42237 ( .A(n40002), .Z(n40005) );
  NANDN U42238 ( .A(n113), .B(n114), .Z(n40002) );
  XOR U42239 ( .A(n40009), .B(n40010), .Z(n114) );
  NAND U42240 ( .A(a[49]), .B(b[0]), .Z(n113) );
  XNOR U42241 ( .A(n39990), .B(n39994), .Z(n40011) );
  XNOR U42242 ( .A(n39985), .B(n39989), .Z(n40012) );
  XNOR U42243 ( .A(n39980), .B(n39984), .Z(n40013) );
  XNOR U42244 ( .A(n39975), .B(n39979), .Z(n40014) );
  XNOR U42245 ( .A(n39970), .B(n39974), .Z(n40015) );
  XNOR U42246 ( .A(n39965), .B(n39969), .Z(n40016) );
  XNOR U42247 ( .A(n39960), .B(n39964), .Z(n40017) );
  XNOR U42248 ( .A(n39955), .B(n39959), .Z(n40018) );
  XNOR U42249 ( .A(n39950), .B(n39954), .Z(n40019) );
  XNOR U42250 ( .A(n39945), .B(n39949), .Z(n40020) );
  XNOR U42251 ( .A(n39940), .B(n39944), .Z(n40021) );
  XNOR U42252 ( .A(n39935), .B(n39939), .Z(n40022) );
  XNOR U42253 ( .A(n39930), .B(n39934), .Z(n40023) );
  XNOR U42254 ( .A(n39925), .B(n39929), .Z(n40024) );
  XNOR U42255 ( .A(n39920), .B(n39924), .Z(n40025) );
  XNOR U42256 ( .A(n39915), .B(n39919), .Z(n40026) );
  XNOR U42257 ( .A(n39910), .B(n39914), .Z(n40027) );
  XNOR U42258 ( .A(n39905), .B(n39909), .Z(n40028) );
  XNOR U42259 ( .A(n39900), .B(n39904), .Z(n40029) );
  XNOR U42260 ( .A(n39895), .B(n39899), .Z(n40030) );
  XNOR U42261 ( .A(n39890), .B(n39894), .Z(n40031) );
  XNOR U42262 ( .A(n39885), .B(n39889), .Z(n40032) );
  XNOR U42263 ( .A(n39880), .B(n39884), .Z(n40033) );
  XNOR U42264 ( .A(n39875), .B(n39879), .Z(n40034) );
  XNOR U42265 ( .A(n39870), .B(n39874), .Z(n40035) );
  XNOR U42266 ( .A(n39865), .B(n39869), .Z(n40036) );
  XNOR U42267 ( .A(n39860), .B(n39864), .Z(n40037) );
  XNOR U42268 ( .A(n39855), .B(n39859), .Z(n40038) );
  XNOR U42269 ( .A(n39850), .B(n39854), .Z(n40039) );
  XNOR U42270 ( .A(n39845), .B(n39849), .Z(n40040) );
  XNOR U42271 ( .A(n39840), .B(n39844), .Z(n40041) );
  XNOR U42272 ( .A(n39835), .B(n39839), .Z(n40042) );
  XNOR U42273 ( .A(n39830), .B(n39834), .Z(n40043) );
  XNOR U42274 ( .A(n39825), .B(n39829), .Z(n40044) );
  XNOR U42275 ( .A(n39820), .B(n39824), .Z(n40045) );
  XNOR U42276 ( .A(n39815), .B(n39819), .Z(n40046) );
  XNOR U42277 ( .A(n39810), .B(n39814), .Z(n40047) );
  XNOR U42278 ( .A(n39805), .B(n39809), .Z(n40048) );
  XNOR U42279 ( .A(n39800), .B(n39804), .Z(n40049) );
  XNOR U42280 ( .A(n39795), .B(n39799), .Z(n40050) );
  XNOR U42281 ( .A(n39790), .B(n39794), .Z(n40051) );
  XNOR U42282 ( .A(n39785), .B(n39789), .Z(n40052) );
  XNOR U42283 ( .A(n39780), .B(n39784), .Z(n40053) );
  XNOR U42284 ( .A(n39775), .B(n39779), .Z(n40054) );
  XNOR U42285 ( .A(n39770), .B(n39774), .Z(n40055) );
  XNOR U42286 ( .A(n39765), .B(n39769), .Z(n40056) );
  XNOR U42287 ( .A(n39760), .B(n39764), .Z(n40057) );
  XNOR U42288 ( .A(n40058), .B(n39759), .Z(n39760) );
  AND U42289 ( .A(a[0]), .B(b[51]), .Z(n40058) );
  XOR U42290 ( .A(n40059), .B(n39759), .Z(n39761) );
  XNOR U42291 ( .A(n40060), .B(n40061), .Z(n39759) );
  ANDN U42292 ( .B(n40062), .A(n40063), .Z(n40060) );
  AND U42293 ( .A(a[1]), .B(b[50]), .Z(n40059) );
  XOR U42294 ( .A(n40065), .B(n40066), .Z(n39764) );
  ANDN U42295 ( .B(n40067), .A(n40068), .Z(n40065) );
  AND U42296 ( .A(a[2]), .B(b[49]), .Z(n40064) );
  XOR U42297 ( .A(n40070), .B(n40071), .Z(n39769) );
  ANDN U42298 ( .B(n40072), .A(n40073), .Z(n40070) );
  AND U42299 ( .A(a[3]), .B(b[48]), .Z(n40069) );
  XOR U42300 ( .A(n40075), .B(n40076), .Z(n39774) );
  ANDN U42301 ( .B(n40077), .A(n40078), .Z(n40075) );
  AND U42302 ( .A(a[4]), .B(b[47]), .Z(n40074) );
  XOR U42303 ( .A(n40080), .B(n40081), .Z(n39779) );
  ANDN U42304 ( .B(n40082), .A(n40083), .Z(n40080) );
  AND U42305 ( .A(a[5]), .B(b[46]), .Z(n40079) );
  XOR U42306 ( .A(n40085), .B(n40086), .Z(n39784) );
  ANDN U42307 ( .B(n40087), .A(n40088), .Z(n40085) );
  AND U42308 ( .A(a[6]), .B(b[45]), .Z(n40084) );
  XOR U42309 ( .A(n40090), .B(n40091), .Z(n39789) );
  ANDN U42310 ( .B(n40092), .A(n40093), .Z(n40090) );
  AND U42311 ( .A(a[7]), .B(b[44]), .Z(n40089) );
  XOR U42312 ( .A(n40095), .B(n40096), .Z(n39794) );
  ANDN U42313 ( .B(n40097), .A(n40098), .Z(n40095) );
  AND U42314 ( .A(a[8]), .B(b[43]), .Z(n40094) );
  XOR U42315 ( .A(n40100), .B(n40101), .Z(n39799) );
  ANDN U42316 ( .B(n40102), .A(n40103), .Z(n40100) );
  AND U42317 ( .A(a[9]), .B(b[42]), .Z(n40099) );
  XOR U42318 ( .A(n40105), .B(n40106), .Z(n39804) );
  ANDN U42319 ( .B(n40107), .A(n40108), .Z(n40105) );
  AND U42320 ( .A(a[10]), .B(b[41]), .Z(n40104) );
  XOR U42321 ( .A(n40110), .B(n40111), .Z(n39809) );
  ANDN U42322 ( .B(n40112), .A(n40113), .Z(n40110) );
  AND U42323 ( .A(a[11]), .B(b[40]), .Z(n40109) );
  XOR U42324 ( .A(n40115), .B(n40116), .Z(n39814) );
  ANDN U42325 ( .B(n40117), .A(n40118), .Z(n40115) );
  AND U42326 ( .A(a[12]), .B(b[39]), .Z(n40114) );
  XOR U42327 ( .A(n40120), .B(n40121), .Z(n39819) );
  ANDN U42328 ( .B(n40122), .A(n40123), .Z(n40120) );
  AND U42329 ( .A(a[13]), .B(b[38]), .Z(n40119) );
  XOR U42330 ( .A(n40125), .B(n40126), .Z(n39824) );
  ANDN U42331 ( .B(n40127), .A(n40128), .Z(n40125) );
  AND U42332 ( .A(a[14]), .B(b[37]), .Z(n40124) );
  XOR U42333 ( .A(n40130), .B(n40131), .Z(n39829) );
  ANDN U42334 ( .B(n40132), .A(n40133), .Z(n40130) );
  AND U42335 ( .A(a[15]), .B(b[36]), .Z(n40129) );
  XOR U42336 ( .A(n40135), .B(n40136), .Z(n39834) );
  ANDN U42337 ( .B(n40137), .A(n40138), .Z(n40135) );
  AND U42338 ( .A(a[16]), .B(b[35]), .Z(n40134) );
  XOR U42339 ( .A(n40140), .B(n40141), .Z(n39839) );
  ANDN U42340 ( .B(n40142), .A(n40143), .Z(n40140) );
  AND U42341 ( .A(a[17]), .B(b[34]), .Z(n40139) );
  XOR U42342 ( .A(n40145), .B(n40146), .Z(n39844) );
  ANDN U42343 ( .B(n40147), .A(n40148), .Z(n40145) );
  AND U42344 ( .A(a[18]), .B(b[33]), .Z(n40144) );
  XOR U42345 ( .A(n40150), .B(n40151), .Z(n39849) );
  ANDN U42346 ( .B(n40152), .A(n40153), .Z(n40150) );
  AND U42347 ( .A(a[19]), .B(b[32]), .Z(n40149) );
  XOR U42348 ( .A(n40155), .B(n40156), .Z(n39854) );
  ANDN U42349 ( .B(n40157), .A(n40158), .Z(n40155) );
  AND U42350 ( .A(a[20]), .B(b[31]), .Z(n40154) );
  XOR U42351 ( .A(n40160), .B(n40161), .Z(n39859) );
  ANDN U42352 ( .B(n40162), .A(n40163), .Z(n40160) );
  AND U42353 ( .A(a[21]), .B(b[30]), .Z(n40159) );
  XOR U42354 ( .A(n40165), .B(n40166), .Z(n39864) );
  ANDN U42355 ( .B(n40167), .A(n40168), .Z(n40165) );
  AND U42356 ( .A(a[22]), .B(b[29]), .Z(n40164) );
  XOR U42357 ( .A(n40170), .B(n40171), .Z(n39869) );
  ANDN U42358 ( .B(n40172), .A(n40173), .Z(n40170) );
  AND U42359 ( .A(a[23]), .B(b[28]), .Z(n40169) );
  XOR U42360 ( .A(n40175), .B(n40176), .Z(n39874) );
  ANDN U42361 ( .B(n40177), .A(n40178), .Z(n40175) );
  AND U42362 ( .A(a[24]), .B(b[27]), .Z(n40174) );
  XOR U42363 ( .A(n40180), .B(n40181), .Z(n39879) );
  ANDN U42364 ( .B(n40182), .A(n40183), .Z(n40180) );
  AND U42365 ( .A(a[25]), .B(b[26]), .Z(n40179) );
  XOR U42366 ( .A(n40185), .B(n40186), .Z(n39884) );
  ANDN U42367 ( .B(n40187), .A(n40188), .Z(n40185) );
  AND U42368 ( .A(a[26]), .B(b[25]), .Z(n40184) );
  XOR U42369 ( .A(n40190), .B(n40191), .Z(n39889) );
  ANDN U42370 ( .B(n40192), .A(n40193), .Z(n40190) );
  AND U42371 ( .A(a[27]), .B(b[24]), .Z(n40189) );
  XOR U42372 ( .A(n40195), .B(n40196), .Z(n39894) );
  ANDN U42373 ( .B(n40197), .A(n40198), .Z(n40195) );
  AND U42374 ( .A(a[28]), .B(b[23]), .Z(n40194) );
  XOR U42375 ( .A(n40200), .B(n40201), .Z(n39899) );
  ANDN U42376 ( .B(n40202), .A(n40203), .Z(n40200) );
  AND U42377 ( .A(a[29]), .B(b[22]), .Z(n40199) );
  XOR U42378 ( .A(n40205), .B(n40206), .Z(n39904) );
  ANDN U42379 ( .B(n40207), .A(n40208), .Z(n40205) );
  AND U42380 ( .A(a[30]), .B(b[21]), .Z(n40204) );
  XOR U42381 ( .A(n40210), .B(n40211), .Z(n39909) );
  ANDN U42382 ( .B(n40212), .A(n40213), .Z(n40210) );
  AND U42383 ( .A(a[31]), .B(b[20]), .Z(n40209) );
  XOR U42384 ( .A(n40215), .B(n40216), .Z(n39914) );
  ANDN U42385 ( .B(n40217), .A(n40218), .Z(n40215) );
  AND U42386 ( .A(a[32]), .B(b[19]), .Z(n40214) );
  XOR U42387 ( .A(n40220), .B(n40221), .Z(n39919) );
  ANDN U42388 ( .B(n40222), .A(n40223), .Z(n40220) );
  AND U42389 ( .A(a[33]), .B(b[18]), .Z(n40219) );
  XOR U42390 ( .A(n40225), .B(n40226), .Z(n39924) );
  ANDN U42391 ( .B(n40227), .A(n40228), .Z(n40225) );
  AND U42392 ( .A(a[34]), .B(b[17]), .Z(n40224) );
  XOR U42393 ( .A(n40230), .B(n40231), .Z(n39929) );
  ANDN U42394 ( .B(n40232), .A(n40233), .Z(n40230) );
  AND U42395 ( .A(a[35]), .B(b[16]), .Z(n40229) );
  XOR U42396 ( .A(n40235), .B(n40236), .Z(n39934) );
  ANDN U42397 ( .B(n40237), .A(n40238), .Z(n40235) );
  AND U42398 ( .A(a[36]), .B(b[15]), .Z(n40234) );
  XOR U42399 ( .A(n40240), .B(n40241), .Z(n39939) );
  ANDN U42400 ( .B(n40242), .A(n40243), .Z(n40240) );
  AND U42401 ( .A(a[37]), .B(b[14]), .Z(n40239) );
  XOR U42402 ( .A(n40245), .B(n40246), .Z(n39944) );
  ANDN U42403 ( .B(n40247), .A(n40248), .Z(n40245) );
  AND U42404 ( .A(a[38]), .B(b[13]), .Z(n40244) );
  XOR U42405 ( .A(n40250), .B(n40251), .Z(n39949) );
  ANDN U42406 ( .B(n40252), .A(n40253), .Z(n40250) );
  AND U42407 ( .A(a[39]), .B(b[12]), .Z(n40249) );
  XOR U42408 ( .A(n40255), .B(n40256), .Z(n39954) );
  ANDN U42409 ( .B(n40257), .A(n40258), .Z(n40255) );
  AND U42410 ( .A(a[40]), .B(b[11]), .Z(n40254) );
  XOR U42411 ( .A(n40260), .B(n40261), .Z(n39959) );
  ANDN U42412 ( .B(n40262), .A(n40263), .Z(n40260) );
  AND U42413 ( .A(a[41]), .B(b[10]), .Z(n40259) );
  XOR U42414 ( .A(n40265), .B(n40266), .Z(n39964) );
  ANDN U42415 ( .B(n40267), .A(n40268), .Z(n40265) );
  AND U42416 ( .A(b[9]), .B(a[42]), .Z(n40264) );
  XOR U42417 ( .A(n40270), .B(n40271), .Z(n39969) );
  ANDN U42418 ( .B(n40272), .A(n40273), .Z(n40270) );
  AND U42419 ( .A(b[8]), .B(a[43]), .Z(n40269) );
  XOR U42420 ( .A(n40275), .B(n40276), .Z(n39974) );
  ANDN U42421 ( .B(n40277), .A(n40278), .Z(n40275) );
  AND U42422 ( .A(b[7]), .B(a[44]), .Z(n40274) );
  XOR U42423 ( .A(n40280), .B(n40281), .Z(n39979) );
  ANDN U42424 ( .B(n40282), .A(n40283), .Z(n40280) );
  AND U42425 ( .A(b[6]), .B(a[45]), .Z(n40279) );
  XOR U42426 ( .A(n40285), .B(n40286), .Z(n39984) );
  ANDN U42427 ( .B(n40287), .A(n40288), .Z(n40285) );
  AND U42428 ( .A(b[5]), .B(a[46]), .Z(n40284) );
  XOR U42429 ( .A(n40290), .B(n40291), .Z(n39989) );
  ANDN U42430 ( .B(n40292), .A(n40293), .Z(n40290) );
  AND U42431 ( .A(b[4]), .B(a[47]), .Z(n40289) );
  XOR U42432 ( .A(n40295), .B(n40296), .Z(n39994) );
  ANDN U42433 ( .B(n40006), .A(n40007), .Z(n40295) );
  AND U42434 ( .A(b[2]), .B(a[48]), .Z(n40297) );
  XNOR U42435 ( .A(n40292), .B(n40296), .Z(n40298) );
  XOR U42436 ( .A(n40299), .B(n40300), .Z(n40296) );
  OR U42437 ( .A(n40009), .B(n40010), .Z(n40300) );
  XNOR U42438 ( .A(n40302), .B(n40303), .Z(n40301) );
  XOR U42439 ( .A(n40302), .B(n40305), .Z(n40009) );
  NAND U42440 ( .A(b[1]), .B(a[48]), .Z(n40305) );
  IV U42441 ( .A(n40299), .Z(n40302) );
  NANDN U42442 ( .A(n115), .B(n116), .Z(n40299) );
  XOR U42443 ( .A(n40306), .B(n40307), .Z(n116) );
  NAND U42444 ( .A(a[48]), .B(b[0]), .Z(n115) );
  XNOR U42445 ( .A(n40287), .B(n40291), .Z(n40308) );
  XNOR U42446 ( .A(n40282), .B(n40286), .Z(n40309) );
  XNOR U42447 ( .A(n40277), .B(n40281), .Z(n40310) );
  XNOR U42448 ( .A(n40272), .B(n40276), .Z(n40311) );
  XNOR U42449 ( .A(n40267), .B(n40271), .Z(n40312) );
  XNOR U42450 ( .A(n40262), .B(n40266), .Z(n40313) );
  XNOR U42451 ( .A(n40257), .B(n40261), .Z(n40314) );
  XNOR U42452 ( .A(n40252), .B(n40256), .Z(n40315) );
  XNOR U42453 ( .A(n40247), .B(n40251), .Z(n40316) );
  XNOR U42454 ( .A(n40242), .B(n40246), .Z(n40317) );
  XNOR U42455 ( .A(n40237), .B(n40241), .Z(n40318) );
  XNOR U42456 ( .A(n40232), .B(n40236), .Z(n40319) );
  XNOR U42457 ( .A(n40227), .B(n40231), .Z(n40320) );
  XNOR U42458 ( .A(n40222), .B(n40226), .Z(n40321) );
  XNOR U42459 ( .A(n40217), .B(n40221), .Z(n40322) );
  XNOR U42460 ( .A(n40212), .B(n40216), .Z(n40323) );
  XNOR U42461 ( .A(n40207), .B(n40211), .Z(n40324) );
  XNOR U42462 ( .A(n40202), .B(n40206), .Z(n40325) );
  XNOR U42463 ( .A(n40197), .B(n40201), .Z(n40326) );
  XNOR U42464 ( .A(n40192), .B(n40196), .Z(n40327) );
  XNOR U42465 ( .A(n40187), .B(n40191), .Z(n40328) );
  XNOR U42466 ( .A(n40182), .B(n40186), .Z(n40329) );
  XNOR U42467 ( .A(n40177), .B(n40181), .Z(n40330) );
  XNOR U42468 ( .A(n40172), .B(n40176), .Z(n40331) );
  XNOR U42469 ( .A(n40167), .B(n40171), .Z(n40332) );
  XNOR U42470 ( .A(n40162), .B(n40166), .Z(n40333) );
  XNOR U42471 ( .A(n40157), .B(n40161), .Z(n40334) );
  XNOR U42472 ( .A(n40152), .B(n40156), .Z(n40335) );
  XNOR U42473 ( .A(n40147), .B(n40151), .Z(n40336) );
  XNOR U42474 ( .A(n40142), .B(n40146), .Z(n40337) );
  XNOR U42475 ( .A(n40137), .B(n40141), .Z(n40338) );
  XNOR U42476 ( .A(n40132), .B(n40136), .Z(n40339) );
  XNOR U42477 ( .A(n40127), .B(n40131), .Z(n40340) );
  XNOR U42478 ( .A(n40122), .B(n40126), .Z(n40341) );
  XNOR U42479 ( .A(n40117), .B(n40121), .Z(n40342) );
  XNOR U42480 ( .A(n40112), .B(n40116), .Z(n40343) );
  XNOR U42481 ( .A(n40107), .B(n40111), .Z(n40344) );
  XNOR U42482 ( .A(n40102), .B(n40106), .Z(n40345) );
  XNOR U42483 ( .A(n40097), .B(n40101), .Z(n40346) );
  XNOR U42484 ( .A(n40092), .B(n40096), .Z(n40347) );
  XNOR U42485 ( .A(n40087), .B(n40091), .Z(n40348) );
  XNOR U42486 ( .A(n40082), .B(n40086), .Z(n40349) );
  XNOR U42487 ( .A(n40077), .B(n40081), .Z(n40350) );
  XNOR U42488 ( .A(n40072), .B(n40076), .Z(n40351) );
  XNOR U42489 ( .A(n40067), .B(n40071), .Z(n40352) );
  XNOR U42490 ( .A(n40062), .B(n40066), .Z(n40353) );
  XOR U42491 ( .A(n40354), .B(n40061), .Z(n40062) );
  AND U42492 ( .A(a[0]), .B(b[50]), .Z(n40354) );
  XNOR U42493 ( .A(n40355), .B(n40061), .Z(n40063) );
  XNOR U42494 ( .A(n40356), .B(n40357), .Z(n40061) );
  ANDN U42495 ( .B(n40358), .A(n40359), .Z(n40356) );
  AND U42496 ( .A(a[1]), .B(b[49]), .Z(n40355) );
  XOR U42497 ( .A(n40361), .B(n40362), .Z(n40066) );
  ANDN U42498 ( .B(n40363), .A(n40364), .Z(n40361) );
  AND U42499 ( .A(a[2]), .B(b[48]), .Z(n40360) );
  XOR U42500 ( .A(n40366), .B(n40367), .Z(n40071) );
  ANDN U42501 ( .B(n40368), .A(n40369), .Z(n40366) );
  AND U42502 ( .A(a[3]), .B(b[47]), .Z(n40365) );
  XOR U42503 ( .A(n40371), .B(n40372), .Z(n40076) );
  ANDN U42504 ( .B(n40373), .A(n40374), .Z(n40371) );
  AND U42505 ( .A(a[4]), .B(b[46]), .Z(n40370) );
  XOR U42506 ( .A(n40376), .B(n40377), .Z(n40081) );
  ANDN U42507 ( .B(n40378), .A(n40379), .Z(n40376) );
  AND U42508 ( .A(a[5]), .B(b[45]), .Z(n40375) );
  XOR U42509 ( .A(n40381), .B(n40382), .Z(n40086) );
  ANDN U42510 ( .B(n40383), .A(n40384), .Z(n40381) );
  AND U42511 ( .A(a[6]), .B(b[44]), .Z(n40380) );
  XOR U42512 ( .A(n40386), .B(n40387), .Z(n40091) );
  ANDN U42513 ( .B(n40388), .A(n40389), .Z(n40386) );
  AND U42514 ( .A(a[7]), .B(b[43]), .Z(n40385) );
  XOR U42515 ( .A(n40391), .B(n40392), .Z(n40096) );
  ANDN U42516 ( .B(n40393), .A(n40394), .Z(n40391) );
  AND U42517 ( .A(a[8]), .B(b[42]), .Z(n40390) );
  XOR U42518 ( .A(n40396), .B(n40397), .Z(n40101) );
  ANDN U42519 ( .B(n40398), .A(n40399), .Z(n40396) );
  AND U42520 ( .A(a[9]), .B(b[41]), .Z(n40395) );
  XOR U42521 ( .A(n40401), .B(n40402), .Z(n40106) );
  ANDN U42522 ( .B(n40403), .A(n40404), .Z(n40401) );
  AND U42523 ( .A(a[10]), .B(b[40]), .Z(n40400) );
  XOR U42524 ( .A(n40406), .B(n40407), .Z(n40111) );
  ANDN U42525 ( .B(n40408), .A(n40409), .Z(n40406) );
  AND U42526 ( .A(a[11]), .B(b[39]), .Z(n40405) );
  XOR U42527 ( .A(n40411), .B(n40412), .Z(n40116) );
  ANDN U42528 ( .B(n40413), .A(n40414), .Z(n40411) );
  AND U42529 ( .A(a[12]), .B(b[38]), .Z(n40410) );
  XOR U42530 ( .A(n40416), .B(n40417), .Z(n40121) );
  ANDN U42531 ( .B(n40418), .A(n40419), .Z(n40416) );
  AND U42532 ( .A(a[13]), .B(b[37]), .Z(n40415) );
  XOR U42533 ( .A(n40421), .B(n40422), .Z(n40126) );
  ANDN U42534 ( .B(n40423), .A(n40424), .Z(n40421) );
  AND U42535 ( .A(a[14]), .B(b[36]), .Z(n40420) );
  XOR U42536 ( .A(n40426), .B(n40427), .Z(n40131) );
  ANDN U42537 ( .B(n40428), .A(n40429), .Z(n40426) );
  AND U42538 ( .A(a[15]), .B(b[35]), .Z(n40425) );
  XOR U42539 ( .A(n40431), .B(n40432), .Z(n40136) );
  ANDN U42540 ( .B(n40433), .A(n40434), .Z(n40431) );
  AND U42541 ( .A(a[16]), .B(b[34]), .Z(n40430) );
  XOR U42542 ( .A(n40436), .B(n40437), .Z(n40141) );
  ANDN U42543 ( .B(n40438), .A(n40439), .Z(n40436) );
  AND U42544 ( .A(a[17]), .B(b[33]), .Z(n40435) );
  XOR U42545 ( .A(n40441), .B(n40442), .Z(n40146) );
  ANDN U42546 ( .B(n40443), .A(n40444), .Z(n40441) );
  AND U42547 ( .A(a[18]), .B(b[32]), .Z(n40440) );
  XOR U42548 ( .A(n40446), .B(n40447), .Z(n40151) );
  ANDN U42549 ( .B(n40448), .A(n40449), .Z(n40446) );
  AND U42550 ( .A(a[19]), .B(b[31]), .Z(n40445) );
  XOR U42551 ( .A(n40451), .B(n40452), .Z(n40156) );
  ANDN U42552 ( .B(n40453), .A(n40454), .Z(n40451) );
  AND U42553 ( .A(a[20]), .B(b[30]), .Z(n40450) );
  XOR U42554 ( .A(n40456), .B(n40457), .Z(n40161) );
  ANDN U42555 ( .B(n40458), .A(n40459), .Z(n40456) );
  AND U42556 ( .A(a[21]), .B(b[29]), .Z(n40455) );
  XOR U42557 ( .A(n40461), .B(n40462), .Z(n40166) );
  ANDN U42558 ( .B(n40463), .A(n40464), .Z(n40461) );
  AND U42559 ( .A(a[22]), .B(b[28]), .Z(n40460) );
  XOR U42560 ( .A(n40466), .B(n40467), .Z(n40171) );
  ANDN U42561 ( .B(n40468), .A(n40469), .Z(n40466) );
  AND U42562 ( .A(a[23]), .B(b[27]), .Z(n40465) );
  XOR U42563 ( .A(n40471), .B(n40472), .Z(n40176) );
  ANDN U42564 ( .B(n40473), .A(n40474), .Z(n40471) );
  AND U42565 ( .A(a[24]), .B(b[26]), .Z(n40470) );
  XOR U42566 ( .A(n40476), .B(n40477), .Z(n40181) );
  ANDN U42567 ( .B(n40478), .A(n40479), .Z(n40476) );
  AND U42568 ( .A(a[25]), .B(b[25]), .Z(n40475) );
  XOR U42569 ( .A(n40481), .B(n40482), .Z(n40186) );
  ANDN U42570 ( .B(n40483), .A(n40484), .Z(n40481) );
  AND U42571 ( .A(a[26]), .B(b[24]), .Z(n40480) );
  XOR U42572 ( .A(n40486), .B(n40487), .Z(n40191) );
  ANDN U42573 ( .B(n40488), .A(n40489), .Z(n40486) );
  AND U42574 ( .A(a[27]), .B(b[23]), .Z(n40485) );
  XOR U42575 ( .A(n40491), .B(n40492), .Z(n40196) );
  ANDN U42576 ( .B(n40493), .A(n40494), .Z(n40491) );
  AND U42577 ( .A(a[28]), .B(b[22]), .Z(n40490) );
  XOR U42578 ( .A(n40496), .B(n40497), .Z(n40201) );
  ANDN U42579 ( .B(n40498), .A(n40499), .Z(n40496) );
  AND U42580 ( .A(a[29]), .B(b[21]), .Z(n40495) );
  XOR U42581 ( .A(n40501), .B(n40502), .Z(n40206) );
  ANDN U42582 ( .B(n40503), .A(n40504), .Z(n40501) );
  AND U42583 ( .A(a[30]), .B(b[20]), .Z(n40500) );
  XOR U42584 ( .A(n40506), .B(n40507), .Z(n40211) );
  ANDN U42585 ( .B(n40508), .A(n40509), .Z(n40506) );
  AND U42586 ( .A(a[31]), .B(b[19]), .Z(n40505) );
  XOR U42587 ( .A(n40511), .B(n40512), .Z(n40216) );
  ANDN U42588 ( .B(n40513), .A(n40514), .Z(n40511) );
  AND U42589 ( .A(a[32]), .B(b[18]), .Z(n40510) );
  XOR U42590 ( .A(n40516), .B(n40517), .Z(n40221) );
  ANDN U42591 ( .B(n40518), .A(n40519), .Z(n40516) );
  AND U42592 ( .A(a[33]), .B(b[17]), .Z(n40515) );
  XOR U42593 ( .A(n40521), .B(n40522), .Z(n40226) );
  ANDN U42594 ( .B(n40523), .A(n40524), .Z(n40521) );
  AND U42595 ( .A(a[34]), .B(b[16]), .Z(n40520) );
  XOR U42596 ( .A(n40526), .B(n40527), .Z(n40231) );
  ANDN U42597 ( .B(n40528), .A(n40529), .Z(n40526) );
  AND U42598 ( .A(a[35]), .B(b[15]), .Z(n40525) );
  XOR U42599 ( .A(n40531), .B(n40532), .Z(n40236) );
  ANDN U42600 ( .B(n40533), .A(n40534), .Z(n40531) );
  AND U42601 ( .A(a[36]), .B(b[14]), .Z(n40530) );
  XOR U42602 ( .A(n40536), .B(n40537), .Z(n40241) );
  ANDN U42603 ( .B(n40538), .A(n40539), .Z(n40536) );
  AND U42604 ( .A(a[37]), .B(b[13]), .Z(n40535) );
  XOR U42605 ( .A(n40541), .B(n40542), .Z(n40246) );
  ANDN U42606 ( .B(n40543), .A(n40544), .Z(n40541) );
  AND U42607 ( .A(a[38]), .B(b[12]), .Z(n40540) );
  XOR U42608 ( .A(n40546), .B(n40547), .Z(n40251) );
  ANDN U42609 ( .B(n40548), .A(n40549), .Z(n40546) );
  AND U42610 ( .A(a[39]), .B(b[11]), .Z(n40545) );
  XOR U42611 ( .A(n40551), .B(n40552), .Z(n40256) );
  ANDN U42612 ( .B(n40553), .A(n40554), .Z(n40551) );
  AND U42613 ( .A(a[40]), .B(b[10]), .Z(n40550) );
  XOR U42614 ( .A(n40556), .B(n40557), .Z(n40261) );
  ANDN U42615 ( .B(n40558), .A(n40559), .Z(n40556) );
  AND U42616 ( .A(b[9]), .B(a[41]), .Z(n40555) );
  XOR U42617 ( .A(n40561), .B(n40562), .Z(n40266) );
  ANDN U42618 ( .B(n40563), .A(n40564), .Z(n40561) );
  AND U42619 ( .A(b[8]), .B(a[42]), .Z(n40560) );
  XOR U42620 ( .A(n40566), .B(n40567), .Z(n40271) );
  ANDN U42621 ( .B(n40568), .A(n40569), .Z(n40566) );
  AND U42622 ( .A(b[7]), .B(a[43]), .Z(n40565) );
  XOR U42623 ( .A(n40571), .B(n40572), .Z(n40276) );
  ANDN U42624 ( .B(n40573), .A(n40574), .Z(n40571) );
  AND U42625 ( .A(b[6]), .B(a[44]), .Z(n40570) );
  XOR U42626 ( .A(n40576), .B(n40577), .Z(n40281) );
  ANDN U42627 ( .B(n40578), .A(n40579), .Z(n40576) );
  AND U42628 ( .A(b[5]), .B(a[45]), .Z(n40575) );
  XOR U42629 ( .A(n40581), .B(n40582), .Z(n40286) );
  ANDN U42630 ( .B(n40583), .A(n40584), .Z(n40581) );
  AND U42631 ( .A(b[4]), .B(a[46]), .Z(n40580) );
  XOR U42632 ( .A(n40586), .B(n40587), .Z(n40291) );
  ANDN U42633 ( .B(n40303), .A(n40304), .Z(n40586) );
  AND U42634 ( .A(b[2]), .B(a[47]), .Z(n40588) );
  XNOR U42635 ( .A(n40583), .B(n40587), .Z(n40589) );
  XOR U42636 ( .A(n40590), .B(n40591), .Z(n40587) );
  OR U42637 ( .A(n40306), .B(n40307), .Z(n40591) );
  XNOR U42638 ( .A(n40593), .B(n40594), .Z(n40592) );
  XOR U42639 ( .A(n40593), .B(n40596), .Z(n40306) );
  NAND U42640 ( .A(b[1]), .B(a[47]), .Z(n40596) );
  IV U42641 ( .A(n40590), .Z(n40593) );
  NANDN U42642 ( .A(n117), .B(n118), .Z(n40590) );
  XOR U42643 ( .A(n40597), .B(n40598), .Z(n118) );
  NAND U42644 ( .A(a[47]), .B(b[0]), .Z(n117) );
  XNOR U42645 ( .A(n40578), .B(n40582), .Z(n40599) );
  XNOR U42646 ( .A(n40573), .B(n40577), .Z(n40600) );
  XNOR U42647 ( .A(n40568), .B(n40572), .Z(n40601) );
  XNOR U42648 ( .A(n40563), .B(n40567), .Z(n40602) );
  XNOR U42649 ( .A(n40558), .B(n40562), .Z(n40603) );
  XNOR U42650 ( .A(n40553), .B(n40557), .Z(n40604) );
  XNOR U42651 ( .A(n40548), .B(n40552), .Z(n40605) );
  XNOR U42652 ( .A(n40543), .B(n40547), .Z(n40606) );
  XNOR U42653 ( .A(n40538), .B(n40542), .Z(n40607) );
  XNOR U42654 ( .A(n40533), .B(n40537), .Z(n40608) );
  XNOR U42655 ( .A(n40528), .B(n40532), .Z(n40609) );
  XNOR U42656 ( .A(n40523), .B(n40527), .Z(n40610) );
  XNOR U42657 ( .A(n40518), .B(n40522), .Z(n40611) );
  XNOR U42658 ( .A(n40513), .B(n40517), .Z(n40612) );
  XNOR U42659 ( .A(n40508), .B(n40512), .Z(n40613) );
  XNOR U42660 ( .A(n40503), .B(n40507), .Z(n40614) );
  XNOR U42661 ( .A(n40498), .B(n40502), .Z(n40615) );
  XNOR U42662 ( .A(n40493), .B(n40497), .Z(n40616) );
  XNOR U42663 ( .A(n40488), .B(n40492), .Z(n40617) );
  XNOR U42664 ( .A(n40483), .B(n40487), .Z(n40618) );
  XNOR U42665 ( .A(n40478), .B(n40482), .Z(n40619) );
  XNOR U42666 ( .A(n40473), .B(n40477), .Z(n40620) );
  XNOR U42667 ( .A(n40468), .B(n40472), .Z(n40621) );
  XNOR U42668 ( .A(n40463), .B(n40467), .Z(n40622) );
  XNOR U42669 ( .A(n40458), .B(n40462), .Z(n40623) );
  XNOR U42670 ( .A(n40453), .B(n40457), .Z(n40624) );
  XNOR U42671 ( .A(n40448), .B(n40452), .Z(n40625) );
  XNOR U42672 ( .A(n40443), .B(n40447), .Z(n40626) );
  XNOR U42673 ( .A(n40438), .B(n40442), .Z(n40627) );
  XNOR U42674 ( .A(n40433), .B(n40437), .Z(n40628) );
  XNOR U42675 ( .A(n40428), .B(n40432), .Z(n40629) );
  XNOR U42676 ( .A(n40423), .B(n40427), .Z(n40630) );
  XNOR U42677 ( .A(n40418), .B(n40422), .Z(n40631) );
  XNOR U42678 ( .A(n40413), .B(n40417), .Z(n40632) );
  XNOR U42679 ( .A(n40408), .B(n40412), .Z(n40633) );
  XNOR U42680 ( .A(n40403), .B(n40407), .Z(n40634) );
  XNOR U42681 ( .A(n40398), .B(n40402), .Z(n40635) );
  XNOR U42682 ( .A(n40393), .B(n40397), .Z(n40636) );
  XNOR U42683 ( .A(n40388), .B(n40392), .Z(n40637) );
  XNOR U42684 ( .A(n40383), .B(n40387), .Z(n40638) );
  XNOR U42685 ( .A(n40378), .B(n40382), .Z(n40639) );
  XNOR U42686 ( .A(n40373), .B(n40377), .Z(n40640) );
  XNOR U42687 ( .A(n40368), .B(n40372), .Z(n40641) );
  XNOR U42688 ( .A(n40363), .B(n40367), .Z(n40642) );
  XNOR U42689 ( .A(n40358), .B(n40362), .Z(n40643) );
  XNOR U42690 ( .A(n40644), .B(n40357), .Z(n40358) );
  AND U42691 ( .A(a[0]), .B(b[49]), .Z(n40644) );
  XOR U42692 ( .A(n40645), .B(n40357), .Z(n40359) );
  XNOR U42693 ( .A(n40646), .B(n40647), .Z(n40357) );
  ANDN U42694 ( .B(n40648), .A(n40649), .Z(n40646) );
  AND U42695 ( .A(a[1]), .B(b[48]), .Z(n40645) );
  XOR U42696 ( .A(n40651), .B(n40652), .Z(n40362) );
  ANDN U42697 ( .B(n40653), .A(n40654), .Z(n40651) );
  AND U42698 ( .A(a[2]), .B(b[47]), .Z(n40650) );
  XOR U42699 ( .A(n40656), .B(n40657), .Z(n40367) );
  ANDN U42700 ( .B(n40658), .A(n40659), .Z(n40656) );
  AND U42701 ( .A(a[3]), .B(b[46]), .Z(n40655) );
  XOR U42702 ( .A(n40661), .B(n40662), .Z(n40372) );
  ANDN U42703 ( .B(n40663), .A(n40664), .Z(n40661) );
  AND U42704 ( .A(a[4]), .B(b[45]), .Z(n40660) );
  XOR U42705 ( .A(n40666), .B(n40667), .Z(n40377) );
  ANDN U42706 ( .B(n40668), .A(n40669), .Z(n40666) );
  AND U42707 ( .A(a[5]), .B(b[44]), .Z(n40665) );
  XOR U42708 ( .A(n40671), .B(n40672), .Z(n40382) );
  ANDN U42709 ( .B(n40673), .A(n40674), .Z(n40671) );
  AND U42710 ( .A(a[6]), .B(b[43]), .Z(n40670) );
  XOR U42711 ( .A(n40676), .B(n40677), .Z(n40387) );
  ANDN U42712 ( .B(n40678), .A(n40679), .Z(n40676) );
  AND U42713 ( .A(a[7]), .B(b[42]), .Z(n40675) );
  XOR U42714 ( .A(n40681), .B(n40682), .Z(n40392) );
  ANDN U42715 ( .B(n40683), .A(n40684), .Z(n40681) );
  AND U42716 ( .A(a[8]), .B(b[41]), .Z(n40680) );
  XOR U42717 ( .A(n40686), .B(n40687), .Z(n40397) );
  ANDN U42718 ( .B(n40688), .A(n40689), .Z(n40686) );
  AND U42719 ( .A(a[9]), .B(b[40]), .Z(n40685) );
  XOR U42720 ( .A(n40691), .B(n40692), .Z(n40402) );
  ANDN U42721 ( .B(n40693), .A(n40694), .Z(n40691) );
  AND U42722 ( .A(a[10]), .B(b[39]), .Z(n40690) );
  XOR U42723 ( .A(n40696), .B(n40697), .Z(n40407) );
  ANDN U42724 ( .B(n40698), .A(n40699), .Z(n40696) );
  AND U42725 ( .A(a[11]), .B(b[38]), .Z(n40695) );
  XOR U42726 ( .A(n40701), .B(n40702), .Z(n40412) );
  ANDN U42727 ( .B(n40703), .A(n40704), .Z(n40701) );
  AND U42728 ( .A(a[12]), .B(b[37]), .Z(n40700) );
  XOR U42729 ( .A(n40706), .B(n40707), .Z(n40417) );
  ANDN U42730 ( .B(n40708), .A(n40709), .Z(n40706) );
  AND U42731 ( .A(a[13]), .B(b[36]), .Z(n40705) );
  XOR U42732 ( .A(n40711), .B(n40712), .Z(n40422) );
  ANDN U42733 ( .B(n40713), .A(n40714), .Z(n40711) );
  AND U42734 ( .A(a[14]), .B(b[35]), .Z(n40710) );
  XOR U42735 ( .A(n40716), .B(n40717), .Z(n40427) );
  ANDN U42736 ( .B(n40718), .A(n40719), .Z(n40716) );
  AND U42737 ( .A(a[15]), .B(b[34]), .Z(n40715) );
  XOR U42738 ( .A(n40721), .B(n40722), .Z(n40432) );
  ANDN U42739 ( .B(n40723), .A(n40724), .Z(n40721) );
  AND U42740 ( .A(a[16]), .B(b[33]), .Z(n40720) );
  XOR U42741 ( .A(n40726), .B(n40727), .Z(n40437) );
  ANDN U42742 ( .B(n40728), .A(n40729), .Z(n40726) );
  AND U42743 ( .A(a[17]), .B(b[32]), .Z(n40725) );
  XOR U42744 ( .A(n40731), .B(n40732), .Z(n40442) );
  ANDN U42745 ( .B(n40733), .A(n40734), .Z(n40731) );
  AND U42746 ( .A(a[18]), .B(b[31]), .Z(n40730) );
  XOR U42747 ( .A(n40736), .B(n40737), .Z(n40447) );
  ANDN U42748 ( .B(n40738), .A(n40739), .Z(n40736) );
  AND U42749 ( .A(a[19]), .B(b[30]), .Z(n40735) );
  XOR U42750 ( .A(n40741), .B(n40742), .Z(n40452) );
  ANDN U42751 ( .B(n40743), .A(n40744), .Z(n40741) );
  AND U42752 ( .A(a[20]), .B(b[29]), .Z(n40740) );
  XOR U42753 ( .A(n40746), .B(n40747), .Z(n40457) );
  ANDN U42754 ( .B(n40748), .A(n40749), .Z(n40746) );
  AND U42755 ( .A(a[21]), .B(b[28]), .Z(n40745) );
  XOR U42756 ( .A(n40751), .B(n40752), .Z(n40462) );
  ANDN U42757 ( .B(n40753), .A(n40754), .Z(n40751) );
  AND U42758 ( .A(a[22]), .B(b[27]), .Z(n40750) );
  XOR U42759 ( .A(n40756), .B(n40757), .Z(n40467) );
  ANDN U42760 ( .B(n40758), .A(n40759), .Z(n40756) );
  AND U42761 ( .A(a[23]), .B(b[26]), .Z(n40755) );
  XOR U42762 ( .A(n40761), .B(n40762), .Z(n40472) );
  ANDN U42763 ( .B(n40763), .A(n40764), .Z(n40761) );
  AND U42764 ( .A(a[24]), .B(b[25]), .Z(n40760) );
  XOR U42765 ( .A(n40766), .B(n40767), .Z(n40477) );
  ANDN U42766 ( .B(n40768), .A(n40769), .Z(n40766) );
  AND U42767 ( .A(a[25]), .B(b[24]), .Z(n40765) );
  XOR U42768 ( .A(n40771), .B(n40772), .Z(n40482) );
  ANDN U42769 ( .B(n40773), .A(n40774), .Z(n40771) );
  AND U42770 ( .A(a[26]), .B(b[23]), .Z(n40770) );
  XOR U42771 ( .A(n40776), .B(n40777), .Z(n40487) );
  ANDN U42772 ( .B(n40778), .A(n40779), .Z(n40776) );
  AND U42773 ( .A(a[27]), .B(b[22]), .Z(n40775) );
  XOR U42774 ( .A(n40781), .B(n40782), .Z(n40492) );
  ANDN U42775 ( .B(n40783), .A(n40784), .Z(n40781) );
  AND U42776 ( .A(a[28]), .B(b[21]), .Z(n40780) );
  XOR U42777 ( .A(n40786), .B(n40787), .Z(n40497) );
  ANDN U42778 ( .B(n40788), .A(n40789), .Z(n40786) );
  AND U42779 ( .A(a[29]), .B(b[20]), .Z(n40785) );
  XOR U42780 ( .A(n40791), .B(n40792), .Z(n40502) );
  ANDN U42781 ( .B(n40793), .A(n40794), .Z(n40791) );
  AND U42782 ( .A(a[30]), .B(b[19]), .Z(n40790) );
  XOR U42783 ( .A(n40796), .B(n40797), .Z(n40507) );
  ANDN U42784 ( .B(n40798), .A(n40799), .Z(n40796) );
  AND U42785 ( .A(a[31]), .B(b[18]), .Z(n40795) );
  XOR U42786 ( .A(n40801), .B(n40802), .Z(n40512) );
  ANDN U42787 ( .B(n40803), .A(n40804), .Z(n40801) );
  AND U42788 ( .A(a[32]), .B(b[17]), .Z(n40800) );
  XOR U42789 ( .A(n40806), .B(n40807), .Z(n40517) );
  ANDN U42790 ( .B(n40808), .A(n40809), .Z(n40806) );
  AND U42791 ( .A(a[33]), .B(b[16]), .Z(n40805) );
  XOR U42792 ( .A(n40811), .B(n40812), .Z(n40522) );
  ANDN U42793 ( .B(n40813), .A(n40814), .Z(n40811) );
  AND U42794 ( .A(a[34]), .B(b[15]), .Z(n40810) );
  XOR U42795 ( .A(n40816), .B(n40817), .Z(n40527) );
  ANDN U42796 ( .B(n40818), .A(n40819), .Z(n40816) );
  AND U42797 ( .A(a[35]), .B(b[14]), .Z(n40815) );
  XOR U42798 ( .A(n40821), .B(n40822), .Z(n40532) );
  ANDN U42799 ( .B(n40823), .A(n40824), .Z(n40821) );
  AND U42800 ( .A(a[36]), .B(b[13]), .Z(n40820) );
  XOR U42801 ( .A(n40826), .B(n40827), .Z(n40537) );
  ANDN U42802 ( .B(n40828), .A(n40829), .Z(n40826) );
  AND U42803 ( .A(a[37]), .B(b[12]), .Z(n40825) );
  XOR U42804 ( .A(n40831), .B(n40832), .Z(n40542) );
  ANDN U42805 ( .B(n40833), .A(n40834), .Z(n40831) );
  AND U42806 ( .A(a[38]), .B(b[11]), .Z(n40830) );
  XOR U42807 ( .A(n40836), .B(n40837), .Z(n40547) );
  ANDN U42808 ( .B(n40838), .A(n40839), .Z(n40836) );
  AND U42809 ( .A(a[39]), .B(b[10]), .Z(n40835) );
  XOR U42810 ( .A(n40841), .B(n40842), .Z(n40552) );
  ANDN U42811 ( .B(n40843), .A(n40844), .Z(n40841) );
  AND U42812 ( .A(b[9]), .B(a[40]), .Z(n40840) );
  XOR U42813 ( .A(n40846), .B(n40847), .Z(n40557) );
  ANDN U42814 ( .B(n40848), .A(n40849), .Z(n40846) );
  AND U42815 ( .A(b[8]), .B(a[41]), .Z(n40845) );
  XOR U42816 ( .A(n40851), .B(n40852), .Z(n40562) );
  ANDN U42817 ( .B(n40853), .A(n40854), .Z(n40851) );
  AND U42818 ( .A(b[7]), .B(a[42]), .Z(n40850) );
  XOR U42819 ( .A(n40856), .B(n40857), .Z(n40567) );
  ANDN U42820 ( .B(n40858), .A(n40859), .Z(n40856) );
  AND U42821 ( .A(b[6]), .B(a[43]), .Z(n40855) );
  XOR U42822 ( .A(n40861), .B(n40862), .Z(n40572) );
  ANDN U42823 ( .B(n40863), .A(n40864), .Z(n40861) );
  AND U42824 ( .A(b[5]), .B(a[44]), .Z(n40860) );
  XOR U42825 ( .A(n40866), .B(n40867), .Z(n40577) );
  ANDN U42826 ( .B(n40868), .A(n40869), .Z(n40866) );
  AND U42827 ( .A(b[4]), .B(a[45]), .Z(n40865) );
  XOR U42828 ( .A(n40871), .B(n40872), .Z(n40582) );
  ANDN U42829 ( .B(n40594), .A(n40595), .Z(n40871) );
  AND U42830 ( .A(b[2]), .B(a[46]), .Z(n40873) );
  XNOR U42831 ( .A(n40868), .B(n40872), .Z(n40874) );
  XOR U42832 ( .A(n40875), .B(n40876), .Z(n40872) );
  OR U42833 ( .A(n40597), .B(n40598), .Z(n40876) );
  XNOR U42834 ( .A(n40878), .B(n40879), .Z(n40877) );
  XOR U42835 ( .A(n40878), .B(n40881), .Z(n40597) );
  NAND U42836 ( .A(b[1]), .B(a[46]), .Z(n40881) );
  IV U42837 ( .A(n40875), .Z(n40878) );
  NANDN U42838 ( .A(n119), .B(n120), .Z(n40875) );
  XOR U42839 ( .A(n40882), .B(n40883), .Z(n120) );
  NAND U42840 ( .A(a[46]), .B(b[0]), .Z(n119) );
  XNOR U42841 ( .A(n40863), .B(n40867), .Z(n40884) );
  XNOR U42842 ( .A(n40858), .B(n40862), .Z(n40885) );
  XNOR U42843 ( .A(n40853), .B(n40857), .Z(n40886) );
  XNOR U42844 ( .A(n40848), .B(n40852), .Z(n40887) );
  XNOR U42845 ( .A(n40843), .B(n40847), .Z(n40888) );
  XNOR U42846 ( .A(n40838), .B(n40842), .Z(n40889) );
  XNOR U42847 ( .A(n40833), .B(n40837), .Z(n40890) );
  XNOR U42848 ( .A(n40828), .B(n40832), .Z(n40891) );
  XNOR U42849 ( .A(n40823), .B(n40827), .Z(n40892) );
  XNOR U42850 ( .A(n40818), .B(n40822), .Z(n40893) );
  XNOR U42851 ( .A(n40813), .B(n40817), .Z(n40894) );
  XNOR U42852 ( .A(n40808), .B(n40812), .Z(n40895) );
  XNOR U42853 ( .A(n40803), .B(n40807), .Z(n40896) );
  XNOR U42854 ( .A(n40798), .B(n40802), .Z(n40897) );
  XNOR U42855 ( .A(n40793), .B(n40797), .Z(n40898) );
  XNOR U42856 ( .A(n40788), .B(n40792), .Z(n40899) );
  XNOR U42857 ( .A(n40783), .B(n40787), .Z(n40900) );
  XNOR U42858 ( .A(n40778), .B(n40782), .Z(n40901) );
  XNOR U42859 ( .A(n40773), .B(n40777), .Z(n40902) );
  XNOR U42860 ( .A(n40768), .B(n40772), .Z(n40903) );
  XNOR U42861 ( .A(n40763), .B(n40767), .Z(n40904) );
  XNOR U42862 ( .A(n40758), .B(n40762), .Z(n40905) );
  XNOR U42863 ( .A(n40753), .B(n40757), .Z(n40906) );
  XNOR U42864 ( .A(n40748), .B(n40752), .Z(n40907) );
  XNOR U42865 ( .A(n40743), .B(n40747), .Z(n40908) );
  XNOR U42866 ( .A(n40738), .B(n40742), .Z(n40909) );
  XNOR U42867 ( .A(n40733), .B(n40737), .Z(n40910) );
  XNOR U42868 ( .A(n40728), .B(n40732), .Z(n40911) );
  XNOR U42869 ( .A(n40723), .B(n40727), .Z(n40912) );
  XNOR U42870 ( .A(n40718), .B(n40722), .Z(n40913) );
  XNOR U42871 ( .A(n40713), .B(n40717), .Z(n40914) );
  XNOR U42872 ( .A(n40708), .B(n40712), .Z(n40915) );
  XNOR U42873 ( .A(n40703), .B(n40707), .Z(n40916) );
  XNOR U42874 ( .A(n40698), .B(n40702), .Z(n40917) );
  XNOR U42875 ( .A(n40693), .B(n40697), .Z(n40918) );
  XNOR U42876 ( .A(n40688), .B(n40692), .Z(n40919) );
  XNOR U42877 ( .A(n40683), .B(n40687), .Z(n40920) );
  XNOR U42878 ( .A(n40678), .B(n40682), .Z(n40921) );
  XNOR U42879 ( .A(n40673), .B(n40677), .Z(n40922) );
  XNOR U42880 ( .A(n40668), .B(n40672), .Z(n40923) );
  XNOR U42881 ( .A(n40663), .B(n40667), .Z(n40924) );
  XNOR U42882 ( .A(n40658), .B(n40662), .Z(n40925) );
  XNOR U42883 ( .A(n40653), .B(n40657), .Z(n40926) );
  XNOR U42884 ( .A(n40648), .B(n40652), .Z(n40927) );
  XOR U42885 ( .A(n40928), .B(n40647), .Z(n40648) );
  AND U42886 ( .A(a[0]), .B(b[48]), .Z(n40928) );
  XNOR U42887 ( .A(n40929), .B(n40647), .Z(n40649) );
  XNOR U42888 ( .A(n40930), .B(n40931), .Z(n40647) );
  ANDN U42889 ( .B(n40932), .A(n40933), .Z(n40930) );
  AND U42890 ( .A(a[1]), .B(b[47]), .Z(n40929) );
  XOR U42891 ( .A(n40935), .B(n40936), .Z(n40652) );
  ANDN U42892 ( .B(n40937), .A(n40938), .Z(n40935) );
  AND U42893 ( .A(a[2]), .B(b[46]), .Z(n40934) );
  XOR U42894 ( .A(n40940), .B(n40941), .Z(n40657) );
  ANDN U42895 ( .B(n40942), .A(n40943), .Z(n40940) );
  AND U42896 ( .A(a[3]), .B(b[45]), .Z(n40939) );
  XOR U42897 ( .A(n40945), .B(n40946), .Z(n40662) );
  ANDN U42898 ( .B(n40947), .A(n40948), .Z(n40945) );
  AND U42899 ( .A(a[4]), .B(b[44]), .Z(n40944) );
  XOR U42900 ( .A(n40950), .B(n40951), .Z(n40667) );
  ANDN U42901 ( .B(n40952), .A(n40953), .Z(n40950) );
  AND U42902 ( .A(a[5]), .B(b[43]), .Z(n40949) );
  XOR U42903 ( .A(n40955), .B(n40956), .Z(n40672) );
  ANDN U42904 ( .B(n40957), .A(n40958), .Z(n40955) );
  AND U42905 ( .A(a[6]), .B(b[42]), .Z(n40954) );
  XOR U42906 ( .A(n40960), .B(n40961), .Z(n40677) );
  ANDN U42907 ( .B(n40962), .A(n40963), .Z(n40960) );
  AND U42908 ( .A(a[7]), .B(b[41]), .Z(n40959) );
  XOR U42909 ( .A(n40965), .B(n40966), .Z(n40682) );
  ANDN U42910 ( .B(n40967), .A(n40968), .Z(n40965) );
  AND U42911 ( .A(a[8]), .B(b[40]), .Z(n40964) );
  XOR U42912 ( .A(n40970), .B(n40971), .Z(n40687) );
  ANDN U42913 ( .B(n40972), .A(n40973), .Z(n40970) );
  AND U42914 ( .A(a[9]), .B(b[39]), .Z(n40969) );
  XOR U42915 ( .A(n40975), .B(n40976), .Z(n40692) );
  ANDN U42916 ( .B(n40977), .A(n40978), .Z(n40975) );
  AND U42917 ( .A(a[10]), .B(b[38]), .Z(n40974) );
  XOR U42918 ( .A(n40980), .B(n40981), .Z(n40697) );
  ANDN U42919 ( .B(n40982), .A(n40983), .Z(n40980) );
  AND U42920 ( .A(a[11]), .B(b[37]), .Z(n40979) );
  XOR U42921 ( .A(n40985), .B(n40986), .Z(n40702) );
  ANDN U42922 ( .B(n40987), .A(n40988), .Z(n40985) );
  AND U42923 ( .A(a[12]), .B(b[36]), .Z(n40984) );
  XOR U42924 ( .A(n40990), .B(n40991), .Z(n40707) );
  ANDN U42925 ( .B(n40992), .A(n40993), .Z(n40990) );
  AND U42926 ( .A(a[13]), .B(b[35]), .Z(n40989) );
  XOR U42927 ( .A(n40995), .B(n40996), .Z(n40712) );
  ANDN U42928 ( .B(n40997), .A(n40998), .Z(n40995) );
  AND U42929 ( .A(a[14]), .B(b[34]), .Z(n40994) );
  XOR U42930 ( .A(n41000), .B(n41001), .Z(n40717) );
  ANDN U42931 ( .B(n41002), .A(n41003), .Z(n41000) );
  AND U42932 ( .A(a[15]), .B(b[33]), .Z(n40999) );
  XOR U42933 ( .A(n41005), .B(n41006), .Z(n40722) );
  ANDN U42934 ( .B(n41007), .A(n41008), .Z(n41005) );
  AND U42935 ( .A(a[16]), .B(b[32]), .Z(n41004) );
  XOR U42936 ( .A(n41010), .B(n41011), .Z(n40727) );
  ANDN U42937 ( .B(n41012), .A(n41013), .Z(n41010) );
  AND U42938 ( .A(a[17]), .B(b[31]), .Z(n41009) );
  XOR U42939 ( .A(n41015), .B(n41016), .Z(n40732) );
  ANDN U42940 ( .B(n41017), .A(n41018), .Z(n41015) );
  AND U42941 ( .A(a[18]), .B(b[30]), .Z(n41014) );
  XOR U42942 ( .A(n41020), .B(n41021), .Z(n40737) );
  ANDN U42943 ( .B(n41022), .A(n41023), .Z(n41020) );
  AND U42944 ( .A(a[19]), .B(b[29]), .Z(n41019) );
  XOR U42945 ( .A(n41025), .B(n41026), .Z(n40742) );
  ANDN U42946 ( .B(n41027), .A(n41028), .Z(n41025) );
  AND U42947 ( .A(a[20]), .B(b[28]), .Z(n41024) );
  XOR U42948 ( .A(n41030), .B(n41031), .Z(n40747) );
  ANDN U42949 ( .B(n41032), .A(n41033), .Z(n41030) );
  AND U42950 ( .A(a[21]), .B(b[27]), .Z(n41029) );
  XOR U42951 ( .A(n41035), .B(n41036), .Z(n40752) );
  ANDN U42952 ( .B(n41037), .A(n41038), .Z(n41035) );
  AND U42953 ( .A(a[22]), .B(b[26]), .Z(n41034) );
  XOR U42954 ( .A(n41040), .B(n41041), .Z(n40757) );
  ANDN U42955 ( .B(n41042), .A(n41043), .Z(n41040) );
  AND U42956 ( .A(a[23]), .B(b[25]), .Z(n41039) );
  XOR U42957 ( .A(n41045), .B(n41046), .Z(n40762) );
  ANDN U42958 ( .B(n41047), .A(n41048), .Z(n41045) );
  AND U42959 ( .A(a[24]), .B(b[24]), .Z(n41044) );
  XOR U42960 ( .A(n41050), .B(n41051), .Z(n40767) );
  ANDN U42961 ( .B(n41052), .A(n41053), .Z(n41050) );
  AND U42962 ( .A(a[25]), .B(b[23]), .Z(n41049) );
  XOR U42963 ( .A(n41055), .B(n41056), .Z(n40772) );
  ANDN U42964 ( .B(n41057), .A(n41058), .Z(n41055) );
  AND U42965 ( .A(a[26]), .B(b[22]), .Z(n41054) );
  XOR U42966 ( .A(n41060), .B(n41061), .Z(n40777) );
  ANDN U42967 ( .B(n41062), .A(n41063), .Z(n41060) );
  AND U42968 ( .A(a[27]), .B(b[21]), .Z(n41059) );
  XOR U42969 ( .A(n41065), .B(n41066), .Z(n40782) );
  ANDN U42970 ( .B(n41067), .A(n41068), .Z(n41065) );
  AND U42971 ( .A(a[28]), .B(b[20]), .Z(n41064) );
  XOR U42972 ( .A(n41070), .B(n41071), .Z(n40787) );
  ANDN U42973 ( .B(n41072), .A(n41073), .Z(n41070) );
  AND U42974 ( .A(a[29]), .B(b[19]), .Z(n41069) );
  XOR U42975 ( .A(n41075), .B(n41076), .Z(n40792) );
  ANDN U42976 ( .B(n41077), .A(n41078), .Z(n41075) );
  AND U42977 ( .A(a[30]), .B(b[18]), .Z(n41074) );
  XOR U42978 ( .A(n41080), .B(n41081), .Z(n40797) );
  ANDN U42979 ( .B(n41082), .A(n41083), .Z(n41080) );
  AND U42980 ( .A(a[31]), .B(b[17]), .Z(n41079) );
  XOR U42981 ( .A(n41085), .B(n41086), .Z(n40802) );
  ANDN U42982 ( .B(n41087), .A(n41088), .Z(n41085) );
  AND U42983 ( .A(a[32]), .B(b[16]), .Z(n41084) );
  XOR U42984 ( .A(n41090), .B(n41091), .Z(n40807) );
  ANDN U42985 ( .B(n41092), .A(n41093), .Z(n41090) );
  AND U42986 ( .A(a[33]), .B(b[15]), .Z(n41089) );
  XOR U42987 ( .A(n41095), .B(n41096), .Z(n40812) );
  ANDN U42988 ( .B(n41097), .A(n41098), .Z(n41095) );
  AND U42989 ( .A(a[34]), .B(b[14]), .Z(n41094) );
  XOR U42990 ( .A(n41100), .B(n41101), .Z(n40817) );
  ANDN U42991 ( .B(n41102), .A(n41103), .Z(n41100) );
  AND U42992 ( .A(a[35]), .B(b[13]), .Z(n41099) );
  XOR U42993 ( .A(n41105), .B(n41106), .Z(n40822) );
  ANDN U42994 ( .B(n41107), .A(n41108), .Z(n41105) );
  AND U42995 ( .A(a[36]), .B(b[12]), .Z(n41104) );
  XOR U42996 ( .A(n41110), .B(n41111), .Z(n40827) );
  ANDN U42997 ( .B(n41112), .A(n41113), .Z(n41110) );
  AND U42998 ( .A(a[37]), .B(b[11]), .Z(n41109) );
  XOR U42999 ( .A(n41115), .B(n41116), .Z(n40832) );
  ANDN U43000 ( .B(n41117), .A(n41118), .Z(n41115) );
  AND U43001 ( .A(a[38]), .B(b[10]), .Z(n41114) );
  XOR U43002 ( .A(n41120), .B(n41121), .Z(n40837) );
  ANDN U43003 ( .B(n41122), .A(n41123), .Z(n41120) );
  AND U43004 ( .A(b[9]), .B(a[39]), .Z(n41119) );
  XOR U43005 ( .A(n41125), .B(n41126), .Z(n40842) );
  ANDN U43006 ( .B(n41127), .A(n41128), .Z(n41125) );
  AND U43007 ( .A(b[8]), .B(a[40]), .Z(n41124) );
  XOR U43008 ( .A(n41130), .B(n41131), .Z(n40847) );
  ANDN U43009 ( .B(n41132), .A(n41133), .Z(n41130) );
  AND U43010 ( .A(b[7]), .B(a[41]), .Z(n41129) );
  XOR U43011 ( .A(n41135), .B(n41136), .Z(n40852) );
  ANDN U43012 ( .B(n41137), .A(n41138), .Z(n41135) );
  AND U43013 ( .A(b[6]), .B(a[42]), .Z(n41134) );
  XOR U43014 ( .A(n41140), .B(n41141), .Z(n40857) );
  ANDN U43015 ( .B(n41142), .A(n41143), .Z(n41140) );
  AND U43016 ( .A(b[5]), .B(a[43]), .Z(n41139) );
  XOR U43017 ( .A(n41145), .B(n41146), .Z(n40862) );
  ANDN U43018 ( .B(n41147), .A(n41148), .Z(n41145) );
  AND U43019 ( .A(b[4]), .B(a[44]), .Z(n41144) );
  XOR U43020 ( .A(n41150), .B(n41151), .Z(n40867) );
  ANDN U43021 ( .B(n40879), .A(n40880), .Z(n41150) );
  AND U43022 ( .A(b[2]), .B(a[45]), .Z(n41152) );
  XNOR U43023 ( .A(n41147), .B(n41151), .Z(n41153) );
  XOR U43024 ( .A(n41154), .B(n41155), .Z(n41151) );
  OR U43025 ( .A(n40882), .B(n40883), .Z(n41155) );
  XNOR U43026 ( .A(n41157), .B(n41158), .Z(n41156) );
  XOR U43027 ( .A(n41157), .B(n41160), .Z(n40882) );
  NAND U43028 ( .A(b[1]), .B(a[45]), .Z(n41160) );
  IV U43029 ( .A(n41154), .Z(n41157) );
  NANDN U43030 ( .A(n121), .B(n122), .Z(n41154) );
  XOR U43031 ( .A(n41161), .B(n41162), .Z(n122) );
  NAND U43032 ( .A(a[45]), .B(b[0]), .Z(n121) );
  XNOR U43033 ( .A(n41142), .B(n41146), .Z(n41163) );
  XNOR U43034 ( .A(n41137), .B(n41141), .Z(n41164) );
  XNOR U43035 ( .A(n41132), .B(n41136), .Z(n41165) );
  XNOR U43036 ( .A(n41127), .B(n41131), .Z(n41166) );
  XNOR U43037 ( .A(n41122), .B(n41126), .Z(n41167) );
  XNOR U43038 ( .A(n41117), .B(n41121), .Z(n41168) );
  XNOR U43039 ( .A(n41112), .B(n41116), .Z(n41169) );
  XNOR U43040 ( .A(n41107), .B(n41111), .Z(n41170) );
  XNOR U43041 ( .A(n41102), .B(n41106), .Z(n41171) );
  XNOR U43042 ( .A(n41097), .B(n41101), .Z(n41172) );
  XNOR U43043 ( .A(n41092), .B(n41096), .Z(n41173) );
  XNOR U43044 ( .A(n41087), .B(n41091), .Z(n41174) );
  XNOR U43045 ( .A(n41082), .B(n41086), .Z(n41175) );
  XNOR U43046 ( .A(n41077), .B(n41081), .Z(n41176) );
  XNOR U43047 ( .A(n41072), .B(n41076), .Z(n41177) );
  XNOR U43048 ( .A(n41067), .B(n41071), .Z(n41178) );
  XNOR U43049 ( .A(n41062), .B(n41066), .Z(n41179) );
  XNOR U43050 ( .A(n41057), .B(n41061), .Z(n41180) );
  XNOR U43051 ( .A(n41052), .B(n41056), .Z(n41181) );
  XNOR U43052 ( .A(n41047), .B(n41051), .Z(n41182) );
  XNOR U43053 ( .A(n41042), .B(n41046), .Z(n41183) );
  XNOR U43054 ( .A(n41037), .B(n41041), .Z(n41184) );
  XNOR U43055 ( .A(n41032), .B(n41036), .Z(n41185) );
  XNOR U43056 ( .A(n41027), .B(n41031), .Z(n41186) );
  XNOR U43057 ( .A(n41022), .B(n41026), .Z(n41187) );
  XNOR U43058 ( .A(n41017), .B(n41021), .Z(n41188) );
  XNOR U43059 ( .A(n41012), .B(n41016), .Z(n41189) );
  XNOR U43060 ( .A(n41007), .B(n41011), .Z(n41190) );
  XNOR U43061 ( .A(n41002), .B(n41006), .Z(n41191) );
  XNOR U43062 ( .A(n40997), .B(n41001), .Z(n41192) );
  XNOR U43063 ( .A(n40992), .B(n40996), .Z(n41193) );
  XNOR U43064 ( .A(n40987), .B(n40991), .Z(n41194) );
  XNOR U43065 ( .A(n40982), .B(n40986), .Z(n41195) );
  XNOR U43066 ( .A(n40977), .B(n40981), .Z(n41196) );
  XNOR U43067 ( .A(n40972), .B(n40976), .Z(n41197) );
  XNOR U43068 ( .A(n40967), .B(n40971), .Z(n41198) );
  XNOR U43069 ( .A(n40962), .B(n40966), .Z(n41199) );
  XNOR U43070 ( .A(n40957), .B(n40961), .Z(n41200) );
  XNOR U43071 ( .A(n40952), .B(n40956), .Z(n41201) );
  XNOR U43072 ( .A(n40947), .B(n40951), .Z(n41202) );
  XNOR U43073 ( .A(n40942), .B(n40946), .Z(n41203) );
  XNOR U43074 ( .A(n40937), .B(n40941), .Z(n41204) );
  XNOR U43075 ( .A(n40932), .B(n40936), .Z(n41205) );
  XNOR U43076 ( .A(n41206), .B(n40931), .Z(n40932) );
  AND U43077 ( .A(a[0]), .B(b[47]), .Z(n41206) );
  XOR U43078 ( .A(n41207), .B(n40931), .Z(n40933) );
  XNOR U43079 ( .A(n41208), .B(n41209), .Z(n40931) );
  ANDN U43080 ( .B(n41210), .A(n41211), .Z(n41208) );
  AND U43081 ( .A(a[1]), .B(b[46]), .Z(n41207) );
  XOR U43082 ( .A(n41213), .B(n41214), .Z(n40936) );
  ANDN U43083 ( .B(n41215), .A(n41216), .Z(n41213) );
  AND U43084 ( .A(a[2]), .B(b[45]), .Z(n41212) );
  XOR U43085 ( .A(n41218), .B(n41219), .Z(n40941) );
  ANDN U43086 ( .B(n41220), .A(n41221), .Z(n41218) );
  AND U43087 ( .A(a[3]), .B(b[44]), .Z(n41217) );
  XOR U43088 ( .A(n41223), .B(n41224), .Z(n40946) );
  ANDN U43089 ( .B(n41225), .A(n41226), .Z(n41223) );
  AND U43090 ( .A(a[4]), .B(b[43]), .Z(n41222) );
  XOR U43091 ( .A(n41228), .B(n41229), .Z(n40951) );
  ANDN U43092 ( .B(n41230), .A(n41231), .Z(n41228) );
  AND U43093 ( .A(a[5]), .B(b[42]), .Z(n41227) );
  XOR U43094 ( .A(n41233), .B(n41234), .Z(n40956) );
  ANDN U43095 ( .B(n41235), .A(n41236), .Z(n41233) );
  AND U43096 ( .A(a[6]), .B(b[41]), .Z(n41232) );
  XOR U43097 ( .A(n41238), .B(n41239), .Z(n40961) );
  ANDN U43098 ( .B(n41240), .A(n41241), .Z(n41238) );
  AND U43099 ( .A(a[7]), .B(b[40]), .Z(n41237) );
  XOR U43100 ( .A(n41243), .B(n41244), .Z(n40966) );
  ANDN U43101 ( .B(n41245), .A(n41246), .Z(n41243) );
  AND U43102 ( .A(a[8]), .B(b[39]), .Z(n41242) );
  XOR U43103 ( .A(n41248), .B(n41249), .Z(n40971) );
  ANDN U43104 ( .B(n41250), .A(n41251), .Z(n41248) );
  AND U43105 ( .A(a[9]), .B(b[38]), .Z(n41247) );
  XOR U43106 ( .A(n41253), .B(n41254), .Z(n40976) );
  ANDN U43107 ( .B(n41255), .A(n41256), .Z(n41253) );
  AND U43108 ( .A(a[10]), .B(b[37]), .Z(n41252) );
  XOR U43109 ( .A(n41258), .B(n41259), .Z(n40981) );
  ANDN U43110 ( .B(n41260), .A(n41261), .Z(n41258) );
  AND U43111 ( .A(a[11]), .B(b[36]), .Z(n41257) );
  XOR U43112 ( .A(n41263), .B(n41264), .Z(n40986) );
  ANDN U43113 ( .B(n41265), .A(n41266), .Z(n41263) );
  AND U43114 ( .A(a[12]), .B(b[35]), .Z(n41262) );
  XOR U43115 ( .A(n41268), .B(n41269), .Z(n40991) );
  ANDN U43116 ( .B(n41270), .A(n41271), .Z(n41268) );
  AND U43117 ( .A(a[13]), .B(b[34]), .Z(n41267) );
  XOR U43118 ( .A(n41273), .B(n41274), .Z(n40996) );
  ANDN U43119 ( .B(n41275), .A(n41276), .Z(n41273) );
  AND U43120 ( .A(a[14]), .B(b[33]), .Z(n41272) );
  XOR U43121 ( .A(n41278), .B(n41279), .Z(n41001) );
  ANDN U43122 ( .B(n41280), .A(n41281), .Z(n41278) );
  AND U43123 ( .A(a[15]), .B(b[32]), .Z(n41277) );
  XOR U43124 ( .A(n41283), .B(n41284), .Z(n41006) );
  ANDN U43125 ( .B(n41285), .A(n41286), .Z(n41283) );
  AND U43126 ( .A(a[16]), .B(b[31]), .Z(n41282) );
  XOR U43127 ( .A(n41288), .B(n41289), .Z(n41011) );
  ANDN U43128 ( .B(n41290), .A(n41291), .Z(n41288) );
  AND U43129 ( .A(a[17]), .B(b[30]), .Z(n41287) );
  XOR U43130 ( .A(n41293), .B(n41294), .Z(n41016) );
  ANDN U43131 ( .B(n41295), .A(n41296), .Z(n41293) );
  AND U43132 ( .A(a[18]), .B(b[29]), .Z(n41292) );
  XOR U43133 ( .A(n41298), .B(n41299), .Z(n41021) );
  ANDN U43134 ( .B(n41300), .A(n41301), .Z(n41298) );
  AND U43135 ( .A(a[19]), .B(b[28]), .Z(n41297) );
  XOR U43136 ( .A(n41303), .B(n41304), .Z(n41026) );
  ANDN U43137 ( .B(n41305), .A(n41306), .Z(n41303) );
  AND U43138 ( .A(a[20]), .B(b[27]), .Z(n41302) );
  XOR U43139 ( .A(n41308), .B(n41309), .Z(n41031) );
  ANDN U43140 ( .B(n41310), .A(n41311), .Z(n41308) );
  AND U43141 ( .A(a[21]), .B(b[26]), .Z(n41307) );
  XOR U43142 ( .A(n41313), .B(n41314), .Z(n41036) );
  ANDN U43143 ( .B(n41315), .A(n41316), .Z(n41313) );
  AND U43144 ( .A(a[22]), .B(b[25]), .Z(n41312) );
  XOR U43145 ( .A(n41318), .B(n41319), .Z(n41041) );
  ANDN U43146 ( .B(n41320), .A(n41321), .Z(n41318) );
  AND U43147 ( .A(a[23]), .B(b[24]), .Z(n41317) );
  XOR U43148 ( .A(n41323), .B(n41324), .Z(n41046) );
  ANDN U43149 ( .B(n41325), .A(n41326), .Z(n41323) );
  AND U43150 ( .A(a[24]), .B(b[23]), .Z(n41322) );
  XOR U43151 ( .A(n41328), .B(n41329), .Z(n41051) );
  ANDN U43152 ( .B(n41330), .A(n41331), .Z(n41328) );
  AND U43153 ( .A(a[25]), .B(b[22]), .Z(n41327) );
  XOR U43154 ( .A(n41333), .B(n41334), .Z(n41056) );
  ANDN U43155 ( .B(n41335), .A(n41336), .Z(n41333) );
  AND U43156 ( .A(a[26]), .B(b[21]), .Z(n41332) );
  XOR U43157 ( .A(n41338), .B(n41339), .Z(n41061) );
  ANDN U43158 ( .B(n41340), .A(n41341), .Z(n41338) );
  AND U43159 ( .A(a[27]), .B(b[20]), .Z(n41337) );
  XOR U43160 ( .A(n41343), .B(n41344), .Z(n41066) );
  ANDN U43161 ( .B(n41345), .A(n41346), .Z(n41343) );
  AND U43162 ( .A(a[28]), .B(b[19]), .Z(n41342) );
  XOR U43163 ( .A(n41348), .B(n41349), .Z(n41071) );
  ANDN U43164 ( .B(n41350), .A(n41351), .Z(n41348) );
  AND U43165 ( .A(a[29]), .B(b[18]), .Z(n41347) );
  XOR U43166 ( .A(n41353), .B(n41354), .Z(n41076) );
  ANDN U43167 ( .B(n41355), .A(n41356), .Z(n41353) );
  AND U43168 ( .A(a[30]), .B(b[17]), .Z(n41352) );
  XOR U43169 ( .A(n41358), .B(n41359), .Z(n41081) );
  ANDN U43170 ( .B(n41360), .A(n41361), .Z(n41358) );
  AND U43171 ( .A(a[31]), .B(b[16]), .Z(n41357) );
  XOR U43172 ( .A(n41363), .B(n41364), .Z(n41086) );
  ANDN U43173 ( .B(n41365), .A(n41366), .Z(n41363) );
  AND U43174 ( .A(a[32]), .B(b[15]), .Z(n41362) );
  XOR U43175 ( .A(n41368), .B(n41369), .Z(n41091) );
  ANDN U43176 ( .B(n41370), .A(n41371), .Z(n41368) );
  AND U43177 ( .A(a[33]), .B(b[14]), .Z(n41367) );
  XOR U43178 ( .A(n41373), .B(n41374), .Z(n41096) );
  ANDN U43179 ( .B(n41375), .A(n41376), .Z(n41373) );
  AND U43180 ( .A(a[34]), .B(b[13]), .Z(n41372) );
  XOR U43181 ( .A(n41378), .B(n41379), .Z(n41101) );
  ANDN U43182 ( .B(n41380), .A(n41381), .Z(n41378) );
  AND U43183 ( .A(a[35]), .B(b[12]), .Z(n41377) );
  XOR U43184 ( .A(n41383), .B(n41384), .Z(n41106) );
  ANDN U43185 ( .B(n41385), .A(n41386), .Z(n41383) );
  AND U43186 ( .A(a[36]), .B(b[11]), .Z(n41382) );
  XOR U43187 ( .A(n41388), .B(n41389), .Z(n41111) );
  ANDN U43188 ( .B(n41390), .A(n41391), .Z(n41388) );
  AND U43189 ( .A(a[37]), .B(b[10]), .Z(n41387) );
  XOR U43190 ( .A(n41393), .B(n41394), .Z(n41116) );
  ANDN U43191 ( .B(n41395), .A(n41396), .Z(n41393) );
  AND U43192 ( .A(b[9]), .B(a[38]), .Z(n41392) );
  XOR U43193 ( .A(n41398), .B(n41399), .Z(n41121) );
  ANDN U43194 ( .B(n41400), .A(n41401), .Z(n41398) );
  AND U43195 ( .A(b[8]), .B(a[39]), .Z(n41397) );
  XOR U43196 ( .A(n41403), .B(n41404), .Z(n41126) );
  ANDN U43197 ( .B(n41405), .A(n41406), .Z(n41403) );
  AND U43198 ( .A(b[7]), .B(a[40]), .Z(n41402) );
  XOR U43199 ( .A(n41408), .B(n41409), .Z(n41131) );
  ANDN U43200 ( .B(n41410), .A(n41411), .Z(n41408) );
  AND U43201 ( .A(b[6]), .B(a[41]), .Z(n41407) );
  XOR U43202 ( .A(n41413), .B(n41414), .Z(n41136) );
  ANDN U43203 ( .B(n41415), .A(n41416), .Z(n41413) );
  AND U43204 ( .A(b[5]), .B(a[42]), .Z(n41412) );
  XOR U43205 ( .A(n41418), .B(n41419), .Z(n41141) );
  ANDN U43206 ( .B(n41420), .A(n41421), .Z(n41418) );
  AND U43207 ( .A(b[4]), .B(a[43]), .Z(n41417) );
  XOR U43208 ( .A(n41423), .B(n41424), .Z(n41146) );
  ANDN U43209 ( .B(n41158), .A(n41159), .Z(n41423) );
  AND U43210 ( .A(b[2]), .B(a[44]), .Z(n41425) );
  XNOR U43211 ( .A(n41420), .B(n41424), .Z(n41426) );
  XOR U43212 ( .A(n41427), .B(n41428), .Z(n41424) );
  OR U43213 ( .A(n41161), .B(n41162), .Z(n41428) );
  XNOR U43214 ( .A(n41430), .B(n41431), .Z(n41429) );
  XOR U43215 ( .A(n41430), .B(n41433), .Z(n41161) );
  NAND U43216 ( .A(b[1]), .B(a[44]), .Z(n41433) );
  IV U43217 ( .A(n41427), .Z(n41430) );
  NANDN U43218 ( .A(n123), .B(n124), .Z(n41427) );
  XOR U43219 ( .A(n41434), .B(n41435), .Z(n124) );
  NAND U43220 ( .A(a[44]), .B(b[0]), .Z(n123) );
  XNOR U43221 ( .A(n41415), .B(n41419), .Z(n41436) );
  XNOR U43222 ( .A(n41410), .B(n41414), .Z(n41437) );
  XNOR U43223 ( .A(n41405), .B(n41409), .Z(n41438) );
  XNOR U43224 ( .A(n41400), .B(n41404), .Z(n41439) );
  XNOR U43225 ( .A(n41395), .B(n41399), .Z(n41440) );
  XNOR U43226 ( .A(n41390), .B(n41394), .Z(n41441) );
  XNOR U43227 ( .A(n41385), .B(n41389), .Z(n41442) );
  XNOR U43228 ( .A(n41380), .B(n41384), .Z(n41443) );
  XNOR U43229 ( .A(n41375), .B(n41379), .Z(n41444) );
  XNOR U43230 ( .A(n41370), .B(n41374), .Z(n41445) );
  XNOR U43231 ( .A(n41365), .B(n41369), .Z(n41446) );
  XNOR U43232 ( .A(n41360), .B(n41364), .Z(n41447) );
  XNOR U43233 ( .A(n41355), .B(n41359), .Z(n41448) );
  XNOR U43234 ( .A(n41350), .B(n41354), .Z(n41449) );
  XNOR U43235 ( .A(n41345), .B(n41349), .Z(n41450) );
  XNOR U43236 ( .A(n41340), .B(n41344), .Z(n41451) );
  XNOR U43237 ( .A(n41335), .B(n41339), .Z(n41452) );
  XNOR U43238 ( .A(n41330), .B(n41334), .Z(n41453) );
  XNOR U43239 ( .A(n41325), .B(n41329), .Z(n41454) );
  XNOR U43240 ( .A(n41320), .B(n41324), .Z(n41455) );
  XNOR U43241 ( .A(n41315), .B(n41319), .Z(n41456) );
  XNOR U43242 ( .A(n41310), .B(n41314), .Z(n41457) );
  XNOR U43243 ( .A(n41305), .B(n41309), .Z(n41458) );
  XNOR U43244 ( .A(n41300), .B(n41304), .Z(n41459) );
  XNOR U43245 ( .A(n41295), .B(n41299), .Z(n41460) );
  XNOR U43246 ( .A(n41290), .B(n41294), .Z(n41461) );
  XNOR U43247 ( .A(n41285), .B(n41289), .Z(n41462) );
  XNOR U43248 ( .A(n41280), .B(n41284), .Z(n41463) );
  XNOR U43249 ( .A(n41275), .B(n41279), .Z(n41464) );
  XNOR U43250 ( .A(n41270), .B(n41274), .Z(n41465) );
  XNOR U43251 ( .A(n41265), .B(n41269), .Z(n41466) );
  XNOR U43252 ( .A(n41260), .B(n41264), .Z(n41467) );
  XNOR U43253 ( .A(n41255), .B(n41259), .Z(n41468) );
  XNOR U43254 ( .A(n41250), .B(n41254), .Z(n41469) );
  XNOR U43255 ( .A(n41245), .B(n41249), .Z(n41470) );
  XNOR U43256 ( .A(n41240), .B(n41244), .Z(n41471) );
  XNOR U43257 ( .A(n41235), .B(n41239), .Z(n41472) );
  XNOR U43258 ( .A(n41230), .B(n41234), .Z(n41473) );
  XNOR U43259 ( .A(n41225), .B(n41229), .Z(n41474) );
  XNOR U43260 ( .A(n41220), .B(n41224), .Z(n41475) );
  XNOR U43261 ( .A(n41215), .B(n41219), .Z(n41476) );
  XNOR U43262 ( .A(n41210), .B(n41214), .Z(n41477) );
  XOR U43263 ( .A(n41478), .B(n41209), .Z(n41210) );
  AND U43264 ( .A(a[0]), .B(b[46]), .Z(n41478) );
  XNOR U43265 ( .A(n41479), .B(n41209), .Z(n41211) );
  XNOR U43266 ( .A(n41480), .B(n41481), .Z(n41209) );
  ANDN U43267 ( .B(n41482), .A(n41483), .Z(n41480) );
  AND U43268 ( .A(a[1]), .B(b[45]), .Z(n41479) );
  XOR U43269 ( .A(n41485), .B(n41486), .Z(n41214) );
  ANDN U43270 ( .B(n41487), .A(n41488), .Z(n41485) );
  AND U43271 ( .A(a[2]), .B(b[44]), .Z(n41484) );
  XOR U43272 ( .A(n41490), .B(n41491), .Z(n41219) );
  ANDN U43273 ( .B(n41492), .A(n41493), .Z(n41490) );
  AND U43274 ( .A(a[3]), .B(b[43]), .Z(n41489) );
  XOR U43275 ( .A(n41495), .B(n41496), .Z(n41224) );
  ANDN U43276 ( .B(n41497), .A(n41498), .Z(n41495) );
  AND U43277 ( .A(a[4]), .B(b[42]), .Z(n41494) );
  XOR U43278 ( .A(n41500), .B(n41501), .Z(n41229) );
  ANDN U43279 ( .B(n41502), .A(n41503), .Z(n41500) );
  AND U43280 ( .A(a[5]), .B(b[41]), .Z(n41499) );
  XOR U43281 ( .A(n41505), .B(n41506), .Z(n41234) );
  ANDN U43282 ( .B(n41507), .A(n41508), .Z(n41505) );
  AND U43283 ( .A(a[6]), .B(b[40]), .Z(n41504) );
  XOR U43284 ( .A(n41510), .B(n41511), .Z(n41239) );
  ANDN U43285 ( .B(n41512), .A(n41513), .Z(n41510) );
  AND U43286 ( .A(a[7]), .B(b[39]), .Z(n41509) );
  XOR U43287 ( .A(n41515), .B(n41516), .Z(n41244) );
  ANDN U43288 ( .B(n41517), .A(n41518), .Z(n41515) );
  AND U43289 ( .A(a[8]), .B(b[38]), .Z(n41514) );
  XOR U43290 ( .A(n41520), .B(n41521), .Z(n41249) );
  ANDN U43291 ( .B(n41522), .A(n41523), .Z(n41520) );
  AND U43292 ( .A(a[9]), .B(b[37]), .Z(n41519) );
  XOR U43293 ( .A(n41525), .B(n41526), .Z(n41254) );
  ANDN U43294 ( .B(n41527), .A(n41528), .Z(n41525) );
  AND U43295 ( .A(a[10]), .B(b[36]), .Z(n41524) );
  XOR U43296 ( .A(n41530), .B(n41531), .Z(n41259) );
  ANDN U43297 ( .B(n41532), .A(n41533), .Z(n41530) );
  AND U43298 ( .A(a[11]), .B(b[35]), .Z(n41529) );
  XOR U43299 ( .A(n41535), .B(n41536), .Z(n41264) );
  ANDN U43300 ( .B(n41537), .A(n41538), .Z(n41535) );
  AND U43301 ( .A(a[12]), .B(b[34]), .Z(n41534) );
  XOR U43302 ( .A(n41540), .B(n41541), .Z(n41269) );
  ANDN U43303 ( .B(n41542), .A(n41543), .Z(n41540) );
  AND U43304 ( .A(a[13]), .B(b[33]), .Z(n41539) );
  XOR U43305 ( .A(n41545), .B(n41546), .Z(n41274) );
  ANDN U43306 ( .B(n41547), .A(n41548), .Z(n41545) );
  AND U43307 ( .A(a[14]), .B(b[32]), .Z(n41544) );
  XOR U43308 ( .A(n41550), .B(n41551), .Z(n41279) );
  ANDN U43309 ( .B(n41552), .A(n41553), .Z(n41550) );
  AND U43310 ( .A(a[15]), .B(b[31]), .Z(n41549) );
  XOR U43311 ( .A(n41555), .B(n41556), .Z(n41284) );
  ANDN U43312 ( .B(n41557), .A(n41558), .Z(n41555) );
  AND U43313 ( .A(a[16]), .B(b[30]), .Z(n41554) );
  XOR U43314 ( .A(n41560), .B(n41561), .Z(n41289) );
  ANDN U43315 ( .B(n41562), .A(n41563), .Z(n41560) );
  AND U43316 ( .A(a[17]), .B(b[29]), .Z(n41559) );
  XOR U43317 ( .A(n41565), .B(n41566), .Z(n41294) );
  ANDN U43318 ( .B(n41567), .A(n41568), .Z(n41565) );
  AND U43319 ( .A(a[18]), .B(b[28]), .Z(n41564) );
  XOR U43320 ( .A(n41570), .B(n41571), .Z(n41299) );
  ANDN U43321 ( .B(n41572), .A(n41573), .Z(n41570) );
  AND U43322 ( .A(a[19]), .B(b[27]), .Z(n41569) );
  XOR U43323 ( .A(n41575), .B(n41576), .Z(n41304) );
  ANDN U43324 ( .B(n41577), .A(n41578), .Z(n41575) );
  AND U43325 ( .A(a[20]), .B(b[26]), .Z(n41574) );
  XOR U43326 ( .A(n41580), .B(n41581), .Z(n41309) );
  ANDN U43327 ( .B(n41582), .A(n41583), .Z(n41580) );
  AND U43328 ( .A(a[21]), .B(b[25]), .Z(n41579) );
  XOR U43329 ( .A(n41585), .B(n41586), .Z(n41314) );
  ANDN U43330 ( .B(n41587), .A(n41588), .Z(n41585) );
  AND U43331 ( .A(a[22]), .B(b[24]), .Z(n41584) );
  XOR U43332 ( .A(n41590), .B(n41591), .Z(n41319) );
  ANDN U43333 ( .B(n41592), .A(n41593), .Z(n41590) );
  AND U43334 ( .A(a[23]), .B(b[23]), .Z(n41589) );
  XOR U43335 ( .A(n41595), .B(n41596), .Z(n41324) );
  ANDN U43336 ( .B(n41597), .A(n41598), .Z(n41595) );
  AND U43337 ( .A(a[24]), .B(b[22]), .Z(n41594) );
  XOR U43338 ( .A(n41600), .B(n41601), .Z(n41329) );
  ANDN U43339 ( .B(n41602), .A(n41603), .Z(n41600) );
  AND U43340 ( .A(a[25]), .B(b[21]), .Z(n41599) );
  XOR U43341 ( .A(n41605), .B(n41606), .Z(n41334) );
  ANDN U43342 ( .B(n41607), .A(n41608), .Z(n41605) );
  AND U43343 ( .A(a[26]), .B(b[20]), .Z(n41604) );
  XOR U43344 ( .A(n41610), .B(n41611), .Z(n41339) );
  ANDN U43345 ( .B(n41612), .A(n41613), .Z(n41610) );
  AND U43346 ( .A(a[27]), .B(b[19]), .Z(n41609) );
  XOR U43347 ( .A(n41615), .B(n41616), .Z(n41344) );
  ANDN U43348 ( .B(n41617), .A(n41618), .Z(n41615) );
  AND U43349 ( .A(a[28]), .B(b[18]), .Z(n41614) );
  XOR U43350 ( .A(n41620), .B(n41621), .Z(n41349) );
  ANDN U43351 ( .B(n41622), .A(n41623), .Z(n41620) );
  AND U43352 ( .A(a[29]), .B(b[17]), .Z(n41619) );
  XOR U43353 ( .A(n41625), .B(n41626), .Z(n41354) );
  ANDN U43354 ( .B(n41627), .A(n41628), .Z(n41625) );
  AND U43355 ( .A(a[30]), .B(b[16]), .Z(n41624) );
  XOR U43356 ( .A(n41630), .B(n41631), .Z(n41359) );
  ANDN U43357 ( .B(n41632), .A(n41633), .Z(n41630) );
  AND U43358 ( .A(a[31]), .B(b[15]), .Z(n41629) );
  XOR U43359 ( .A(n41635), .B(n41636), .Z(n41364) );
  ANDN U43360 ( .B(n41637), .A(n41638), .Z(n41635) );
  AND U43361 ( .A(a[32]), .B(b[14]), .Z(n41634) );
  XOR U43362 ( .A(n41640), .B(n41641), .Z(n41369) );
  ANDN U43363 ( .B(n41642), .A(n41643), .Z(n41640) );
  AND U43364 ( .A(a[33]), .B(b[13]), .Z(n41639) );
  XOR U43365 ( .A(n41645), .B(n41646), .Z(n41374) );
  ANDN U43366 ( .B(n41647), .A(n41648), .Z(n41645) );
  AND U43367 ( .A(a[34]), .B(b[12]), .Z(n41644) );
  XOR U43368 ( .A(n41650), .B(n41651), .Z(n41379) );
  ANDN U43369 ( .B(n41652), .A(n41653), .Z(n41650) );
  AND U43370 ( .A(a[35]), .B(b[11]), .Z(n41649) );
  XOR U43371 ( .A(n41655), .B(n41656), .Z(n41384) );
  ANDN U43372 ( .B(n41657), .A(n41658), .Z(n41655) );
  AND U43373 ( .A(a[36]), .B(b[10]), .Z(n41654) );
  XOR U43374 ( .A(n41660), .B(n41661), .Z(n41389) );
  ANDN U43375 ( .B(n41662), .A(n41663), .Z(n41660) );
  AND U43376 ( .A(b[9]), .B(a[37]), .Z(n41659) );
  XOR U43377 ( .A(n41665), .B(n41666), .Z(n41394) );
  ANDN U43378 ( .B(n41667), .A(n41668), .Z(n41665) );
  AND U43379 ( .A(b[8]), .B(a[38]), .Z(n41664) );
  XOR U43380 ( .A(n41670), .B(n41671), .Z(n41399) );
  ANDN U43381 ( .B(n41672), .A(n41673), .Z(n41670) );
  AND U43382 ( .A(b[7]), .B(a[39]), .Z(n41669) );
  XOR U43383 ( .A(n41675), .B(n41676), .Z(n41404) );
  ANDN U43384 ( .B(n41677), .A(n41678), .Z(n41675) );
  AND U43385 ( .A(b[6]), .B(a[40]), .Z(n41674) );
  XOR U43386 ( .A(n41680), .B(n41681), .Z(n41409) );
  ANDN U43387 ( .B(n41682), .A(n41683), .Z(n41680) );
  AND U43388 ( .A(b[5]), .B(a[41]), .Z(n41679) );
  XOR U43389 ( .A(n41685), .B(n41686), .Z(n41414) );
  ANDN U43390 ( .B(n41687), .A(n41688), .Z(n41685) );
  AND U43391 ( .A(b[4]), .B(a[42]), .Z(n41684) );
  XOR U43392 ( .A(n41690), .B(n41691), .Z(n41419) );
  ANDN U43393 ( .B(n41431), .A(n41432), .Z(n41690) );
  AND U43394 ( .A(b[2]), .B(a[43]), .Z(n41692) );
  XNOR U43395 ( .A(n41687), .B(n41691), .Z(n41693) );
  XOR U43396 ( .A(n41694), .B(n41695), .Z(n41691) );
  OR U43397 ( .A(n41434), .B(n41435), .Z(n41695) );
  XNOR U43398 ( .A(n41697), .B(n41698), .Z(n41696) );
  XOR U43399 ( .A(n41697), .B(n41700), .Z(n41434) );
  NAND U43400 ( .A(b[1]), .B(a[43]), .Z(n41700) );
  IV U43401 ( .A(n41694), .Z(n41697) );
  NANDN U43402 ( .A(n125), .B(n126), .Z(n41694) );
  XOR U43403 ( .A(n41701), .B(n41702), .Z(n126) );
  NAND U43404 ( .A(a[43]), .B(b[0]), .Z(n125) );
  XNOR U43405 ( .A(n41682), .B(n41686), .Z(n41703) );
  XNOR U43406 ( .A(n41677), .B(n41681), .Z(n41704) );
  XNOR U43407 ( .A(n41672), .B(n41676), .Z(n41705) );
  XNOR U43408 ( .A(n41667), .B(n41671), .Z(n41706) );
  XNOR U43409 ( .A(n41662), .B(n41666), .Z(n41707) );
  XNOR U43410 ( .A(n41657), .B(n41661), .Z(n41708) );
  XNOR U43411 ( .A(n41652), .B(n41656), .Z(n41709) );
  XNOR U43412 ( .A(n41647), .B(n41651), .Z(n41710) );
  XNOR U43413 ( .A(n41642), .B(n41646), .Z(n41711) );
  XNOR U43414 ( .A(n41637), .B(n41641), .Z(n41712) );
  XNOR U43415 ( .A(n41632), .B(n41636), .Z(n41713) );
  XNOR U43416 ( .A(n41627), .B(n41631), .Z(n41714) );
  XNOR U43417 ( .A(n41622), .B(n41626), .Z(n41715) );
  XNOR U43418 ( .A(n41617), .B(n41621), .Z(n41716) );
  XNOR U43419 ( .A(n41612), .B(n41616), .Z(n41717) );
  XNOR U43420 ( .A(n41607), .B(n41611), .Z(n41718) );
  XNOR U43421 ( .A(n41602), .B(n41606), .Z(n41719) );
  XNOR U43422 ( .A(n41597), .B(n41601), .Z(n41720) );
  XNOR U43423 ( .A(n41592), .B(n41596), .Z(n41721) );
  XNOR U43424 ( .A(n41587), .B(n41591), .Z(n41722) );
  XNOR U43425 ( .A(n41582), .B(n41586), .Z(n41723) );
  XNOR U43426 ( .A(n41577), .B(n41581), .Z(n41724) );
  XNOR U43427 ( .A(n41572), .B(n41576), .Z(n41725) );
  XNOR U43428 ( .A(n41567), .B(n41571), .Z(n41726) );
  XNOR U43429 ( .A(n41562), .B(n41566), .Z(n41727) );
  XNOR U43430 ( .A(n41557), .B(n41561), .Z(n41728) );
  XNOR U43431 ( .A(n41552), .B(n41556), .Z(n41729) );
  XNOR U43432 ( .A(n41547), .B(n41551), .Z(n41730) );
  XNOR U43433 ( .A(n41542), .B(n41546), .Z(n41731) );
  XNOR U43434 ( .A(n41537), .B(n41541), .Z(n41732) );
  XNOR U43435 ( .A(n41532), .B(n41536), .Z(n41733) );
  XNOR U43436 ( .A(n41527), .B(n41531), .Z(n41734) );
  XNOR U43437 ( .A(n41522), .B(n41526), .Z(n41735) );
  XNOR U43438 ( .A(n41517), .B(n41521), .Z(n41736) );
  XNOR U43439 ( .A(n41512), .B(n41516), .Z(n41737) );
  XNOR U43440 ( .A(n41507), .B(n41511), .Z(n41738) );
  XNOR U43441 ( .A(n41502), .B(n41506), .Z(n41739) );
  XNOR U43442 ( .A(n41497), .B(n41501), .Z(n41740) );
  XNOR U43443 ( .A(n41492), .B(n41496), .Z(n41741) );
  XNOR U43444 ( .A(n41487), .B(n41491), .Z(n41742) );
  XNOR U43445 ( .A(n41482), .B(n41486), .Z(n41743) );
  XNOR U43446 ( .A(n41744), .B(n41481), .Z(n41482) );
  AND U43447 ( .A(a[0]), .B(b[45]), .Z(n41744) );
  XOR U43448 ( .A(n41745), .B(n41481), .Z(n41483) );
  XNOR U43449 ( .A(n41746), .B(n41747), .Z(n41481) );
  ANDN U43450 ( .B(n41748), .A(n41749), .Z(n41746) );
  AND U43451 ( .A(a[1]), .B(b[44]), .Z(n41745) );
  XOR U43452 ( .A(n41751), .B(n41752), .Z(n41486) );
  ANDN U43453 ( .B(n41753), .A(n41754), .Z(n41751) );
  AND U43454 ( .A(a[2]), .B(b[43]), .Z(n41750) );
  XOR U43455 ( .A(n41756), .B(n41757), .Z(n41491) );
  ANDN U43456 ( .B(n41758), .A(n41759), .Z(n41756) );
  AND U43457 ( .A(a[3]), .B(b[42]), .Z(n41755) );
  XOR U43458 ( .A(n41761), .B(n41762), .Z(n41496) );
  ANDN U43459 ( .B(n41763), .A(n41764), .Z(n41761) );
  AND U43460 ( .A(a[4]), .B(b[41]), .Z(n41760) );
  XOR U43461 ( .A(n41766), .B(n41767), .Z(n41501) );
  ANDN U43462 ( .B(n41768), .A(n41769), .Z(n41766) );
  AND U43463 ( .A(a[5]), .B(b[40]), .Z(n41765) );
  XOR U43464 ( .A(n41771), .B(n41772), .Z(n41506) );
  ANDN U43465 ( .B(n41773), .A(n41774), .Z(n41771) );
  AND U43466 ( .A(a[6]), .B(b[39]), .Z(n41770) );
  XOR U43467 ( .A(n41776), .B(n41777), .Z(n41511) );
  ANDN U43468 ( .B(n41778), .A(n41779), .Z(n41776) );
  AND U43469 ( .A(a[7]), .B(b[38]), .Z(n41775) );
  XOR U43470 ( .A(n41781), .B(n41782), .Z(n41516) );
  ANDN U43471 ( .B(n41783), .A(n41784), .Z(n41781) );
  AND U43472 ( .A(a[8]), .B(b[37]), .Z(n41780) );
  XOR U43473 ( .A(n41786), .B(n41787), .Z(n41521) );
  ANDN U43474 ( .B(n41788), .A(n41789), .Z(n41786) );
  AND U43475 ( .A(a[9]), .B(b[36]), .Z(n41785) );
  XOR U43476 ( .A(n41791), .B(n41792), .Z(n41526) );
  ANDN U43477 ( .B(n41793), .A(n41794), .Z(n41791) );
  AND U43478 ( .A(a[10]), .B(b[35]), .Z(n41790) );
  XOR U43479 ( .A(n41796), .B(n41797), .Z(n41531) );
  ANDN U43480 ( .B(n41798), .A(n41799), .Z(n41796) );
  AND U43481 ( .A(a[11]), .B(b[34]), .Z(n41795) );
  XOR U43482 ( .A(n41801), .B(n41802), .Z(n41536) );
  ANDN U43483 ( .B(n41803), .A(n41804), .Z(n41801) );
  AND U43484 ( .A(a[12]), .B(b[33]), .Z(n41800) );
  XOR U43485 ( .A(n41806), .B(n41807), .Z(n41541) );
  ANDN U43486 ( .B(n41808), .A(n41809), .Z(n41806) );
  AND U43487 ( .A(a[13]), .B(b[32]), .Z(n41805) );
  XOR U43488 ( .A(n41811), .B(n41812), .Z(n41546) );
  ANDN U43489 ( .B(n41813), .A(n41814), .Z(n41811) );
  AND U43490 ( .A(a[14]), .B(b[31]), .Z(n41810) );
  XOR U43491 ( .A(n41816), .B(n41817), .Z(n41551) );
  ANDN U43492 ( .B(n41818), .A(n41819), .Z(n41816) );
  AND U43493 ( .A(a[15]), .B(b[30]), .Z(n41815) );
  XOR U43494 ( .A(n41821), .B(n41822), .Z(n41556) );
  ANDN U43495 ( .B(n41823), .A(n41824), .Z(n41821) );
  AND U43496 ( .A(a[16]), .B(b[29]), .Z(n41820) );
  XOR U43497 ( .A(n41826), .B(n41827), .Z(n41561) );
  ANDN U43498 ( .B(n41828), .A(n41829), .Z(n41826) );
  AND U43499 ( .A(a[17]), .B(b[28]), .Z(n41825) );
  XOR U43500 ( .A(n41831), .B(n41832), .Z(n41566) );
  ANDN U43501 ( .B(n41833), .A(n41834), .Z(n41831) );
  AND U43502 ( .A(a[18]), .B(b[27]), .Z(n41830) );
  XOR U43503 ( .A(n41836), .B(n41837), .Z(n41571) );
  ANDN U43504 ( .B(n41838), .A(n41839), .Z(n41836) );
  AND U43505 ( .A(a[19]), .B(b[26]), .Z(n41835) );
  XOR U43506 ( .A(n41841), .B(n41842), .Z(n41576) );
  ANDN U43507 ( .B(n41843), .A(n41844), .Z(n41841) );
  AND U43508 ( .A(a[20]), .B(b[25]), .Z(n41840) );
  XOR U43509 ( .A(n41846), .B(n41847), .Z(n41581) );
  ANDN U43510 ( .B(n41848), .A(n41849), .Z(n41846) );
  AND U43511 ( .A(a[21]), .B(b[24]), .Z(n41845) );
  XOR U43512 ( .A(n41851), .B(n41852), .Z(n41586) );
  ANDN U43513 ( .B(n41853), .A(n41854), .Z(n41851) );
  AND U43514 ( .A(a[22]), .B(b[23]), .Z(n41850) );
  XOR U43515 ( .A(n41856), .B(n41857), .Z(n41591) );
  ANDN U43516 ( .B(n41858), .A(n41859), .Z(n41856) );
  AND U43517 ( .A(a[23]), .B(b[22]), .Z(n41855) );
  XOR U43518 ( .A(n41861), .B(n41862), .Z(n41596) );
  ANDN U43519 ( .B(n41863), .A(n41864), .Z(n41861) );
  AND U43520 ( .A(a[24]), .B(b[21]), .Z(n41860) );
  XOR U43521 ( .A(n41866), .B(n41867), .Z(n41601) );
  ANDN U43522 ( .B(n41868), .A(n41869), .Z(n41866) );
  AND U43523 ( .A(a[25]), .B(b[20]), .Z(n41865) );
  XOR U43524 ( .A(n41871), .B(n41872), .Z(n41606) );
  ANDN U43525 ( .B(n41873), .A(n41874), .Z(n41871) );
  AND U43526 ( .A(a[26]), .B(b[19]), .Z(n41870) );
  XOR U43527 ( .A(n41876), .B(n41877), .Z(n41611) );
  ANDN U43528 ( .B(n41878), .A(n41879), .Z(n41876) );
  AND U43529 ( .A(a[27]), .B(b[18]), .Z(n41875) );
  XOR U43530 ( .A(n41881), .B(n41882), .Z(n41616) );
  ANDN U43531 ( .B(n41883), .A(n41884), .Z(n41881) );
  AND U43532 ( .A(a[28]), .B(b[17]), .Z(n41880) );
  XOR U43533 ( .A(n41886), .B(n41887), .Z(n41621) );
  ANDN U43534 ( .B(n41888), .A(n41889), .Z(n41886) );
  AND U43535 ( .A(a[29]), .B(b[16]), .Z(n41885) );
  XOR U43536 ( .A(n41891), .B(n41892), .Z(n41626) );
  ANDN U43537 ( .B(n41893), .A(n41894), .Z(n41891) );
  AND U43538 ( .A(a[30]), .B(b[15]), .Z(n41890) );
  XOR U43539 ( .A(n41896), .B(n41897), .Z(n41631) );
  ANDN U43540 ( .B(n41898), .A(n41899), .Z(n41896) );
  AND U43541 ( .A(a[31]), .B(b[14]), .Z(n41895) );
  XOR U43542 ( .A(n41901), .B(n41902), .Z(n41636) );
  ANDN U43543 ( .B(n41903), .A(n41904), .Z(n41901) );
  AND U43544 ( .A(a[32]), .B(b[13]), .Z(n41900) );
  XOR U43545 ( .A(n41906), .B(n41907), .Z(n41641) );
  ANDN U43546 ( .B(n41908), .A(n41909), .Z(n41906) );
  AND U43547 ( .A(a[33]), .B(b[12]), .Z(n41905) );
  XOR U43548 ( .A(n41911), .B(n41912), .Z(n41646) );
  ANDN U43549 ( .B(n41913), .A(n41914), .Z(n41911) );
  AND U43550 ( .A(a[34]), .B(b[11]), .Z(n41910) );
  XOR U43551 ( .A(n41916), .B(n41917), .Z(n41651) );
  ANDN U43552 ( .B(n41918), .A(n41919), .Z(n41916) );
  AND U43553 ( .A(a[35]), .B(b[10]), .Z(n41915) );
  XOR U43554 ( .A(n41921), .B(n41922), .Z(n41656) );
  ANDN U43555 ( .B(n41923), .A(n41924), .Z(n41921) );
  AND U43556 ( .A(b[9]), .B(a[36]), .Z(n41920) );
  XOR U43557 ( .A(n41926), .B(n41927), .Z(n41661) );
  ANDN U43558 ( .B(n41928), .A(n41929), .Z(n41926) );
  AND U43559 ( .A(b[8]), .B(a[37]), .Z(n41925) );
  XOR U43560 ( .A(n41931), .B(n41932), .Z(n41666) );
  ANDN U43561 ( .B(n41933), .A(n41934), .Z(n41931) );
  AND U43562 ( .A(b[7]), .B(a[38]), .Z(n41930) );
  XOR U43563 ( .A(n41936), .B(n41937), .Z(n41671) );
  ANDN U43564 ( .B(n41938), .A(n41939), .Z(n41936) );
  AND U43565 ( .A(b[6]), .B(a[39]), .Z(n41935) );
  XOR U43566 ( .A(n41941), .B(n41942), .Z(n41676) );
  ANDN U43567 ( .B(n41943), .A(n41944), .Z(n41941) );
  AND U43568 ( .A(b[5]), .B(a[40]), .Z(n41940) );
  XOR U43569 ( .A(n41946), .B(n41947), .Z(n41681) );
  ANDN U43570 ( .B(n41948), .A(n41949), .Z(n41946) );
  AND U43571 ( .A(b[4]), .B(a[41]), .Z(n41945) );
  XOR U43572 ( .A(n41951), .B(n41952), .Z(n41686) );
  ANDN U43573 ( .B(n41698), .A(n41699), .Z(n41951) );
  AND U43574 ( .A(b[2]), .B(a[42]), .Z(n41953) );
  XNOR U43575 ( .A(n41948), .B(n41952), .Z(n41954) );
  XOR U43576 ( .A(n41955), .B(n41956), .Z(n41952) );
  OR U43577 ( .A(n41701), .B(n41702), .Z(n41956) );
  XNOR U43578 ( .A(n41958), .B(n41959), .Z(n41957) );
  XOR U43579 ( .A(n41958), .B(n41961), .Z(n41701) );
  NAND U43580 ( .A(b[1]), .B(a[42]), .Z(n41961) );
  IV U43581 ( .A(n41955), .Z(n41958) );
  NANDN U43582 ( .A(n127), .B(n128), .Z(n41955) );
  XOR U43583 ( .A(n41962), .B(n41963), .Z(n128) );
  NAND U43584 ( .A(a[42]), .B(b[0]), .Z(n127) );
  XNOR U43585 ( .A(n41943), .B(n41947), .Z(n41964) );
  XNOR U43586 ( .A(n41938), .B(n41942), .Z(n41965) );
  XNOR U43587 ( .A(n41933), .B(n41937), .Z(n41966) );
  XNOR U43588 ( .A(n41928), .B(n41932), .Z(n41967) );
  XNOR U43589 ( .A(n41923), .B(n41927), .Z(n41968) );
  XNOR U43590 ( .A(n41918), .B(n41922), .Z(n41969) );
  XNOR U43591 ( .A(n41913), .B(n41917), .Z(n41970) );
  XNOR U43592 ( .A(n41908), .B(n41912), .Z(n41971) );
  XNOR U43593 ( .A(n41903), .B(n41907), .Z(n41972) );
  XNOR U43594 ( .A(n41898), .B(n41902), .Z(n41973) );
  XNOR U43595 ( .A(n41893), .B(n41897), .Z(n41974) );
  XNOR U43596 ( .A(n41888), .B(n41892), .Z(n41975) );
  XNOR U43597 ( .A(n41883), .B(n41887), .Z(n41976) );
  XNOR U43598 ( .A(n41878), .B(n41882), .Z(n41977) );
  XNOR U43599 ( .A(n41873), .B(n41877), .Z(n41978) );
  XNOR U43600 ( .A(n41868), .B(n41872), .Z(n41979) );
  XNOR U43601 ( .A(n41863), .B(n41867), .Z(n41980) );
  XNOR U43602 ( .A(n41858), .B(n41862), .Z(n41981) );
  XNOR U43603 ( .A(n41853), .B(n41857), .Z(n41982) );
  XNOR U43604 ( .A(n41848), .B(n41852), .Z(n41983) );
  XNOR U43605 ( .A(n41843), .B(n41847), .Z(n41984) );
  XNOR U43606 ( .A(n41838), .B(n41842), .Z(n41985) );
  XNOR U43607 ( .A(n41833), .B(n41837), .Z(n41986) );
  XNOR U43608 ( .A(n41828), .B(n41832), .Z(n41987) );
  XNOR U43609 ( .A(n41823), .B(n41827), .Z(n41988) );
  XNOR U43610 ( .A(n41818), .B(n41822), .Z(n41989) );
  XNOR U43611 ( .A(n41813), .B(n41817), .Z(n41990) );
  XNOR U43612 ( .A(n41808), .B(n41812), .Z(n41991) );
  XNOR U43613 ( .A(n41803), .B(n41807), .Z(n41992) );
  XNOR U43614 ( .A(n41798), .B(n41802), .Z(n41993) );
  XNOR U43615 ( .A(n41793), .B(n41797), .Z(n41994) );
  XNOR U43616 ( .A(n41788), .B(n41792), .Z(n41995) );
  XNOR U43617 ( .A(n41783), .B(n41787), .Z(n41996) );
  XNOR U43618 ( .A(n41778), .B(n41782), .Z(n41997) );
  XNOR U43619 ( .A(n41773), .B(n41777), .Z(n41998) );
  XNOR U43620 ( .A(n41768), .B(n41772), .Z(n41999) );
  XNOR U43621 ( .A(n41763), .B(n41767), .Z(n42000) );
  XNOR U43622 ( .A(n41758), .B(n41762), .Z(n42001) );
  XNOR U43623 ( .A(n41753), .B(n41757), .Z(n42002) );
  XNOR U43624 ( .A(n41748), .B(n41752), .Z(n42003) );
  XOR U43625 ( .A(n42004), .B(n41747), .Z(n41748) );
  AND U43626 ( .A(a[0]), .B(b[44]), .Z(n42004) );
  XNOR U43627 ( .A(n42005), .B(n41747), .Z(n41749) );
  XNOR U43628 ( .A(n42006), .B(n42007), .Z(n41747) );
  ANDN U43629 ( .B(n42008), .A(n42009), .Z(n42006) );
  AND U43630 ( .A(a[1]), .B(b[43]), .Z(n42005) );
  XOR U43631 ( .A(n42011), .B(n42012), .Z(n41752) );
  ANDN U43632 ( .B(n42013), .A(n42014), .Z(n42011) );
  AND U43633 ( .A(a[2]), .B(b[42]), .Z(n42010) );
  XOR U43634 ( .A(n42016), .B(n42017), .Z(n41757) );
  ANDN U43635 ( .B(n42018), .A(n42019), .Z(n42016) );
  AND U43636 ( .A(a[3]), .B(b[41]), .Z(n42015) );
  XOR U43637 ( .A(n42021), .B(n42022), .Z(n41762) );
  ANDN U43638 ( .B(n42023), .A(n42024), .Z(n42021) );
  AND U43639 ( .A(a[4]), .B(b[40]), .Z(n42020) );
  XOR U43640 ( .A(n42026), .B(n42027), .Z(n41767) );
  ANDN U43641 ( .B(n42028), .A(n42029), .Z(n42026) );
  AND U43642 ( .A(a[5]), .B(b[39]), .Z(n42025) );
  XOR U43643 ( .A(n42031), .B(n42032), .Z(n41772) );
  ANDN U43644 ( .B(n42033), .A(n42034), .Z(n42031) );
  AND U43645 ( .A(a[6]), .B(b[38]), .Z(n42030) );
  XOR U43646 ( .A(n42036), .B(n42037), .Z(n41777) );
  ANDN U43647 ( .B(n42038), .A(n42039), .Z(n42036) );
  AND U43648 ( .A(a[7]), .B(b[37]), .Z(n42035) );
  XOR U43649 ( .A(n42041), .B(n42042), .Z(n41782) );
  ANDN U43650 ( .B(n42043), .A(n42044), .Z(n42041) );
  AND U43651 ( .A(a[8]), .B(b[36]), .Z(n42040) );
  XOR U43652 ( .A(n42046), .B(n42047), .Z(n41787) );
  ANDN U43653 ( .B(n42048), .A(n42049), .Z(n42046) );
  AND U43654 ( .A(a[9]), .B(b[35]), .Z(n42045) );
  XOR U43655 ( .A(n42051), .B(n42052), .Z(n41792) );
  ANDN U43656 ( .B(n42053), .A(n42054), .Z(n42051) );
  AND U43657 ( .A(a[10]), .B(b[34]), .Z(n42050) );
  XOR U43658 ( .A(n42056), .B(n42057), .Z(n41797) );
  ANDN U43659 ( .B(n42058), .A(n42059), .Z(n42056) );
  AND U43660 ( .A(a[11]), .B(b[33]), .Z(n42055) );
  XOR U43661 ( .A(n42061), .B(n42062), .Z(n41802) );
  ANDN U43662 ( .B(n42063), .A(n42064), .Z(n42061) );
  AND U43663 ( .A(a[12]), .B(b[32]), .Z(n42060) );
  XOR U43664 ( .A(n42066), .B(n42067), .Z(n41807) );
  ANDN U43665 ( .B(n42068), .A(n42069), .Z(n42066) );
  AND U43666 ( .A(a[13]), .B(b[31]), .Z(n42065) );
  XOR U43667 ( .A(n42071), .B(n42072), .Z(n41812) );
  ANDN U43668 ( .B(n42073), .A(n42074), .Z(n42071) );
  AND U43669 ( .A(a[14]), .B(b[30]), .Z(n42070) );
  XOR U43670 ( .A(n42076), .B(n42077), .Z(n41817) );
  ANDN U43671 ( .B(n42078), .A(n42079), .Z(n42076) );
  AND U43672 ( .A(a[15]), .B(b[29]), .Z(n42075) );
  XOR U43673 ( .A(n42081), .B(n42082), .Z(n41822) );
  ANDN U43674 ( .B(n42083), .A(n42084), .Z(n42081) );
  AND U43675 ( .A(a[16]), .B(b[28]), .Z(n42080) );
  XOR U43676 ( .A(n42086), .B(n42087), .Z(n41827) );
  ANDN U43677 ( .B(n42088), .A(n42089), .Z(n42086) );
  AND U43678 ( .A(a[17]), .B(b[27]), .Z(n42085) );
  XOR U43679 ( .A(n42091), .B(n42092), .Z(n41832) );
  ANDN U43680 ( .B(n42093), .A(n42094), .Z(n42091) );
  AND U43681 ( .A(a[18]), .B(b[26]), .Z(n42090) );
  XOR U43682 ( .A(n42096), .B(n42097), .Z(n41837) );
  ANDN U43683 ( .B(n42098), .A(n42099), .Z(n42096) );
  AND U43684 ( .A(a[19]), .B(b[25]), .Z(n42095) );
  XOR U43685 ( .A(n42101), .B(n42102), .Z(n41842) );
  ANDN U43686 ( .B(n42103), .A(n42104), .Z(n42101) );
  AND U43687 ( .A(a[20]), .B(b[24]), .Z(n42100) );
  XOR U43688 ( .A(n42106), .B(n42107), .Z(n41847) );
  ANDN U43689 ( .B(n42108), .A(n42109), .Z(n42106) );
  AND U43690 ( .A(a[21]), .B(b[23]), .Z(n42105) );
  XOR U43691 ( .A(n42111), .B(n42112), .Z(n41852) );
  ANDN U43692 ( .B(n42113), .A(n42114), .Z(n42111) );
  AND U43693 ( .A(a[22]), .B(b[22]), .Z(n42110) );
  XOR U43694 ( .A(n42116), .B(n42117), .Z(n41857) );
  ANDN U43695 ( .B(n42118), .A(n42119), .Z(n42116) );
  AND U43696 ( .A(a[23]), .B(b[21]), .Z(n42115) );
  XOR U43697 ( .A(n42121), .B(n42122), .Z(n41862) );
  ANDN U43698 ( .B(n42123), .A(n42124), .Z(n42121) );
  AND U43699 ( .A(a[24]), .B(b[20]), .Z(n42120) );
  XOR U43700 ( .A(n42126), .B(n42127), .Z(n41867) );
  ANDN U43701 ( .B(n42128), .A(n42129), .Z(n42126) );
  AND U43702 ( .A(a[25]), .B(b[19]), .Z(n42125) );
  XOR U43703 ( .A(n42131), .B(n42132), .Z(n41872) );
  ANDN U43704 ( .B(n42133), .A(n42134), .Z(n42131) );
  AND U43705 ( .A(a[26]), .B(b[18]), .Z(n42130) );
  XOR U43706 ( .A(n42136), .B(n42137), .Z(n41877) );
  ANDN U43707 ( .B(n42138), .A(n42139), .Z(n42136) );
  AND U43708 ( .A(a[27]), .B(b[17]), .Z(n42135) );
  XOR U43709 ( .A(n42141), .B(n42142), .Z(n41882) );
  ANDN U43710 ( .B(n42143), .A(n42144), .Z(n42141) );
  AND U43711 ( .A(a[28]), .B(b[16]), .Z(n42140) );
  XOR U43712 ( .A(n42146), .B(n42147), .Z(n41887) );
  ANDN U43713 ( .B(n42148), .A(n42149), .Z(n42146) );
  AND U43714 ( .A(a[29]), .B(b[15]), .Z(n42145) );
  XOR U43715 ( .A(n42151), .B(n42152), .Z(n41892) );
  ANDN U43716 ( .B(n42153), .A(n42154), .Z(n42151) );
  AND U43717 ( .A(a[30]), .B(b[14]), .Z(n42150) );
  XOR U43718 ( .A(n42156), .B(n42157), .Z(n41897) );
  ANDN U43719 ( .B(n42158), .A(n42159), .Z(n42156) );
  AND U43720 ( .A(a[31]), .B(b[13]), .Z(n42155) );
  XOR U43721 ( .A(n42161), .B(n42162), .Z(n41902) );
  ANDN U43722 ( .B(n42163), .A(n42164), .Z(n42161) );
  AND U43723 ( .A(a[32]), .B(b[12]), .Z(n42160) );
  XOR U43724 ( .A(n42166), .B(n42167), .Z(n41907) );
  ANDN U43725 ( .B(n42168), .A(n42169), .Z(n42166) );
  AND U43726 ( .A(a[33]), .B(b[11]), .Z(n42165) );
  XOR U43727 ( .A(n42171), .B(n42172), .Z(n41912) );
  ANDN U43728 ( .B(n42173), .A(n42174), .Z(n42171) );
  AND U43729 ( .A(a[34]), .B(b[10]), .Z(n42170) );
  XOR U43730 ( .A(n42176), .B(n42177), .Z(n41917) );
  ANDN U43731 ( .B(n42178), .A(n42179), .Z(n42176) );
  AND U43732 ( .A(b[9]), .B(a[35]), .Z(n42175) );
  XOR U43733 ( .A(n42181), .B(n42182), .Z(n41922) );
  ANDN U43734 ( .B(n42183), .A(n42184), .Z(n42181) );
  AND U43735 ( .A(b[8]), .B(a[36]), .Z(n42180) );
  XOR U43736 ( .A(n42186), .B(n42187), .Z(n41927) );
  ANDN U43737 ( .B(n42188), .A(n42189), .Z(n42186) );
  AND U43738 ( .A(b[7]), .B(a[37]), .Z(n42185) );
  XOR U43739 ( .A(n42191), .B(n42192), .Z(n41932) );
  ANDN U43740 ( .B(n42193), .A(n42194), .Z(n42191) );
  AND U43741 ( .A(b[6]), .B(a[38]), .Z(n42190) );
  XOR U43742 ( .A(n42196), .B(n42197), .Z(n41937) );
  ANDN U43743 ( .B(n42198), .A(n42199), .Z(n42196) );
  AND U43744 ( .A(b[5]), .B(a[39]), .Z(n42195) );
  XOR U43745 ( .A(n42201), .B(n42202), .Z(n41942) );
  ANDN U43746 ( .B(n42203), .A(n42204), .Z(n42201) );
  AND U43747 ( .A(b[4]), .B(a[40]), .Z(n42200) );
  XOR U43748 ( .A(n42206), .B(n42207), .Z(n41947) );
  ANDN U43749 ( .B(n41959), .A(n41960), .Z(n42206) );
  AND U43750 ( .A(b[2]), .B(a[41]), .Z(n42208) );
  XNOR U43751 ( .A(n42203), .B(n42207), .Z(n42209) );
  XOR U43752 ( .A(n42210), .B(n42211), .Z(n42207) );
  OR U43753 ( .A(n41962), .B(n41963), .Z(n42211) );
  XNOR U43754 ( .A(n42213), .B(n42214), .Z(n42212) );
  XOR U43755 ( .A(n42213), .B(n42216), .Z(n41962) );
  NAND U43756 ( .A(b[1]), .B(a[41]), .Z(n42216) );
  IV U43757 ( .A(n42210), .Z(n42213) );
  NANDN U43758 ( .A(n129), .B(n130), .Z(n42210) );
  XOR U43759 ( .A(n42217), .B(n42218), .Z(n130) );
  NAND U43760 ( .A(a[41]), .B(b[0]), .Z(n129) );
  XNOR U43761 ( .A(n42198), .B(n42202), .Z(n42219) );
  XNOR U43762 ( .A(n42193), .B(n42197), .Z(n42220) );
  XNOR U43763 ( .A(n42188), .B(n42192), .Z(n42221) );
  XNOR U43764 ( .A(n42183), .B(n42187), .Z(n42222) );
  XNOR U43765 ( .A(n42178), .B(n42182), .Z(n42223) );
  XNOR U43766 ( .A(n42173), .B(n42177), .Z(n42224) );
  XNOR U43767 ( .A(n42168), .B(n42172), .Z(n42225) );
  XNOR U43768 ( .A(n42163), .B(n42167), .Z(n42226) );
  XNOR U43769 ( .A(n42158), .B(n42162), .Z(n42227) );
  XNOR U43770 ( .A(n42153), .B(n42157), .Z(n42228) );
  XNOR U43771 ( .A(n42148), .B(n42152), .Z(n42229) );
  XNOR U43772 ( .A(n42143), .B(n42147), .Z(n42230) );
  XNOR U43773 ( .A(n42138), .B(n42142), .Z(n42231) );
  XNOR U43774 ( .A(n42133), .B(n42137), .Z(n42232) );
  XNOR U43775 ( .A(n42128), .B(n42132), .Z(n42233) );
  XNOR U43776 ( .A(n42123), .B(n42127), .Z(n42234) );
  XNOR U43777 ( .A(n42118), .B(n42122), .Z(n42235) );
  XNOR U43778 ( .A(n42113), .B(n42117), .Z(n42236) );
  XNOR U43779 ( .A(n42108), .B(n42112), .Z(n42237) );
  XNOR U43780 ( .A(n42103), .B(n42107), .Z(n42238) );
  XNOR U43781 ( .A(n42098), .B(n42102), .Z(n42239) );
  XNOR U43782 ( .A(n42093), .B(n42097), .Z(n42240) );
  XNOR U43783 ( .A(n42088), .B(n42092), .Z(n42241) );
  XNOR U43784 ( .A(n42083), .B(n42087), .Z(n42242) );
  XNOR U43785 ( .A(n42078), .B(n42082), .Z(n42243) );
  XNOR U43786 ( .A(n42073), .B(n42077), .Z(n42244) );
  XNOR U43787 ( .A(n42068), .B(n42072), .Z(n42245) );
  XNOR U43788 ( .A(n42063), .B(n42067), .Z(n42246) );
  XNOR U43789 ( .A(n42058), .B(n42062), .Z(n42247) );
  XNOR U43790 ( .A(n42053), .B(n42057), .Z(n42248) );
  XNOR U43791 ( .A(n42048), .B(n42052), .Z(n42249) );
  XNOR U43792 ( .A(n42043), .B(n42047), .Z(n42250) );
  XNOR U43793 ( .A(n42038), .B(n42042), .Z(n42251) );
  XNOR U43794 ( .A(n42033), .B(n42037), .Z(n42252) );
  XNOR U43795 ( .A(n42028), .B(n42032), .Z(n42253) );
  XNOR U43796 ( .A(n42023), .B(n42027), .Z(n42254) );
  XNOR U43797 ( .A(n42018), .B(n42022), .Z(n42255) );
  XNOR U43798 ( .A(n42013), .B(n42017), .Z(n42256) );
  XNOR U43799 ( .A(n42008), .B(n42012), .Z(n42257) );
  XNOR U43800 ( .A(n42258), .B(n42007), .Z(n42008) );
  AND U43801 ( .A(a[0]), .B(b[43]), .Z(n42258) );
  XOR U43802 ( .A(n42259), .B(n42007), .Z(n42009) );
  XNOR U43803 ( .A(n42260), .B(n42261), .Z(n42007) );
  ANDN U43804 ( .B(n42262), .A(n42263), .Z(n42260) );
  AND U43805 ( .A(a[1]), .B(b[42]), .Z(n42259) );
  XOR U43806 ( .A(n42265), .B(n42266), .Z(n42012) );
  ANDN U43807 ( .B(n42267), .A(n42268), .Z(n42265) );
  AND U43808 ( .A(a[2]), .B(b[41]), .Z(n42264) );
  XOR U43809 ( .A(n42270), .B(n42271), .Z(n42017) );
  ANDN U43810 ( .B(n42272), .A(n42273), .Z(n42270) );
  AND U43811 ( .A(a[3]), .B(b[40]), .Z(n42269) );
  XOR U43812 ( .A(n42275), .B(n42276), .Z(n42022) );
  ANDN U43813 ( .B(n42277), .A(n42278), .Z(n42275) );
  AND U43814 ( .A(a[4]), .B(b[39]), .Z(n42274) );
  XOR U43815 ( .A(n42280), .B(n42281), .Z(n42027) );
  ANDN U43816 ( .B(n42282), .A(n42283), .Z(n42280) );
  AND U43817 ( .A(a[5]), .B(b[38]), .Z(n42279) );
  XOR U43818 ( .A(n42285), .B(n42286), .Z(n42032) );
  ANDN U43819 ( .B(n42287), .A(n42288), .Z(n42285) );
  AND U43820 ( .A(a[6]), .B(b[37]), .Z(n42284) );
  XOR U43821 ( .A(n42290), .B(n42291), .Z(n42037) );
  ANDN U43822 ( .B(n42292), .A(n42293), .Z(n42290) );
  AND U43823 ( .A(a[7]), .B(b[36]), .Z(n42289) );
  XOR U43824 ( .A(n42295), .B(n42296), .Z(n42042) );
  ANDN U43825 ( .B(n42297), .A(n42298), .Z(n42295) );
  AND U43826 ( .A(a[8]), .B(b[35]), .Z(n42294) );
  XOR U43827 ( .A(n42300), .B(n42301), .Z(n42047) );
  ANDN U43828 ( .B(n42302), .A(n42303), .Z(n42300) );
  AND U43829 ( .A(a[9]), .B(b[34]), .Z(n42299) );
  XOR U43830 ( .A(n42305), .B(n42306), .Z(n42052) );
  ANDN U43831 ( .B(n42307), .A(n42308), .Z(n42305) );
  AND U43832 ( .A(a[10]), .B(b[33]), .Z(n42304) );
  XOR U43833 ( .A(n42310), .B(n42311), .Z(n42057) );
  ANDN U43834 ( .B(n42312), .A(n42313), .Z(n42310) );
  AND U43835 ( .A(a[11]), .B(b[32]), .Z(n42309) );
  XOR U43836 ( .A(n42315), .B(n42316), .Z(n42062) );
  ANDN U43837 ( .B(n42317), .A(n42318), .Z(n42315) );
  AND U43838 ( .A(a[12]), .B(b[31]), .Z(n42314) );
  XOR U43839 ( .A(n42320), .B(n42321), .Z(n42067) );
  ANDN U43840 ( .B(n42322), .A(n42323), .Z(n42320) );
  AND U43841 ( .A(a[13]), .B(b[30]), .Z(n42319) );
  XOR U43842 ( .A(n42325), .B(n42326), .Z(n42072) );
  ANDN U43843 ( .B(n42327), .A(n42328), .Z(n42325) );
  AND U43844 ( .A(a[14]), .B(b[29]), .Z(n42324) );
  XOR U43845 ( .A(n42330), .B(n42331), .Z(n42077) );
  ANDN U43846 ( .B(n42332), .A(n42333), .Z(n42330) );
  AND U43847 ( .A(a[15]), .B(b[28]), .Z(n42329) );
  XOR U43848 ( .A(n42335), .B(n42336), .Z(n42082) );
  ANDN U43849 ( .B(n42337), .A(n42338), .Z(n42335) );
  AND U43850 ( .A(a[16]), .B(b[27]), .Z(n42334) );
  XOR U43851 ( .A(n42340), .B(n42341), .Z(n42087) );
  ANDN U43852 ( .B(n42342), .A(n42343), .Z(n42340) );
  AND U43853 ( .A(a[17]), .B(b[26]), .Z(n42339) );
  XOR U43854 ( .A(n42345), .B(n42346), .Z(n42092) );
  ANDN U43855 ( .B(n42347), .A(n42348), .Z(n42345) );
  AND U43856 ( .A(a[18]), .B(b[25]), .Z(n42344) );
  XOR U43857 ( .A(n42350), .B(n42351), .Z(n42097) );
  ANDN U43858 ( .B(n42352), .A(n42353), .Z(n42350) );
  AND U43859 ( .A(a[19]), .B(b[24]), .Z(n42349) );
  XOR U43860 ( .A(n42355), .B(n42356), .Z(n42102) );
  ANDN U43861 ( .B(n42357), .A(n42358), .Z(n42355) );
  AND U43862 ( .A(a[20]), .B(b[23]), .Z(n42354) );
  XOR U43863 ( .A(n42360), .B(n42361), .Z(n42107) );
  ANDN U43864 ( .B(n42362), .A(n42363), .Z(n42360) );
  AND U43865 ( .A(a[21]), .B(b[22]), .Z(n42359) );
  XOR U43866 ( .A(n42365), .B(n42366), .Z(n42112) );
  ANDN U43867 ( .B(n42367), .A(n42368), .Z(n42365) );
  AND U43868 ( .A(a[22]), .B(b[21]), .Z(n42364) );
  XOR U43869 ( .A(n42370), .B(n42371), .Z(n42117) );
  ANDN U43870 ( .B(n42372), .A(n42373), .Z(n42370) );
  AND U43871 ( .A(a[23]), .B(b[20]), .Z(n42369) );
  XOR U43872 ( .A(n42375), .B(n42376), .Z(n42122) );
  ANDN U43873 ( .B(n42377), .A(n42378), .Z(n42375) );
  AND U43874 ( .A(a[24]), .B(b[19]), .Z(n42374) );
  XOR U43875 ( .A(n42380), .B(n42381), .Z(n42127) );
  ANDN U43876 ( .B(n42382), .A(n42383), .Z(n42380) );
  AND U43877 ( .A(a[25]), .B(b[18]), .Z(n42379) );
  XOR U43878 ( .A(n42385), .B(n42386), .Z(n42132) );
  ANDN U43879 ( .B(n42387), .A(n42388), .Z(n42385) );
  AND U43880 ( .A(a[26]), .B(b[17]), .Z(n42384) );
  XOR U43881 ( .A(n42390), .B(n42391), .Z(n42137) );
  ANDN U43882 ( .B(n42392), .A(n42393), .Z(n42390) );
  AND U43883 ( .A(a[27]), .B(b[16]), .Z(n42389) );
  XOR U43884 ( .A(n42395), .B(n42396), .Z(n42142) );
  ANDN U43885 ( .B(n42397), .A(n42398), .Z(n42395) );
  AND U43886 ( .A(a[28]), .B(b[15]), .Z(n42394) );
  XOR U43887 ( .A(n42400), .B(n42401), .Z(n42147) );
  ANDN U43888 ( .B(n42402), .A(n42403), .Z(n42400) );
  AND U43889 ( .A(a[29]), .B(b[14]), .Z(n42399) );
  XOR U43890 ( .A(n42405), .B(n42406), .Z(n42152) );
  ANDN U43891 ( .B(n42407), .A(n42408), .Z(n42405) );
  AND U43892 ( .A(a[30]), .B(b[13]), .Z(n42404) );
  XOR U43893 ( .A(n42410), .B(n42411), .Z(n42157) );
  ANDN U43894 ( .B(n42412), .A(n42413), .Z(n42410) );
  AND U43895 ( .A(a[31]), .B(b[12]), .Z(n42409) );
  XOR U43896 ( .A(n42415), .B(n42416), .Z(n42162) );
  ANDN U43897 ( .B(n42417), .A(n42418), .Z(n42415) );
  AND U43898 ( .A(a[32]), .B(b[11]), .Z(n42414) );
  XOR U43899 ( .A(n42420), .B(n42421), .Z(n42167) );
  ANDN U43900 ( .B(n42422), .A(n42423), .Z(n42420) );
  AND U43901 ( .A(a[33]), .B(b[10]), .Z(n42419) );
  XOR U43902 ( .A(n42425), .B(n42426), .Z(n42172) );
  ANDN U43903 ( .B(n42427), .A(n42428), .Z(n42425) );
  AND U43904 ( .A(b[9]), .B(a[34]), .Z(n42424) );
  XOR U43905 ( .A(n42430), .B(n42431), .Z(n42177) );
  ANDN U43906 ( .B(n42432), .A(n42433), .Z(n42430) );
  AND U43907 ( .A(b[8]), .B(a[35]), .Z(n42429) );
  XOR U43908 ( .A(n42435), .B(n42436), .Z(n42182) );
  ANDN U43909 ( .B(n42437), .A(n42438), .Z(n42435) );
  AND U43910 ( .A(b[7]), .B(a[36]), .Z(n42434) );
  XOR U43911 ( .A(n42440), .B(n42441), .Z(n42187) );
  ANDN U43912 ( .B(n42442), .A(n42443), .Z(n42440) );
  AND U43913 ( .A(b[6]), .B(a[37]), .Z(n42439) );
  XOR U43914 ( .A(n42445), .B(n42446), .Z(n42192) );
  ANDN U43915 ( .B(n42447), .A(n42448), .Z(n42445) );
  AND U43916 ( .A(b[5]), .B(a[38]), .Z(n42444) );
  XOR U43917 ( .A(n42450), .B(n42451), .Z(n42197) );
  ANDN U43918 ( .B(n42452), .A(n42453), .Z(n42450) );
  AND U43919 ( .A(b[4]), .B(a[39]), .Z(n42449) );
  XOR U43920 ( .A(n42455), .B(n42456), .Z(n42202) );
  ANDN U43921 ( .B(n42214), .A(n42215), .Z(n42455) );
  AND U43922 ( .A(b[2]), .B(a[40]), .Z(n42457) );
  XNOR U43923 ( .A(n42452), .B(n42456), .Z(n42458) );
  XOR U43924 ( .A(n42459), .B(n42460), .Z(n42456) );
  OR U43925 ( .A(n42217), .B(n42218), .Z(n42460) );
  XNOR U43926 ( .A(n42462), .B(n42463), .Z(n42461) );
  XOR U43927 ( .A(n42462), .B(n42465), .Z(n42217) );
  NAND U43928 ( .A(b[1]), .B(a[40]), .Z(n42465) );
  IV U43929 ( .A(n42459), .Z(n42462) );
  NANDN U43930 ( .A(n131), .B(n132), .Z(n42459) );
  XOR U43931 ( .A(n42466), .B(n42467), .Z(n132) );
  NAND U43932 ( .A(a[40]), .B(b[0]), .Z(n131) );
  XNOR U43933 ( .A(n42447), .B(n42451), .Z(n42468) );
  XNOR U43934 ( .A(n42442), .B(n42446), .Z(n42469) );
  XNOR U43935 ( .A(n42437), .B(n42441), .Z(n42470) );
  XNOR U43936 ( .A(n42432), .B(n42436), .Z(n42471) );
  XNOR U43937 ( .A(n42427), .B(n42431), .Z(n42472) );
  XNOR U43938 ( .A(n42422), .B(n42426), .Z(n42473) );
  XNOR U43939 ( .A(n42417), .B(n42421), .Z(n42474) );
  XNOR U43940 ( .A(n42412), .B(n42416), .Z(n42475) );
  XNOR U43941 ( .A(n42407), .B(n42411), .Z(n42476) );
  XNOR U43942 ( .A(n42402), .B(n42406), .Z(n42477) );
  XNOR U43943 ( .A(n42397), .B(n42401), .Z(n42478) );
  XNOR U43944 ( .A(n42392), .B(n42396), .Z(n42479) );
  XNOR U43945 ( .A(n42387), .B(n42391), .Z(n42480) );
  XNOR U43946 ( .A(n42382), .B(n42386), .Z(n42481) );
  XNOR U43947 ( .A(n42377), .B(n42381), .Z(n42482) );
  XNOR U43948 ( .A(n42372), .B(n42376), .Z(n42483) );
  XNOR U43949 ( .A(n42367), .B(n42371), .Z(n42484) );
  XNOR U43950 ( .A(n42362), .B(n42366), .Z(n42485) );
  XNOR U43951 ( .A(n42357), .B(n42361), .Z(n42486) );
  XNOR U43952 ( .A(n42352), .B(n42356), .Z(n42487) );
  XNOR U43953 ( .A(n42347), .B(n42351), .Z(n42488) );
  XNOR U43954 ( .A(n42342), .B(n42346), .Z(n42489) );
  XNOR U43955 ( .A(n42337), .B(n42341), .Z(n42490) );
  XNOR U43956 ( .A(n42332), .B(n42336), .Z(n42491) );
  XNOR U43957 ( .A(n42327), .B(n42331), .Z(n42492) );
  XNOR U43958 ( .A(n42322), .B(n42326), .Z(n42493) );
  XNOR U43959 ( .A(n42317), .B(n42321), .Z(n42494) );
  XNOR U43960 ( .A(n42312), .B(n42316), .Z(n42495) );
  XNOR U43961 ( .A(n42307), .B(n42311), .Z(n42496) );
  XNOR U43962 ( .A(n42302), .B(n42306), .Z(n42497) );
  XNOR U43963 ( .A(n42297), .B(n42301), .Z(n42498) );
  XNOR U43964 ( .A(n42292), .B(n42296), .Z(n42499) );
  XNOR U43965 ( .A(n42287), .B(n42291), .Z(n42500) );
  XNOR U43966 ( .A(n42282), .B(n42286), .Z(n42501) );
  XNOR U43967 ( .A(n42277), .B(n42281), .Z(n42502) );
  XNOR U43968 ( .A(n42272), .B(n42276), .Z(n42503) );
  XNOR U43969 ( .A(n42267), .B(n42271), .Z(n42504) );
  XNOR U43970 ( .A(n42262), .B(n42266), .Z(n42505) );
  XOR U43971 ( .A(n42506), .B(n42261), .Z(n42262) );
  AND U43972 ( .A(a[0]), .B(b[42]), .Z(n42506) );
  XNOR U43973 ( .A(n42507), .B(n42261), .Z(n42263) );
  XNOR U43974 ( .A(n42508), .B(n42509), .Z(n42261) );
  ANDN U43975 ( .B(n42510), .A(n42511), .Z(n42508) );
  AND U43976 ( .A(a[1]), .B(b[41]), .Z(n42507) );
  XOR U43977 ( .A(n42513), .B(n42514), .Z(n42266) );
  ANDN U43978 ( .B(n42515), .A(n42516), .Z(n42513) );
  AND U43979 ( .A(a[2]), .B(b[40]), .Z(n42512) );
  XOR U43980 ( .A(n42518), .B(n42519), .Z(n42271) );
  ANDN U43981 ( .B(n42520), .A(n42521), .Z(n42518) );
  AND U43982 ( .A(a[3]), .B(b[39]), .Z(n42517) );
  XOR U43983 ( .A(n42523), .B(n42524), .Z(n42276) );
  ANDN U43984 ( .B(n42525), .A(n42526), .Z(n42523) );
  AND U43985 ( .A(a[4]), .B(b[38]), .Z(n42522) );
  XOR U43986 ( .A(n42528), .B(n42529), .Z(n42281) );
  ANDN U43987 ( .B(n42530), .A(n42531), .Z(n42528) );
  AND U43988 ( .A(a[5]), .B(b[37]), .Z(n42527) );
  XOR U43989 ( .A(n42533), .B(n42534), .Z(n42286) );
  ANDN U43990 ( .B(n42535), .A(n42536), .Z(n42533) );
  AND U43991 ( .A(a[6]), .B(b[36]), .Z(n42532) );
  XOR U43992 ( .A(n42538), .B(n42539), .Z(n42291) );
  ANDN U43993 ( .B(n42540), .A(n42541), .Z(n42538) );
  AND U43994 ( .A(a[7]), .B(b[35]), .Z(n42537) );
  XOR U43995 ( .A(n42543), .B(n42544), .Z(n42296) );
  ANDN U43996 ( .B(n42545), .A(n42546), .Z(n42543) );
  AND U43997 ( .A(a[8]), .B(b[34]), .Z(n42542) );
  XOR U43998 ( .A(n42548), .B(n42549), .Z(n42301) );
  ANDN U43999 ( .B(n42550), .A(n42551), .Z(n42548) );
  AND U44000 ( .A(a[9]), .B(b[33]), .Z(n42547) );
  XOR U44001 ( .A(n42553), .B(n42554), .Z(n42306) );
  ANDN U44002 ( .B(n42555), .A(n42556), .Z(n42553) );
  AND U44003 ( .A(a[10]), .B(b[32]), .Z(n42552) );
  XOR U44004 ( .A(n42558), .B(n42559), .Z(n42311) );
  ANDN U44005 ( .B(n42560), .A(n42561), .Z(n42558) );
  AND U44006 ( .A(a[11]), .B(b[31]), .Z(n42557) );
  XOR U44007 ( .A(n42563), .B(n42564), .Z(n42316) );
  ANDN U44008 ( .B(n42565), .A(n42566), .Z(n42563) );
  AND U44009 ( .A(a[12]), .B(b[30]), .Z(n42562) );
  XOR U44010 ( .A(n42568), .B(n42569), .Z(n42321) );
  ANDN U44011 ( .B(n42570), .A(n42571), .Z(n42568) );
  AND U44012 ( .A(a[13]), .B(b[29]), .Z(n42567) );
  XOR U44013 ( .A(n42573), .B(n42574), .Z(n42326) );
  ANDN U44014 ( .B(n42575), .A(n42576), .Z(n42573) );
  AND U44015 ( .A(a[14]), .B(b[28]), .Z(n42572) );
  XOR U44016 ( .A(n42578), .B(n42579), .Z(n42331) );
  ANDN U44017 ( .B(n42580), .A(n42581), .Z(n42578) );
  AND U44018 ( .A(a[15]), .B(b[27]), .Z(n42577) );
  XOR U44019 ( .A(n42583), .B(n42584), .Z(n42336) );
  ANDN U44020 ( .B(n42585), .A(n42586), .Z(n42583) );
  AND U44021 ( .A(a[16]), .B(b[26]), .Z(n42582) );
  XOR U44022 ( .A(n42588), .B(n42589), .Z(n42341) );
  ANDN U44023 ( .B(n42590), .A(n42591), .Z(n42588) );
  AND U44024 ( .A(a[17]), .B(b[25]), .Z(n42587) );
  XOR U44025 ( .A(n42593), .B(n42594), .Z(n42346) );
  ANDN U44026 ( .B(n42595), .A(n42596), .Z(n42593) );
  AND U44027 ( .A(a[18]), .B(b[24]), .Z(n42592) );
  XOR U44028 ( .A(n42598), .B(n42599), .Z(n42351) );
  ANDN U44029 ( .B(n42600), .A(n42601), .Z(n42598) );
  AND U44030 ( .A(a[19]), .B(b[23]), .Z(n42597) );
  XOR U44031 ( .A(n42603), .B(n42604), .Z(n42356) );
  ANDN U44032 ( .B(n42605), .A(n42606), .Z(n42603) );
  AND U44033 ( .A(a[20]), .B(b[22]), .Z(n42602) );
  XOR U44034 ( .A(n42608), .B(n42609), .Z(n42361) );
  ANDN U44035 ( .B(n42610), .A(n42611), .Z(n42608) );
  AND U44036 ( .A(a[21]), .B(b[21]), .Z(n42607) );
  XOR U44037 ( .A(n42613), .B(n42614), .Z(n42366) );
  ANDN U44038 ( .B(n42615), .A(n42616), .Z(n42613) );
  AND U44039 ( .A(a[22]), .B(b[20]), .Z(n42612) );
  XOR U44040 ( .A(n42618), .B(n42619), .Z(n42371) );
  ANDN U44041 ( .B(n42620), .A(n42621), .Z(n42618) );
  AND U44042 ( .A(a[23]), .B(b[19]), .Z(n42617) );
  XOR U44043 ( .A(n42623), .B(n42624), .Z(n42376) );
  ANDN U44044 ( .B(n42625), .A(n42626), .Z(n42623) );
  AND U44045 ( .A(a[24]), .B(b[18]), .Z(n42622) );
  XOR U44046 ( .A(n42628), .B(n42629), .Z(n42381) );
  ANDN U44047 ( .B(n42630), .A(n42631), .Z(n42628) );
  AND U44048 ( .A(a[25]), .B(b[17]), .Z(n42627) );
  XOR U44049 ( .A(n42633), .B(n42634), .Z(n42386) );
  ANDN U44050 ( .B(n42635), .A(n42636), .Z(n42633) );
  AND U44051 ( .A(a[26]), .B(b[16]), .Z(n42632) );
  XOR U44052 ( .A(n42638), .B(n42639), .Z(n42391) );
  ANDN U44053 ( .B(n42640), .A(n42641), .Z(n42638) );
  AND U44054 ( .A(a[27]), .B(b[15]), .Z(n42637) );
  XOR U44055 ( .A(n42643), .B(n42644), .Z(n42396) );
  ANDN U44056 ( .B(n42645), .A(n42646), .Z(n42643) );
  AND U44057 ( .A(a[28]), .B(b[14]), .Z(n42642) );
  XOR U44058 ( .A(n42648), .B(n42649), .Z(n42401) );
  ANDN U44059 ( .B(n42650), .A(n42651), .Z(n42648) );
  AND U44060 ( .A(a[29]), .B(b[13]), .Z(n42647) );
  XOR U44061 ( .A(n42653), .B(n42654), .Z(n42406) );
  ANDN U44062 ( .B(n42655), .A(n42656), .Z(n42653) );
  AND U44063 ( .A(a[30]), .B(b[12]), .Z(n42652) );
  XOR U44064 ( .A(n42658), .B(n42659), .Z(n42411) );
  ANDN U44065 ( .B(n42660), .A(n42661), .Z(n42658) );
  AND U44066 ( .A(a[31]), .B(b[11]), .Z(n42657) );
  XOR U44067 ( .A(n42663), .B(n42664), .Z(n42416) );
  ANDN U44068 ( .B(n42665), .A(n42666), .Z(n42663) );
  AND U44069 ( .A(a[32]), .B(b[10]), .Z(n42662) );
  XOR U44070 ( .A(n42668), .B(n42669), .Z(n42421) );
  ANDN U44071 ( .B(n42670), .A(n42671), .Z(n42668) );
  AND U44072 ( .A(b[9]), .B(a[33]), .Z(n42667) );
  XOR U44073 ( .A(n42673), .B(n42674), .Z(n42426) );
  ANDN U44074 ( .B(n42675), .A(n42676), .Z(n42673) );
  AND U44075 ( .A(b[8]), .B(a[34]), .Z(n42672) );
  XOR U44076 ( .A(n42678), .B(n42679), .Z(n42431) );
  ANDN U44077 ( .B(n42680), .A(n42681), .Z(n42678) );
  AND U44078 ( .A(b[7]), .B(a[35]), .Z(n42677) );
  XOR U44079 ( .A(n42683), .B(n42684), .Z(n42436) );
  ANDN U44080 ( .B(n42685), .A(n42686), .Z(n42683) );
  AND U44081 ( .A(b[6]), .B(a[36]), .Z(n42682) );
  XOR U44082 ( .A(n42688), .B(n42689), .Z(n42441) );
  ANDN U44083 ( .B(n42690), .A(n42691), .Z(n42688) );
  AND U44084 ( .A(b[5]), .B(a[37]), .Z(n42687) );
  XOR U44085 ( .A(n42693), .B(n42694), .Z(n42446) );
  ANDN U44086 ( .B(n42695), .A(n42696), .Z(n42693) );
  AND U44087 ( .A(b[4]), .B(a[38]), .Z(n42692) );
  XOR U44088 ( .A(n42698), .B(n42699), .Z(n42451) );
  ANDN U44089 ( .B(n42463), .A(n42464), .Z(n42698) );
  AND U44090 ( .A(b[2]), .B(a[39]), .Z(n42700) );
  XNOR U44091 ( .A(n42695), .B(n42699), .Z(n42701) );
  XOR U44092 ( .A(n42702), .B(n42703), .Z(n42699) );
  OR U44093 ( .A(n42466), .B(n42467), .Z(n42703) );
  XNOR U44094 ( .A(n42705), .B(n42706), .Z(n42704) );
  XOR U44095 ( .A(n42705), .B(n42708), .Z(n42466) );
  NAND U44096 ( .A(b[1]), .B(a[39]), .Z(n42708) );
  IV U44097 ( .A(n42702), .Z(n42705) );
  NANDN U44098 ( .A(n135), .B(n136), .Z(n42702) );
  XOR U44099 ( .A(n42709), .B(n42710), .Z(n136) );
  NAND U44100 ( .A(a[39]), .B(b[0]), .Z(n135) );
  XNOR U44101 ( .A(n42690), .B(n42694), .Z(n42711) );
  XNOR U44102 ( .A(n42685), .B(n42689), .Z(n42712) );
  XNOR U44103 ( .A(n42680), .B(n42684), .Z(n42713) );
  XNOR U44104 ( .A(n42675), .B(n42679), .Z(n42714) );
  XNOR U44105 ( .A(n42670), .B(n42674), .Z(n42715) );
  XNOR U44106 ( .A(n42665), .B(n42669), .Z(n42716) );
  XNOR U44107 ( .A(n42660), .B(n42664), .Z(n42717) );
  XNOR U44108 ( .A(n42655), .B(n42659), .Z(n42718) );
  XNOR U44109 ( .A(n42650), .B(n42654), .Z(n42719) );
  XNOR U44110 ( .A(n42645), .B(n42649), .Z(n42720) );
  XNOR U44111 ( .A(n42640), .B(n42644), .Z(n42721) );
  XNOR U44112 ( .A(n42635), .B(n42639), .Z(n42722) );
  XNOR U44113 ( .A(n42630), .B(n42634), .Z(n42723) );
  XNOR U44114 ( .A(n42625), .B(n42629), .Z(n42724) );
  XNOR U44115 ( .A(n42620), .B(n42624), .Z(n42725) );
  XNOR U44116 ( .A(n42615), .B(n42619), .Z(n42726) );
  XNOR U44117 ( .A(n42610), .B(n42614), .Z(n42727) );
  XNOR U44118 ( .A(n42605), .B(n42609), .Z(n42728) );
  XNOR U44119 ( .A(n42600), .B(n42604), .Z(n42729) );
  XNOR U44120 ( .A(n42595), .B(n42599), .Z(n42730) );
  XNOR U44121 ( .A(n42590), .B(n42594), .Z(n42731) );
  XNOR U44122 ( .A(n42585), .B(n42589), .Z(n42732) );
  XNOR U44123 ( .A(n42580), .B(n42584), .Z(n42733) );
  XNOR U44124 ( .A(n42575), .B(n42579), .Z(n42734) );
  XNOR U44125 ( .A(n42570), .B(n42574), .Z(n42735) );
  XNOR U44126 ( .A(n42565), .B(n42569), .Z(n42736) );
  XNOR U44127 ( .A(n42560), .B(n42564), .Z(n42737) );
  XNOR U44128 ( .A(n42555), .B(n42559), .Z(n42738) );
  XNOR U44129 ( .A(n42550), .B(n42554), .Z(n42739) );
  XNOR U44130 ( .A(n42545), .B(n42549), .Z(n42740) );
  XNOR U44131 ( .A(n42540), .B(n42544), .Z(n42741) );
  XNOR U44132 ( .A(n42535), .B(n42539), .Z(n42742) );
  XNOR U44133 ( .A(n42530), .B(n42534), .Z(n42743) );
  XNOR U44134 ( .A(n42525), .B(n42529), .Z(n42744) );
  XNOR U44135 ( .A(n42520), .B(n42524), .Z(n42745) );
  XNOR U44136 ( .A(n42515), .B(n42519), .Z(n42746) );
  XNOR U44137 ( .A(n42510), .B(n42514), .Z(n42747) );
  XNOR U44138 ( .A(n42748), .B(n42509), .Z(n42510) );
  AND U44139 ( .A(a[0]), .B(b[41]), .Z(n42748) );
  XOR U44140 ( .A(n42749), .B(n42509), .Z(n42511) );
  XNOR U44141 ( .A(n42750), .B(n42751), .Z(n42509) );
  ANDN U44142 ( .B(n42752), .A(n42753), .Z(n42750) );
  AND U44143 ( .A(a[1]), .B(b[40]), .Z(n42749) );
  XOR U44144 ( .A(n42755), .B(n42756), .Z(n42514) );
  ANDN U44145 ( .B(n42757), .A(n42758), .Z(n42755) );
  AND U44146 ( .A(a[2]), .B(b[39]), .Z(n42754) );
  XOR U44147 ( .A(n42760), .B(n42761), .Z(n42519) );
  ANDN U44148 ( .B(n42762), .A(n42763), .Z(n42760) );
  AND U44149 ( .A(a[3]), .B(b[38]), .Z(n42759) );
  XOR U44150 ( .A(n42765), .B(n42766), .Z(n42524) );
  ANDN U44151 ( .B(n42767), .A(n42768), .Z(n42765) );
  AND U44152 ( .A(a[4]), .B(b[37]), .Z(n42764) );
  XOR U44153 ( .A(n42770), .B(n42771), .Z(n42529) );
  ANDN U44154 ( .B(n42772), .A(n42773), .Z(n42770) );
  AND U44155 ( .A(a[5]), .B(b[36]), .Z(n42769) );
  XOR U44156 ( .A(n42775), .B(n42776), .Z(n42534) );
  ANDN U44157 ( .B(n42777), .A(n42778), .Z(n42775) );
  AND U44158 ( .A(a[6]), .B(b[35]), .Z(n42774) );
  XOR U44159 ( .A(n42780), .B(n42781), .Z(n42539) );
  ANDN U44160 ( .B(n42782), .A(n42783), .Z(n42780) );
  AND U44161 ( .A(a[7]), .B(b[34]), .Z(n42779) );
  XOR U44162 ( .A(n42785), .B(n42786), .Z(n42544) );
  ANDN U44163 ( .B(n42787), .A(n42788), .Z(n42785) );
  AND U44164 ( .A(a[8]), .B(b[33]), .Z(n42784) );
  XOR U44165 ( .A(n42790), .B(n42791), .Z(n42549) );
  ANDN U44166 ( .B(n42792), .A(n42793), .Z(n42790) );
  AND U44167 ( .A(a[9]), .B(b[32]), .Z(n42789) );
  XOR U44168 ( .A(n42795), .B(n42796), .Z(n42554) );
  ANDN U44169 ( .B(n42797), .A(n42798), .Z(n42795) );
  AND U44170 ( .A(a[10]), .B(b[31]), .Z(n42794) );
  XOR U44171 ( .A(n42800), .B(n42801), .Z(n42559) );
  ANDN U44172 ( .B(n42802), .A(n42803), .Z(n42800) );
  AND U44173 ( .A(a[11]), .B(b[30]), .Z(n42799) );
  XOR U44174 ( .A(n42805), .B(n42806), .Z(n42564) );
  ANDN U44175 ( .B(n42807), .A(n42808), .Z(n42805) );
  AND U44176 ( .A(a[12]), .B(b[29]), .Z(n42804) );
  XOR U44177 ( .A(n42810), .B(n42811), .Z(n42569) );
  ANDN U44178 ( .B(n42812), .A(n42813), .Z(n42810) );
  AND U44179 ( .A(a[13]), .B(b[28]), .Z(n42809) );
  XOR U44180 ( .A(n42815), .B(n42816), .Z(n42574) );
  ANDN U44181 ( .B(n42817), .A(n42818), .Z(n42815) );
  AND U44182 ( .A(a[14]), .B(b[27]), .Z(n42814) );
  XOR U44183 ( .A(n42820), .B(n42821), .Z(n42579) );
  ANDN U44184 ( .B(n42822), .A(n42823), .Z(n42820) );
  AND U44185 ( .A(a[15]), .B(b[26]), .Z(n42819) );
  XOR U44186 ( .A(n42825), .B(n42826), .Z(n42584) );
  ANDN U44187 ( .B(n42827), .A(n42828), .Z(n42825) );
  AND U44188 ( .A(a[16]), .B(b[25]), .Z(n42824) );
  XOR U44189 ( .A(n42830), .B(n42831), .Z(n42589) );
  ANDN U44190 ( .B(n42832), .A(n42833), .Z(n42830) );
  AND U44191 ( .A(a[17]), .B(b[24]), .Z(n42829) );
  XOR U44192 ( .A(n42835), .B(n42836), .Z(n42594) );
  ANDN U44193 ( .B(n42837), .A(n42838), .Z(n42835) );
  AND U44194 ( .A(a[18]), .B(b[23]), .Z(n42834) );
  XOR U44195 ( .A(n42840), .B(n42841), .Z(n42599) );
  ANDN U44196 ( .B(n42842), .A(n42843), .Z(n42840) );
  AND U44197 ( .A(a[19]), .B(b[22]), .Z(n42839) );
  XOR U44198 ( .A(n42845), .B(n42846), .Z(n42604) );
  ANDN U44199 ( .B(n42847), .A(n42848), .Z(n42845) );
  AND U44200 ( .A(a[20]), .B(b[21]), .Z(n42844) );
  XOR U44201 ( .A(n42850), .B(n42851), .Z(n42609) );
  ANDN U44202 ( .B(n42852), .A(n42853), .Z(n42850) );
  AND U44203 ( .A(a[21]), .B(b[20]), .Z(n42849) );
  XOR U44204 ( .A(n42855), .B(n42856), .Z(n42614) );
  ANDN U44205 ( .B(n42857), .A(n42858), .Z(n42855) );
  AND U44206 ( .A(a[22]), .B(b[19]), .Z(n42854) );
  XOR U44207 ( .A(n42860), .B(n42861), .Z(n42619) );
  ANDN U44208 ( .B(n42862), .A(n42863), .Z(n42860) );
  AND U44209 ( .A(a[23]), .B(b[18]), .Z(n42859) );
  XOR U44210 ( .A(n42865), .B(n42866), .Z(n42624) );
  ANDN U44211 ( .B(n42867), .A(n42868), .Z(n42865) );
  AND U44212 ( .A(a[24]), .B(b[17]), .Z(n42864) );
  XOR U44213 ( .A(n42870), .B(n42871), .Z(n42629) );
  ANDN U44214 ( .B(n42872), .A(n42873), .Z(n42870) );
  AND U44215 ( .A(a[25]), .B(b[16]), .Z(n42869) );
  XOR U44216 ( .A(n42875), .B(n42876), .Z(n42634) );
  ANDN U44217 ( .B(n42877), .A(n42878), .Z(n42875) );
  AND U44218 ( .A(a[26]), .B(b[15]), .Z(n42874) );
  XOR U44219 ( .A(n42880), .B(n42881), .Z(n42639) );
  ANDN U44220 ( .B(n42882), .A(n42883), .Z(n42880) );
  AND U44221 ( .A(a[27]), .B(b[14]), .Z(n42879) );
  XOR U44222 ( .A(n42885), .B(n42886), .Z(n42644) );
  ANDN U44223 ( .B(n42887), .A(n42888), .Z(n42885) );
  AND U44224 ( .A(a[28]), .B(b[13]), .Z(n42884) );
  XOR U44225 ( .A(n42890), .B(n42891), .Z(n42649) );
  ANDN U44226 ( .B(n42892), .A(n42893), .Z(n42890) );
  AND U44227 ( .A(a[29]), .B(b[12]), .Z(n42889) );
  XOR U44228 ( .A(n42895), .B(n42896), .Z(n42654) );
  ANDN U44229 ( .B(n42897), .A(n42898), .Z(n42895) );
  AND U44230 ( .A(a[30]), .B(b[11]), .Z(n42894) );
  XOR U44231 ( .A(n42900), .B(n42901), .Z(n42659) );
  ANDN U44232 ( .B(n42902), .A(n42903), .Z(n42900) );
  AND U44233 ( .A(a[31]), .B(b[10]), .Z(n42899) );
  XOR U44234 ( .A(n42905), .B(n42906), .Z(n42664) );
  ANDN U44235 ( .B(n42907), .A(n42908), .Z(n42905) );
  AND U44236 ( .A(b[9]), .B(a[32]), .Z(n42904) );
  XOR U44237 ( .A(n42910), .B(n42911), .Z(n42669) );
  ANDN U44238 ( .B(n42912), .A(n42913), .Z(n42910) );
  AND U44239 ( .A(b[8]), .B(a[33]), .Z(n42909) );
  XOR U44240 ( .A(n42915), .B(n42916), .Z(n42674) );
  ANDN U44241 ( .B(n42917), .A(n42918), .Z(n42915) );
  AND U44242 ( .A(b[7]), .B(a[34]), .Z(n42914) );
  XOR U44243 ( .A(n42920), .B(n42921), .Z(n42679) );
  ANDN U44244 ( .B(n42922), .A(n42923), .Z(n42920) );
  AND U44245 ( .A(b[6]), .B(a[35]), .Z(n42919) );
  XOR U44246 ( .A(n42925), .B(n42926), .Z(n42684) );
  ANDN U44247 ( .B(n42927), .A(n42928), .Z(n42925) );
  AND U44248 ( .A(b[5]), .B(a[36]), .Z(n42924) );
  XOR U44249 ( .A(n42930), .B(n42931), .Z(n42689) );
  ANDN U44250 ( .B(n42932), .A(n42933), .Z(n42930) );
  AND U44251 ( .A(b[4]), .B(a[37]), .Z(n42929) );
  XOR U44252 ( .A(n42935), .B(n42936), .Z(n42694) );
  ANDN U44253 ( .B(n42706), .A(n42707), .Z(n42935) );
  AND U44254 ( .A(b[2]), .B(a[38]), .Z(n42937) );
  XNOR U44255 ( .A(n42932), .B(n42936), .Z(n42938) );
  XOR U44256 ( .A(n42939), .B(n42940), .Z(n42936) );
  OR U44257 ( .A(n42709), .B(n42710), .Z(n42940) );
  XNOR U44258 ( .A(n42942), .B(n42943), .Z(n42941) );
  XOR U44259 ( .A(n42942), .B(n42945), .Z(n42709) );
  NAND U44260 ( .A(b[1]), .B(a[38]), .Z(n42945) );
  IV U44261 ( .A(n42939), .Z(n42942) );
  NANDN U44262 ( .A(n137), .B(n138), .Z(n42939) );
  XOR U44263 ( .A(n42946), .B(n42947), .Z(n138) );
  NAND U44264 ( .A(a[38]), .B(b[0]), .Z(n137) );
  XNOR U44265 ( .A(n42927), .B(n42931), .Z(n42948) );
  XNOR U44266 ( .A(n42922), .B(n42926), .Z(n42949) );
  XNOR U44267 ( .A(n42917), .B(n42921), .Z(n42950) );
  XNOR U44268 ( .A(n42912), .B(n42916), .Z(n42951) );
  XNOR U44269 ( .A(n42907), .B(n42911), .Z(n42952) );
  XNOR U44270 ( .A(n42902), .B(n42906), .Z(n42953) );
  XNOR U44271 ( .A(n42897), .B(n42901), .Z(n42954) );
  XNOR U44272 ( .A(n42892), .B(n42896), .Z(n42955) );
  XNOR U44273 ( .A(n42887), .B(n42891), .Z(n42956) );
  XNOR U44274 ( .A(n42882), .B(n42886), .Z(n42957) );
  XNOR U44275 ( .A(n42877), .B(n42881), .Z(n42958) );
  XNOR U44276 ( .A(n42872), .B(n42876), .Z(n42959) );
  XNOR U44277 ( .A(n42867), .B(n42871), .Z(n42960) );
  XNOR U44278 ( .A(n42862), .B(n42866), .Z(n42961) );
  XNOR U44279 ( .A(n42857), .B(n42861), .Z(n42962) );
  XNOR U44280 ( .A(n42852), .B(n42856), .Z(n42963) );
  XNOR U44281 ( .A(n42847), .B(n42851), .Z(n42964) );
  XNOR U44282 ( .A(n42842), .B(n42846), .Z(n42965) );
  XNOR U44283 ( .A(n42837), .B(n42841), .Z(n42966) );
  XNOR U44284 ( .A(n42832), .B(n42836), .Z(n42967) );
  XNOR U44285 ( .A(n42827), .B(n42831), .Z(n42968) );
  XNOR U44286 ( .A(n42822), .B(n42826), .Z(n42969) );
  XNOR U44287 ( .A(n42817), .B(n42821), .Z(n42970) );
  XNOR U44288 ( .A(n42812), .B(n42816), .Z(n42971) );
  XNOR U44289 ( .A(n42807), .B(n42811), .Z(n42972) );
  XNOR U44290 ( .A(n42802), .B(n42806), .Z(n42973) );
  XNOR U44291 ( .A(n42797), .B(n42801), .Z(n42974) );
  XNOR U44292 ( .A(n42792), .B(n42796), .Z(n42975) );
  XNOR U44293 ( .A(n42787), .B(n42791), .Z(n42976) );
  XNOR U44294 ( .A(n42782), .B(n42786), .Z(n42977) );
  XNOR U44295 ( .A(n42777), .B(n42781), .Z(n42978) );
  XNOR U44296 ( .A(n42772), .B(n42776), .Z(n42979) );
  XNOR U44297 ( .A(n42767), .B(n42771), .Z(n42980) );
  XNOR U44298 ( .A(n42762), .B(n42766), .Z(n42981) );
  XNOR U44299 ( .A(n42757), .B(n42761), .Z(n42982) );
  XNOR U44300 ( .A(n42752), .B(n42756), .Z(n42983) );
  XOR U44301 ( .A(n42984), .B(n42751), .Z(n42752) );
  AND U44302 ( .A(a[0]), .B(b[40]), .Z(n42984) );
  XNOR U44303 ( .A(n42985), .B(n42751), .Z(n42753) );
  XNOR U44304 ( .A(n42986), .B(n42987), .Z(n42751) );
  ANDN U44305 ( .B(n42988), .A(n42989), .Z(n42986) );
  AND U44306 ( .A(a[1]), .B(b[39]), .Z(n42985) );
  XOR U44307 ( .A(n42991), .B(n42992), .Z(n42756) );
  ANDN U44308 ( .B(n42993), .A(n42994), .Z(n42991) );
  AND U44309 ( .A(a[2]), .B(b[38]), .Z(n42990) );
  XOR U44310 ( .A(n42996), .B(n42997), .Z(n42761) );
  ANDN U44311 ( .B(n42998), .A(n42999), .Z(n42996) );
  AND U44312 ( .A(a[3]), .B(b[37]), .Z(n42995) );
  XOR U44313 ( .A(n43001), .B(n43002), .Z(n42766) );
  ANDN U44314 ( .B(n43003), .A(n43004), .Z(n43001) );
  AND U44315 ( .A(a[4]), .B(b[36]), .Z(n43000) );
  XOR U44316 ( .A(n43006), .B(n43007), .Z(n42771) );
  ANDN U44317 ( .B(n43008), .A(n43009), .Z(n43006) );
  AND U44318 ( .A(a[5]), .B(b[35]), .Z(n43005) );
  XOR U44319 ( .A(n43011), .B(n43012), .Z(n42776) );
  ANDN U44320 ( .B(n43013), .A(n43014), .Z(n43011) );
  AND U44321 ( .A(a[6]), .B(b[34]), .Z(n43010) );
  XOR U44322 ( .A(n43016), .B(n43017), .Z(n42781) );
  ANDN U44323 ( .B(n43018), .A(n43019), .Z(n43016) );
  AND U44324 ( .A(a[7]), .B(b[33]), .Z(n43015) );
  XOR U44325 ( .A(n43021), .B(n43022), .Z(n42786) );
  ANDN U44326 ( .B(n43023), .A(n43024), .Z(n43021) );
  AND U44327 ( .A(a[8]), .B(b[32]), .Z(n43020) );
  XOR U44328 ( .A(n43026), .B(n43027), .Z(n42791) );
  ANDN U44329 ( .B(n43028), .A(n43029), .Z(n43026) );
  AND U44330 ( .A(a[9]), .B(b[31]), .Z(n43025) );
  XOR U44331 ( .A(n43031), .B(n43032), .Z(n42796) );
  ANDN U44332 ( .B(n43033), .A(n43034), .Z(n43031) );
  AND U44333 ( .A(a[10]), .B(b[30]), .Z(n43030) );
  XOR U44334 ( .A(n43036), .B(n43037), .Z(n42801) );
  ANDN U44335 ( .B(n43038), .A(n43039), .Z(n43036) );
  AND U44336 ( .A(a[11]), .B(b[29]), .Z(n43035) );
  XOR U44337 ( .A(n43041), .B(n43042), .Z(n42806) );
  ANDN U44338 ( .B(n43043), .A(n43044), .Z(n43041) );
  AND U44339 ( .A(a[12]), .B(b[28]), .Z(n43040) );
  XOR U44340 ( .A(n43046), .B(n43047), .Z(n42811) );
  ANDN U44341 ( .B(n43048), .A(n43049), .Z(n43046) );
  AND U44342 ( .A(a[13]), .B(b[27]), .Z(n43045) );
  XOR U44343 ( .A(n43051), .B(n43052), .Z(n42816) );
  ANDN U44344 ( .B(n43053), .A(n43054), .Z(n43051) );
  AND U44345 ( .A(a[14]), .B(b[26]), .Z(n43050) );
  XOR U44346 ( .A(n43056), .B(n43057), .Z(n42821) );
  ANDN U44347 ( .B(n43058), .A(n43059), .Z(n43056) );
  AND U44348 ( .A(a[15]), .B(b[25]), .Z(n43055) );
  XOR U44349 ( .A(n43061), .B(n43062), .Z(n42826) );
  ANDN U44350 ( .B(n43063), .A(n43064), .Z(n43061) );
  AND U44351 ( .A(a[16]), .B(b[24]), .Z(n43060) );
  XOR U44352 ( .A(n43066), .B(n43067), .Z(n42831) );
  ANDN U44353 ( .B(n43068), .A(n43069), .Z(n43066) );
  AND U44354 ( .A(a[17]), .B(b[23]), .Z(n43065) );
  XOR U44355 ( .A(n43071), .B(n43072), .Z(n42836) );
  ANDN U44356 ( .B(n43073), .A(n43074), .Z(n43071) );
  AND U44357 ( .A(a[18]), .B(b[22]), .Z(n43070) );
  XOR U44358 ( .A(n43076), .B(n43077), .Z(n42841) );
  ANDN U44359 ( .B(n43078), .A(n43079), .Z(n43076) );
  AND U44360 ( .A(a[19]), .B(b[21]), .Z(n43075) );
  XOR U44361 ( .A(n43081), .B(n43082), .Z(n42846) );
  ANDN U44362 ( .B(n43083), .A(n43084), .Z(n43081) );
  AND U44363 ( .A(a[20]), .B(b[20]), .Z(n43080) );
  XOR U44364 ( .A(n43086), .B(n43087), .Z(n42851) );
  ANDN U44365 ( .B(n43088), .A(n43089), .Z(n43086) );
  AND U44366 ( .A(a[21]), .B(b[19]), .Z(n43085) );
  XOR U44367 ( .A(n43091), .B(n43092), .Z(n42856) );
  ANDN U44368 ( .B(n43093), .A(n43094), .Z(n43091) );
  AND U44369 ( .A(a[22]), .B(b[18]), .Z(n43090) );
  XOR U44370 ( .A(n43096), .B(n43097), .Z(n42861) );
  ANDN U44371 ( .B(n43098), .A(n43099), .Z(n43096) );
  AND U44372 ( .A(a[23]), .B(b[17]), .Z(n43095) );
  XOR U44373 ( .A(n43101), .B(n43102), .Z(n42866) );
  ANDN U44374 ( .B(n43103), .A(n43104), .Z(n43101) );
  AND U44375 ( .A(a[24]), .B(b[16]), .Z(n43100) );
  XOR U44376 ( .A(n43106), .B(n43107), .Z(n42871) );
  ANDN U44377 ( .B(n43108), .A(n43109), .Z(n43106) );
  AND U44378 ( .A(a[25]), .B(b[15]), .Z(n43105) );
  XOR U44379 ( .A(n43111), .B(n43112), .Z(n42876) );
  ANDN U44380 ( .B(n43113), .A(n43114), .Z(n43111) );
  AND U44381 ( .A(a[26]), .B(b[14]), .Z(n43110) );
  XOR U44382 ( .A(n43116), .B(n43117), .Z(n42881) );
  ANDN U44383 ( .B(n43118), .A(n43119), .Z(n43116) );
  AND U44384 ( .A(a[27]), .B(b[13]), .Z(n43115) );
  XOR U44385 ( .A(n43121), .B(n43122), .Z(n42886) );
  ANDN U44386 ( .B(n43123), .A(n43124), .Z(n43121) );
  AND U44387 ( .A(a[28]), .B(b[12]), .Z(n43120) );
  XOR U44388 ( .A(n43126), .B(n43127), .Z(n42891) );
  ANDN U44389 ( .B(n43128), .A(n43129), .Z(n43126) );
  AND U44390 ( .A(a[29]), .B(b[11]), .Z(n43125) );
  XOR U44391 ( .A(n43131), .B(n43132), .Z(n42896) );
  ANDN U44392 ( .B(n43133), .A(n43134), .Z(n43131) );
  AND U44393 ( .A(a[30]), .B(b[10]), .Z(n43130) );
  XOR U44394 ( .A(n43136), .B(n43137), .Z(n42901) );
  ANDN U44395 ( .B(n43138), .A(n43139), .Z(n43136) );
  AND U44396 ( .A(b[9]), .B(a[31]), .Z(n43135) );
  XOR U44397 ( .A(n43141), .B(n43142), .Z(n42906) );
  ANDN U44398 ( .B(n43143), .A(n43144), .Z(n43141) );
  AND U44399 ( .A(b[8]), .B(a[32]), .Z(n43140) );
  XOR U44400 ( .A(n43146), .B(n43147), .Z(n42911) );
  ANDN U44401 ( .B(n43148), .A(n43149), .Z(n43146) );
  AND U44402 ( .A(b[7]), .B(a[33]), .Z(n43145) );
  XOR U44403 ( .A(n43151), .B(n43152), .Z(n42916) );
  ANDN U44404 ( .B(n43153), .A(n43154), .Z(n43151) );
  AND U44405 ( .A(b[6]), .B(a[34]), .Z(n43150) );
  XOR U44406 ( .A(n43156), .B(n43157), .Z(n42921) );
  ANDN U44407 ( .B(n43158), .A(n43159), .Z(n43156) );
  AND U44408 ( .A(b[5]), .B(a[35]), .Z(n43155) );
  XOR U44409 ( .A(n43161), .B(n43162), .Z(n42926) );
  ANDN U44410 ( .B(n43163), .A(n43164), .Z(n43161) );
  AND U44411 ( .A(b[4]), .B(a[36]), .Z(n43160) );
  XOR U44412 ( .A(n43166), .B(n43167), .Z(n42931) );
  ANDN U44413 ( .B(n42943), .A(n42944), .Z(n43166) );
  AND U44414 ( .A(b[2]), .B(a[37]), .Z(n43168) );
  XNOR U44415 ( .A(n43163), .B(n43167), .Z(n43169) );
  XOR U44416 ( .A(n43170), .B(n43171), .Z(n43167) );
  OR U44417 ( .A(n42946), .B(n42947), .Z(n43171) );
  XNOR U44418 ( .A(n43173), .B(n43174), .Z(n43172) );
  XOR U44419 ( .A(n43173), .B(n43176), .Z(n42946) );
  NAND U44420 ( .A(b[1]), .B(a[37]), .Z(n43176) );
  IV U44421 ( .A(n43170), .Z(n43173) );
  NANDN U44422 ( .A(n139), .B(n140), .Z(n43170) );
  XOR U44423 ( .A(n43177), .B(n43178), .Z(n140) );
  NAND U44424 ( .A(a[37]), .B(b[0]), .Z(n139) );
  XNOR U44425 ( .A(n43158), .B(n43162), .Z(n43179) );
  XNOR U44426 ( .A(n43153), .B(n43157), .Z(n43180) );
  XNOR U44427 ( .A(n43148), .B(n43152), .Z(n43181) );
  XNOR U44428 ( .A(n43143), .B(n43147), .Z(n43182) );
  XNOR U44429 ( .A(n43138), .B(n43142), .Z(n43183) );
  XNOR U44430 ( .A(n43133), .B(n43137), .Z(n43184) );
  XNOR U44431 ( .A(n43128), .B(n43132), .Z(n43185) );
  XNOR U44432 ( .A(n43123), .B(n43127), .Z(n43186) );
  XNOR U44433 ( .A(n43118), .B(n43122), .Z(n43187) );
  XNOR U44434 ( .A(n43113), .B(n43117), .Z(n43188) );
  XNOR U44435 ( .A(n43108), .B(n43112), .Z(n43189) );
  XNOR U44436 ( .A(n43103), .B(n43107), .Z(n43190) );
  XNOR U44437 ( .A(n43098), .B(n43102), .Z(n43191) );
  XNOR U44438 ( .A(n43093), .B(n43097), .Z(n43192) );
  XNOR U44439 ( .A(n43088), .B(n43092), .Z(n43193) );
  XNOR U44440 ( .A(n43083), .B(n43087), .Z(n43194) );
  XNOR U44441 ( .A(n43078), .B(n43082), .Z(n43195) );
  XNOR U44442 ( .A(n43073), .B(n43077), .Z(n43196) );
  XNOR U44443 ( .A(n43068), .B(n43072), .Z(n43197) );
  XNOR U44444 ( .A(n43063), .B(n43067), .Z(n43198) );
  XNOR U44445 ( .A(n43058), .B(n43062), .Z(n43199) );
  XNOR U44446 ( .A(n43053), .B(n43057), .Z(n43200) );
  XNOR U44447 ( .A(n43048), .B(n43052), .Z(n43201) );
  XNOR U44448 ( .A(n43043), .B(n43047), .Z(n43202) );
  XNOR U44449 ( .A(n43038), .B(n43042), .Z(n43203) );
  XNOR U44450 ( .A(n43033), .B(n43037), .Z(n43204) );
  XNOR U44451 ( .A(n43028), .B(n43032), .Z(n43205) );
  XNOR U44452 ( .A(n43023), .B(n43027), .Z(n43206) );
  XNOR U44453 ( .A(n43018), .B(n43022), .Z(n43207) );
  XNOR U44454 ( .A(n43013), .B(n43017), .Z(n43208) );
  XNOR U44455 ( .A(n43008), .B(n43012), .Z(n43209) );
  XNOR U44456 ( .A(n43003), .B(n43007), .Z(n43210) );
  XNOR U44457 ( .A(n42998), .B(n43002), .Z(n43211) );
  XNOR U44458 ( .A(n42993), .B(n42997), .Z(n43212) );
  XNOR U44459 ( .A(n42988), .B(n42992), .Z(n43213) );
  XNOR U44460 ( .A(n43214), .B(n42987), .Z(n42988) );
  AND U44461 ( .A(a[0]), .B(b[39]), .Z(n43214) );
  XOR U44462 ( .A(n43215), .B(n42987), .Z(n42989) );
  XNOR U44463 ( .A(n43216), .B(n43217), .Z(n42987) );
  ANDN U44464 ( .B(n43218), .A(n43219), .Z(n43216) );
  AND U44465 ( .A(a[1]), .B(b[38]), .Z(n43215) );
  XOR U44466 ( .A(n43221), .B(n43222), .Z(n42992) );
  ANDN U44467 ( .B(n43223), .A(n43224), .Z(n43221) );
  AND U44468 ( .A(a[2]), .B(b[37]), .Z(n43220) );
  XOR U44469 ( .A(n43226), .B(n43227), .Z(n42997) );
  ANDN U44470 ( .B(n43228), .A(n43229), .Z(n43226) );
  AND U44471 ( .A(a[3]), .B(b[36]), .Z(n43225) );
  XOR U44472 ( .A(n43231), .B(n43232), .Z(n43002) );
  ANDN U44473 ( .B(n43233), .A(n43234), .Z(n43231) );
  AND U44474 ( .A(a[4]), .B(b[35]), .Z(n43230) );
  XOR U44475 ( .A(n43236), .B(n43237), .Z(n43007) );
  ANDN U44476 ( .B(n43238), .A(n43239), .Z(n43236) );
  AND U44477 ( .A(a[5]), .B(b[34]), .Z(n43235) );
  XOR U44478 ( .A(n43241), .B(n43242), .Z(n43012) );
  ANDN U44479 ( .B(n43243), .A(n43244), .Z(n43241) );
  AND U44480 ( .A(a[6]), .B(b[33]), .Z(n43240) );
  XOR U44481 ( .A(n43246), .B(n43247), .Z(n43017) );
  ANDN U44482 ( .B(n43248), .A(n43249), .Z(n43246) );
  AND U44483 ( .A(a[7]), .B(b[32]), .Z(n43245) );
  XOR U44484 ( .A(n43251), .B(n43252), .Z(n43022) );
  ANDN U44485 ( .B(n43253), .A(n43254), .Z(n43251) );
  AND U44486 ( .A(a[8]), .B(b[31]), .Z(n43250) );
  XOR U44487 ( .A(n43256), .B(n43257), .Z(n43027) );
  ANDN U44488 ( .B(n43258), .A(n43259), .Z(n43256) );
  AND U44489 ( .A(a[9]), .B(b[30]), .Z(n43255) );
  XOR U44490 ( .A(n43261), .B(n43262), .Z(n43032) );
  ANDN U44491 ( .B(n43263), .A(n43264), .Z(n43261) );
  AND U44492 ( .A(a[10]), .B(b[29]), .Z(n43260) );
  XOR U44493 ( .A(n43266), .B(n43267), .Z(n43037) );
  ANDN U44494 ( .B(n43268), .A(n43269), .Z(n43266) );
  AND U44495 ( .A(a[11]), .B(b[28]), .Z(n43265) );
  XOR U44496 ( .A(n43271), .B(n43272), .Z(n43042) );
  ANDN U44497 ( .B(n43273), .A(n43274), .Z(n43271) );
  AND U44498 ( .A(a[12]), .B(b[27]), .Z(n43270) );
  XOR U44499 ( .A(n43276), .B(n43277), .Z(n43047) );
  ANDN U44500 ( .B(n43278), .A(n43279), .Z(n43276) );
  AND U44501 ( .A(a[13]), .B(b[26]), .Z(n43275) );
  XOR U44502 ( .A(n43281), .B(n43282), .Z(n43052) );
  ANDN U44503 ( .B(n43283), .A(n43284), .Z(n43281) );
  AND U44504 ( .A(a[14]), .B(b[25]), .Z(n43280) );
  XOR U44505 ( .A(n43286), .B(n43287), .Z(n43057) );
  ANDN U44506 ( .B(n43288), .A(n43289), .Z(n43286) );
  AND U44507 ( .A(a[15]), .B(b[24]), .Z(n43285) );
  XOR U44508 ( .A(n43291), .B(n43292), .Z(n43062) );
  ANDN U44509 ( .B(n43293), .A(n43294), .Z(n43291) );
  AND U44510 ( .A(a[16]), .B(b[23]), .Z(n43290) );
  XOR U44511 ( .A(n43296), .B(n43297), .Z(n43067) );
  ANDN U44512 ( .B(n43298), .A(n43299), .Z(n43296) );
  AND U44513 ( .A(a[17]), .B(b[22]), .Z(n43295) );
  XOR U44514 ( .A(n43301), .B(n43302), .Z(n43072) );
  ANDN U44515 ( .B(n43303), .A(n43304), .Z(n43301) );
  AND U44516 ( .A(a[18]), .B(b[21]), .Z(n43300) );
  XOR U44517 ( .A(n43306), .B(n43307), .Z(n43077) );
  ANDN U44518 ( .B(n43308), .A(n43309), .Z(n43306) );
  AND U44519 ( .A(a[19]), .B(b[20]), .Z(n43305) );
  XOR U44520 ( .A(n43311), .B(n43312), .Z(n43082) );
  ANDN U44521 ( .B(n43313), .A(n43314), .Z(n43311) );
  AND U44522 ( .A(a[20]), .B(b[19]), .Z(n43310) );
  XOR U44523 ( .A(n43316), .B(n43317), .Z(n43087) );
  ANDN U44524 ( .B(n43318), .A(n43319), .Z(n43316) );
  AND U44525 ( .A(a[21]), .B(b[18]), .Z(n43315) );
  XOR U44526 ( .A(n43321), .B(n43322), .Z(n43092) );
  ANDN U44527 ( .B(n43323), .A(n43324), .Z(n43321) );
  AND U44528 ( .A(a[22]), .B(b[17]), .Z(n43320) );
  XOR U44529 ( .A(n43326), .B(n43327), .Z(n43097) );
  ANDN U44530 ( .B(n43328), .A(n43329), .Z(n43326) );
  AND U44531 ( .A(a[23]), .B(b[16]), .Z(n43325) );
  XOR U44532 ( .A(n43331), .B(n43332), .Z(n43102) );
  ANDN U44533 ( .B(n43333), .A(n43334), .Z(n43331) );
  AND U44534 ( .A(a[24]), .B(b[15]), .Z(n43330) );
  XOR U44535 ( .A(n43336), .B(n43337), .Z(n43107) );
  ANDN U44536 ( .B(n43338), .A(n43339), .Z(n43336) );
  AND U44537 ( .A(a[25]), .B(b[14]), .Z(n43335) );
  XOR U44538 ( .A(n43341), .B(n43342), .Z(n43112) );
  ANDN U44539 ( .B(n43343), .A(n43344), .Z(n43341) );
  AND U44540 ( .A(a[26]), .B(b[13]), .Z(n43340) );
  XOR U44541 ( .A(n43346), .B(n43347), .Z(n43117) );
  ANDN U44542 ( .B(n43348), .A(n43349), .Z(n43346) );
  AND U44543 ( .A(a[27]), .B(b[12]), .Z(n43345) );
  XOR U44544 ( .A(n43351), .B(n43352), .Z(n43122) );
  ANDN U44545 ( .B(n43353), .A(n43354), .Z(n43351) );
  AND U44546 ( .A(a[28]), .B(b[11]), .Z(n43350) );
  XOR U44547 ( .A(n43356), .B(n43357), .Z(n43127) );
  ANDN U44548 ( .B(n43358), .A(n43359), .Z(n43356) );
  AND U44549 ( .A(a[29]), .B(b[10]), .Z(n43355) );
  XOR U44550 ( .A(n43361), .B(n43362), .Z(n43132) );
  ANDN U44551 ( .B(n43363), .A(n43364), .Z(n43361) );
  AND U44552 ( .A(b[9]), .B(a[30]), .Z(n43360) );
  XOR U44553 ( .A(n43366), .B(n43367), .Z(n43137) );
  ANDN U44554 ( .B(n43368), .A(n43369), .Z(n43366) );
  AND U44555 ( .A(b[8]), .B(a[31]), .Z(n43365) );
  XOR U44556 ( .A(n43371), .B(n43372), .Z(n43142) );
  ANDN U44557 ( .B(n43373), .A(n43374), .Z(n43371) );
  AND U44558 ( .A(b[7]), .B(a[32]), .Z(n43370) );
  XOR U44559 ( .A(n43376), .B(n43377), .Z(n43147) );
  ANDN U44560 ( .B(n43378), .A(n43379), .Z(n43376) );
  AND U44561 ( .A(b[6]), .B(a[33]), .Z(n43375) );
  XOR U44562 ( .A(n43381), .B(n43382), .Z(n43152) );
  ANDN U44563 ( .B(n43383), .A(n43384), .Z(n43381) );
  AND U44564 ( .A(b[5]), .B(a[34]), .Z(n43380) );
  XOR U44565 ( .A(n43386), .B(n43387), .Z(n43157) );
  ANDN U44566 ( .B(n43388), .A(n43389), .Z(n43386) );
  AND U44567 ( .A(b[4]), .B(a[35]), .Z(n43385) );
  XOR U44568 ( .A(n43391), .B(n43392), .Z(n43162) );
  ANDN U44569 ( .B(n43174), .A(n43175), .Z(n43391) );
  AND U44570 ( .A(b[2]), .B(a[36]), .Z(n43393) );
  XNOR U44571 ( .A(n43388), .B(n43392), .Z(n43394) );
  XOR U44572 ( .A(n43395), .B(n43396), .Z(n43392) );
  OR U44573 ( .A(n43177), .B(n43178), .Z(n43396) );
  XNOR U44574 ( .A(n43398), .B(n43399), .Z(n43397) );
  XOR U44575 ( .A(n43398), .B(n43401), .Z(n43177) );
  NAND U44576 ( .A(b[1]), .B(a[36]), .Z(n43401) );
  IV U44577 ( .A(n43395), .Z(n43398) );
  NANDN U44578 ( .A(n141), .B(n142), .Z(n43395) );
  XOR U44579 ( .A(n43402), .B(n43403), .Z(n142) );
  NAND U44580 ( .A(a[36]), .B(b[0]), .Z(n141) );
  XNOR U44581 ( .A(n43383), .B(n43387), .Z(n43404) );
  XNOR U44582 ( .A(n43378), .B(n43382), .Z(n43405) );
  XNOR U44583 ( .A(n43373), .B(n43377), .Z(n43406) );
  XNOR U44584 ( .A(n43368), .B(n43372), .Z(n43407) );
  XNOR U44585 ( .A(n43363), .B(n43367), .Z(n43408) );
  XNOR U44586 ( .A(n43358), .B(n43362), .Z(n43409) );
  XNOR U44587 ( .A(n43353), .B(n43357), .Z(n43410) );
  XNOR U44588 ( .A(n43348), .B(n43352), .Z(n43411) );
  XNOR U44589 ( .A(n43343), .B(n43347), .Z(n43412) );
  XNOR U44590 ( .A(n43338), .B(n43342), .Z(n43413) );
  XNOR U44591 ( .A(n43333), .B(n43337), .Z(n43414) );
  XNOR U44592 ( .A(n43328), .B(n43332), .Z(n43415) );
  XNOR U44593 ( .A(n43323), .B(n43327), .Z(n43416) );
  XNOR U44594 ( .A(n43318), .B(n43322), .Z(n43417) );
  XNOR U44595 ( .A(n43313), .B(n43317), .Z(n43418) );
  XNOR U44596 ( .A(n43308), .B(n43312), .Z(n43419) );
  XNOR U44597 ( .A(n43303), .B(n43307), .Z(n43420) );
  XNOR U44598 ( .A(n43298), .B(n43302), .Z(n43421) );
  XNOR U44599 ( .A(n43293), .B(n43297), .Z(n43422) );
  XNOR U44600 ( .A(n43288), .B(n43292), .Z(n43423) );
  XNOR U44601 ( .A(n43283), .B(n43287), .Z(n43424) );
  XNOR U44602 ( .A(n43278), .B(n43282), .Z(n43425) );
  XNOR U44603 ( .A(n43273), .B(n43277), .Z(n43426) );
  XNOR U44604 ( .A(n43268), .B(n43272), .Z(n43427) );
  XNOR U44605 ( .A(n43263), .B(n43267), .Z(n43428) );
  XNOR U44606 ( .A(n43258), .B(n43262), .Z(n43429) );
  XNOR U44607 ( .A(n43253), .B(n43257), .Z(n43430) );
  XNOR U44608 ( .A(n43248), .B(n43252), .Z(n43431) );
  XNOR U44609 ( .A(n43243), .B(n43247), .Z(n43432) );
  XNOR U44610 ( .A(n43238), .B(n43242), .Z(n43433) );
  XNOR U44611 ( .A(n43233), .B(n43237), .Z(n43434) );
  XNOR U44612 ( .A(n43228), .B(n43232), .Z(n43435) );
  XNOR U44613 ( .A(n43223), .B(n43227), .Z(n43436) );
  XNOR U44614 ( .A(n43218), .B(n43222), .Z(n43437) );
  XOR U44615 ( .A(n43438), .B(n43217), .Z(n43218) );
  AND U44616 ( .A(a[0]), .B(b[38]), .Z(n43438) );
  XNOR U44617 ( .A(n43439), .B(n43217), .Z(n43219) );
  XNOR U44618 ( .A(n43440), .B(n43441), .Z(n43217) );
  ANDN U44619 ( .B(n43442), .A(n43443), .Z(n43440) );
  AND U44620 ( .A(a[1]), .B(b[37]), .Z(n43439) );
  XOR U44621 ( .A(n43445), .B(n43446), .Z(n43222) );
  ANDN U44622 ( .B(n43447), .A(n43448), .Z(n43445) );
  AND U44623 ( .A(a[2]), .B(b[36]), .Z(n43444) );
  XOR U44624 ( .A(n43450), .B(n43451), .Z(n43227) );
  ANDN U44625 ( .B(n43452), .A(n43453), .Z(n43450) );
  AND U44626 ( .A(a[3]), .B(b[35]), .Z(n43449) );
  XOR U44627 ( .A(n43455), .B(n43456), .Z(n43232) );
  ANDN U44628 ( .B(n43457), .A(n43458), .Z(n43455) );
  AND U44629 ( .A(a[4]), .B(b[34]), .Z(n43454) );
  XOR U44630 ( .A(n43460), .B(n43461), .Z(n43237) );
  ANDN U44631 ( .B(n43462), .A(n43463), .Z(n43460) );
  AND U44632 ( .A(a[5]), .B(b[33]), .Z(n43459) );
  XOR U44633 ( .A(n43465), .B(n43466), .Z(n43242) );
  ANDN U44634 ( .B(n43467), .A(n43468), .Z(n43465) );
  AND U44635 ( .A(a[6]), .B(b[32]), .Z(n43464) );
  XOR U44636 ( .A(n43470), .B(n43471), .Z(n43247) );
  ANDN U44637 ( .B(n43472), .A(n43473), .Z(n43470) );
  AND U44638 ( .A(a[7]), .B(b[31]), .Z(n43469) );
  XOR U44639 ( .A(n43475), .B(n43476), .Z(n43252) );
  ANDN U44640 ( .B(n43477), .A(n43478), .Z(n43475) );
  AND U44641 ( .A(a[8]), .B(b[30]), .Z(n43474) );
  XOR U44642 ( .A(n43480), .B(n43481), .Z(n43257) );
  ANDN U44643 ( .B(n43482), .A(n43483), .Z(n43480) );
  AND U44644 ( .A(a[9]), .B(b[29]), .Z(n43479) );
  XOR U44645 ( .A(n43485), .B(n43486), .Z(n43262) );
  ANDN U44646 ( .B(n43487), .A(n43488), .Z(n43485) );
  AND U44647 ( .A(a[10]), .B(b[28]), .Z(n43484) );
  XOR U44648 ( .A(n43490), .B(n43491), .Z(n43267) );
  ANDN U44649 ( .B(n43492), .A(n43493), .Z(n43490) );
  AND U44650 ( .A(a[11]), .B(b[27]), .Z(n43489) );
  XOR U44651 ( .A(n43495), .B(n43496), .Z(n43272) );
  ANDN U44652 ( .B(n43497), .A(n43498), .Z(n43495) );
  AND U44653 ( .A(a[12]), .B(b[26]), .Z(n43494) );
  XOR U44654 ( .A(n43500), .B(n43501), .Z(n43277) );
  ANDN U44655 ( .B(n43502), .A(n43503), .Z(n43500) );
  AND U44656 ( .A(a[13]), .B(b[25]), .Z(n43499) );
  XOR U44657 ( .A(n43505), .B(n43506), .Z(n43282) );
  ANDN U44658 ( .B(n43507), .A(n43508), .Z(n43505) );
  AND U44659 ( .A(a[14]), .B(b[24]), .Z(n43504) );
  XOR U44660 ( .A(n43510), .B(n43511), .Z(n43287) );
  ANDN U44661 ( .B(n43512), .A(n43513), .Z(n43510) );
  AND U44662 ( .A(a[15]), .B(b[23]), .Z(n43509) );
  XOR U44663 ( .A(n43515), .B(n43516), .Z(n43292) );
  ANDN U44664 ( .B(n43517), .A(n43518), .Z(n43515) );
  AND U44665 ( .A(a[16]), .B(b[22]), .Z(n43514) );
  XOR U44666 ( .A(n43520), .B(n43521), .Z(n43297) );
  ANDN U44667 ( .B(n43522), .A(n43523), .Z(n43520) );
  AND U44668 ( .A(a[17]), .B(b[21]), .Z(n43519) );
  XOR U44669 ( .A(n43525), .B(n43526), .Z(n43302) );
  ANDN U44670 ( .B(n43527), .A(n43528), .Z(n43525) );
  AND U44671 ( .A(a[18]), .B(b[20]), .Z(n43524) );
  XOR U44672 ( .A(n43530), .B(n43531), .Z(n43307) );
  ANDN U44673 ( .B(n43532), .A(n43533), .Z(n43530) );
  AND U44674 ( .A(a[19]), .B(b[19]), .Z(n43529) );
  XOR U44675 ( .A(n43535), .B(n43536), .Z(n43312) );
  ANDN U44676 ( .B(n43537), .A(n43538), .Z(n43535) );
  AND U44677 ( .A(a[20]), .B(b[18]), .Z(n43534) );
  XOR U44678 ( .A(n43540), .B(n43541), .Z(n43317) );
  ANDN U44679 ( .B(n43542), .A(n43543), .Z(n43540) );
  AND U44680 ( .A(a[21]), .B(b[17]), .Z(n43539) );
  XOR U44681 ( .A(n43545), .B(n43546), .Z(n43322) );
  ANDN U44682 ( .B(n43547), .A(n43548), .Z(n43545) );
  AND U44683 ( .A(a[22]), .B(b[16]), .Z(n43544) );
  XOR U44684 ( .A(n43550), .B(n43551), .Z(n43327) );
  ANDN U44685 ( .B(n43552), .A(n43553), .Z(n43550) );
  AND U44686 ( .A(a[23]), .B(b[15]), .Z(n43549) );
  XOR U44687 ( .A(n43555), .B(n43556), .Z(n43332) );
  ANDN U44688 ( .B(n43557), .A(n43558), .Z(n43555) );
  AND U44689 ( .A(a[24]), .B(b[14]), .Z(n43554) );
  XOR U44690 ( .A(n43560), .B(n43561), .Z(n43337) );
  ANDN U44691 ( .B(n43562), .A(n43563), .Z(n43560) );
  AND U44692 ( .A(a[25]), .B(b[13]), .Z(n43559) );
  XOR U44693 ( .A(n43565), .B(n43566), .Z(n43342) );
  ANDN U44694 ( .B(n43567), .A(n43568), .Z(n43565) );
  AND U44695 ( .A(a[26]), .B(b[12]), .Z(n43564) );
  XOR U44696 ( .A(n43570), .B(n43571), .Z(n43347) );
  ANDN U44697 ( .B(n43572), .A(n43573), .Z(n43570) );
  AND U44698 ( .A(a[27]), .B(b[11]), .Z(n43569) );
  XOR U44699 ( .A(n43575), .B(n43576), .Z(n43352) );
  ANDN U44700 ( .B(n43577), .A(n43578), .Z(n43575) );
  AND U44701 ( .A(a[28]), .B(b[10]), .Z(n43574) );
  XOR U44702 ( .A(n43580), .B(n43581), .Z(n43357) );
  ANDN U44703 ( .B(n43582), .A(n43583), .Z(n43580) );
  AND U44704 ( .A(b[9]), .B(a[29]), .Z(n43579) );
  XOR U44705 ( .A(n43585), .B(n43586), .Z(n43362) );
  ANDN U44706 ( .B(n43587), .A(n43588), .Z(n43585) );
  AND U44707 ( .A(b[8]), .B(a[30]), .Z(n43584) );
  XOR U44708 ( .A(n43590), .B(n43591), .Z(n43367) );
  ANDN U44709 ( .B(n43592), .A(n43593), .Z(n43590) );
  AND U44710 ( .A(b[7]), .B(a[31]), .Z(n43589) );
  XOR U44711 ( .A(n43595), .B(n43596), .Z(n43372) );
  ANDN U44712 ( .B(n43597), .A(n43598), .Z(n43595) );
  AND U44713 ( .A(b[6]), .B(a[32]), .Z(n43594) );
  XOR U44714 ( .A(n43600), .B(n43601), .Z(n43377) );
  ANDN U44715 ( .B(n43602), .A(n43603), .Z(n43600) );
  AND U44716 ( .A(b[5]), .B(a[33]), .Z(n43599) );
  XOR U44717 ( .A(n43605), .B(n43606), .Z(n43382) );
  ANDN U44718 ( .B(n43607), .A(n43608), .Z(n43605) );
  AND U44719 ( .A(b[4]), .B(a[34]), .Z(n43604) );
  XOR U44720 ( .A(n43610), .B(n43611), .Z(n43387) );
  ANDN U44721 ( .B(n43399), .A(n43400), .Z(n43610) );
  AND U44722 ( .A(b[2]), .B(a[35]), .Z(n43612) );
  XNOR U44723 ( .A(n43607), .B(n43611), .Z(n43613) );
  XOR U44724 ( .A(n43614), .B(n43615), .Z(n43611) );
  OR U44725 ( .A(n43402), .B(n43403), .Z(n43615) );
  XNOR U44726 ( .A(n43617), .B(n43618), .Z(n43616) );
  XOR U44727 ( .A(n43617), .B(n43620), .Z(n43402) );
  NAND U44728 ( .A(b[1]), .B(a[35]), .Z(n43620) );
  IV U44729 ( .A(n43614), .Z(n43617) );
  NANDN U44730 ( .A(n143), .B(n144), .Z(n43614) );
  XOR U44731 ( .A(n43621), .B(n43622), .Z(n144) );
  NAND U44732 ( .A(a[35]), .B(b[0]), .Z(n143) );
  XNOR U44733 ( .A(n43602), .B(n43606), .Z(n43623) );
  XNOR U44734 ( .A(n43597), .B(n43601), .Z(n43624) );
  XNOR U44735 ( .A(n43592), .B(n43596), .Z(n43625) );
  XNOR U44736 ( .A(n43587), .B(n43591), .Z(n43626) );
  XNOR U44737 ( .A(n43582), .B(n43586), .Z(n43627) );
  XNOR U44738 ( .A(n43577), .B(n43581), .Z(n43628) );
  XNOR U44739 ( .A(n43572), .B(n43576), .Z(n43629) );
  XNOR U44740 ( .A(n43567), .B(n43571), .Z(n43630) );
  XNOR U44741 ( .A(n43562), .B(n43566), .Z(n43631) );
  XNOR U44742 ( .A(n43557), .B(n43561), .Z(n43632) );
  XNOR U44743 ( .A(n43552), .B(n43556), .Z(n43633) );
  XNOR U44744 ( .A(n43547), .B(n43551), .Z(n43634) );
  XNOR U44745 ( .A(n43542), .B(n43546), .Z(n43635) );
  XNOR U44746 ( .A(n43537), .B(n43541), .Z(n43636) );
  XNOR U44747 ( .A(n43532), .B(n43536), .Z(n43637) );
  XNOR U44748 ( .A(n43527), .B(n43531), .Z(n43638) );
  XNOR U44749 ( .A(n43522), .B(n43526), .Z(n43639) );
  XNOR U44750 ( .A(n43517), .B(n43521), .Z(n43640) );
  XNOR U44751 ( .A(n43512), .B(n43516), .Z(n43641) );
  XNOR U44752 ( .A(n43507), .B(n43511), .Z(n43642) );
  XNOR U44753 ( .A(n43502), .B(n43506), .Z(n43643) );
  XNOR U44754 ( .A(n43497), .B(n43501), .Z(n43644) );
  XNOR U44755 ( .A(n43492), .B(n43496), .Z(n43645) );
  XNOR U44756 ( .A(n43487), .B(n43491), .Z(n43646) );
  XNOR U44757 ( .A(n43482), .B(n43486), .Z(n43647) );
  XNOR U44758 ( .A(n43477), .B(n43481), .Z(n43648) );
  XNOR U44759 ( .A(n43472), .B(n43476), .Z(n43649) );
  XNOR U44760 ( .A(n43467), .B(n43471), .Z(n43650) );
  XNOR U44761 ( .A(n43462), .B(n43466), .Z(n43651) );
  XNOR U44762 ( .A(n43457), .B(n43461), .Z(n43652) );
  XNOR U44763 ( .A(n43452), .B(n43456), .Z(n43653) );
  XNOR U44764 ( .A(n43447), .B(n43451), .Z(n43654) );
  XNOR U44765 ( .A(n43442), .B(n43446), .Z(n43655) );
  XNOR U44766 ( .A(n43656), .B(n43441), .Z(n43442) );
  AND U44767 ( .A(a[0]), .B(b[37]), .Z(n43656) );
  XOR U44768 ( .A(n43657), .B(n43441), .Z(n43443) );
  XNOR U44769 ( .A(n43658), .B(n43659), .Z(n43441) );
  ANDN U44770 ( .B(n43660), .A(n43661), .Z(n43658) );
  AND U44771 ( .A(a[1]), .B(b[36]), .Z(n43657) );
  XOR U44772 ( .A(n43663), .B(n43664), .Z(n43446) );
  ANDN U44773 ( .B(n43665), .A(n43666), .Z(n43663) );
  AND U44774 ( .A(a[2]), .B(b[35]), .Z(n43662) );
  XOR U44775 ( .A(n43668), .B(n43669), .Z(n43451) );
  ANDN U44776 ( .B(n43670), .A(n43671), .Z(n43668) );
  AND U44777 ( .A(a[3]), .B(b[34]), .Z(n43667) );
  XOR U44778 ( .A(n43673), .B(n43674), .Z(n43456) );
  ANDN U44779 ( .B(n43675), .A(n43676), .Z(n43673) );
  AND U44780 ( .A(a[4]), .B(b[33]), .Z(n43672) );
  XOR U44781 ( .A(n43678), .B(n43679), .Z(n43461) );
  ANDN U44782 ( .B(n43680), .A(n43681), .Z(n43678) );
  AND U44783 ( .A(a[5]), .B(b[32]), .Z(n43677) );
  XOR U44784 ( .A(n43683), .B(n43684), .Z(n43466) );
  ANDN U44785 ( .B(n43685), .A(n43686), .Z(n43683) );
  AND U44786 ( .A(a[6]), .B(b[31]), .Z(n43682) );
  XOR U44787 ( .A(n43688), .B(n43689), .Z(n43471) );
  ANDN U44788 ( .B(n43690), .A(n43691), .Z(n43688) );
  AND U44789 ( .A(a[7]), .B(b[30]), .Z(n43687) );
  XOR U44790 ( .A(n43693), .B(n43694), .Z(n43476) );
  ANDN U44791 ( .B(n43695), .A(n43696), .Z(n43693) );
  AND U44792 ( .A(a[8]), .B(b[29]), .Z(n43692) );
  XOR U44793 ( .A(n43698), .B(n43699), .Z(n43481) );
  ANDN U44794 ( .B(n43700), .A(n43701), .Z(n43698) );
  AND U44795 ( .A(a[9]), .B(b[28]), .Z(n43697) );
  XOR U44796 ( .A(n43703), .B(n43704), .Z(n43486) );
  ANDN U44797 ( .B(n43705), .A(n43706), .Z(n43703) );
  AND U44798 ( .A(a[10]), .B(b[27]), .Z(n43702) );
  XOR U44799 ( .A(n43708), .B(n43709), .Z(n43491) );
  ANDN U44800 ( .B(n43710), .A(n43711), .Z(n43708) );
  AND U44801 ( .A(a[11]), .B(b[26]), .Z(n43707) );
  XOR U44802 ( .A(n43713), .B(n43714), .Z(n43496) );
  ANDN U44803 ( .B(n43715), .A(n43716), .Z(n43713) );
  AND U44804 ( .A(a[12]), .B(b[25]), .Z(n43712) );
  XOR U44805 ( .A(n43718), .B(n43719), .Z(n43501) );
  ANDN U44806 ( .B(n43720), .A(n43721), .Z(n43718) );
  AND U44807 ( .A(a[13]), .B(b[24]), .Z(n43717) );
  XOR U44808 ( .A(n43723), .B(n43724), .Z(n43506) );
  ANDN U44809 ( .B(n43725), .A(n43726), .Z(n43723) );
  AND U44810 ( .A(a[14]), .B(b[23]), .Z(n43722) );
  XOR U44811 ( .A(n43728), .B(n43729), .Z(n43511) );
  ANDN U44812 ( .B(n43730), .A(n43731), .Z(n43728) );
  AND U44813 ( .A(a[15]), .B(b[22]), .Z(n43727) );
  XOR U44814 ( .A(n43733), .B(n43734), .Z(n43516) );
  ANDN U44815 ( .B(n43735), .A(n43736), .Z(n43733) );
  AND U44816 ( .A(a[16]), .B(b[21]), .Z(n43732) );
  XOR U44817 ( .A(n43738), .B(n43739), .Z(n43521) );
  ANDN U44818 ( .B(n43740), .A(n43741), .Z(n43738) );
  AND U44819 ( .A(a[17]), .B(b[20]), .Z(n43737) );
  XOR U44820 ( .A(n43743), .B(n43744), .Z(n43526) );
  ANDN U44821 ( .B(n43745), .A(n43746), .Z(n43743) );
  AND U44822 ( .A(a[18]), .B(b[19]), .Z(n43742) );
  XOR U44823 ( .A(n43748), .B(n43749), .Z(n43531) );
  ANDN U44824 ( .B(n43750), .A(n43751), .Z(n43748) );
  AND U44825 ( .A(a[19]), .B(b[18]), .Z(n43747) );
  XOR U44826 ( .A(n43753), .B(n43754), .Z(n43536) );
  ANDN U44827 ( .B(n43755), .A(n43756), .Z(n43753) );
  AND U44828 ( .A(a[20]), .B(b[17]), .Z(n43752) );
  XOR U44829 ( .A(n43758), .B(n43759), .Z(n43541) );
  ANDN U44830 ( .B(n43760), .A(n43761), .Z(n43758) );
  AND U44831 ( .A(a[21]), .B(b[16]), .Z(n43757) );
  XOR U44832 ( .A(n43763), .B(n43764), .Z(n43546) );
  ANDN U44833 ( .B(n43765), .A(n43766), .Z(n43763) );
  AND U44834 ( .A(a[22]), .B(b[15]), .Z(n43762) );
  XOR U44835 ( .A(n43768), .B(n43769), .Z(n43551) );
  ANDN U44836 ( .B(n43770), .A(n43771), .Z(n43768) );
  AND U44837 ( .A(a[23]), .B(b[14]), .Z(n43767) );
  XOR U44838 ( .A(n43773), .B(n43774), .Z(n43556) );
  ANDN U44839 ( .B(n43775), .A(n43776), .Z(n43773) );
  AND U44840 ( .A(a[24]), .B(b[13]), .Z(n43772) );
  XOR U44841 ( .A(n43778), .B(n43779), .Z(n43561) );
  ANDN U44842 ( .B(n43780), .A(n43781), .Z(n43778) );
  AND U44843 ( .A(a[25]), .B(b[12]), .Z(n43777) );
  XOR U44844 ( .A(n43783), .B(n43784), .Z(n43566) );
  ANDN U44845 ( .B(n43785), .A(n43786), .Z(n43783) );
  AND U44846 ( .A(a[26]), .B(b[11]), .Z(n43782) );
  XOR U44847 ( .A(n43788), .B(n43789), .Z(n43571) );
  ANDN U44848 ( .B(n43790), .A(n43791), .Z(n43788) );
  AND U44849 ( .A(a[27]), .B(b[10]), .Z(n43787) );
  XOR U44850 ( .A(n43793), .B(n43794), .Z(n43576) );
  ANDN U44851 ( .B(n43795), .A(n43796), .Z(n43793) );
  AND U44852 ( .A(b[9]), .B(a[28]), .Z(n43792) );
  XOR U44853 ( .A(n43798), .B(n43799), .Z(n43581) );
  ANDN U44854 ( .B(n43800), .A(n43801), .Z(n43798) );
  AND U44855 ( .A(b[8]), .B(a[29]), .Z(n43797) );
  XOR U44856 ( .A(n43803), .B(n43804), .Z(n43586) );
  ANDN U44857 ( .B(n43805), .A(n43806), .Z(n43803) );
  AND U44858 ( .A(b[7]), .B(a[30]), .Z(n43802) );
  XOR U44859 ( .A(n43808), .B(n43809), .Z(n43591) );
  ANDN U44860 ( .B(n43810), .A(n43811), .Z(n43808) );
  AND U44861 ( .A(b[6]), .B(a[31]), .Z(n43807) );
  XOR U44862 ( .A(n43813), .B(n43814), .Z(n43596) );
  ANDN U44863 ( .B(n43815), .A(n43816), .Z(n43813) );
  AND U44864 ( .A(b[5]), .B(a[32]), .Z(n43812) );
  XOR U44865 ( .A(n43818), .B(n43819), .Z(n43601) );
  ANDN U44866 ( .B(n43820), .A(n43821), .Z(n43818) );
  AND U44867 ( .A(b[4]), .B(a[33]), .Z(n43817) );
  XOR U44868 ( .A(n43823), .B(n43824), .Z(n43606) );
  ANDN U44869 ( .B(n43618), .A(n43619), .Z(n43823) );
  AND U44870 ( .A(b[2]), .B(a[34]), .Z(n43825) );
  XNOR U44871 ( .A(n43820), .B(n43824), .Z(n43826) );
  XOR U44872 ( .A(n43827), .B(n43828), .Z(n43824) );
  OR U44873 ( .A(n43621), .B(n43622), .Z(n43828) );
  XNOR U44874 ( .A(n43830), .B(n43831), .Z(n43829) );
  XOR U44875 ( .A(n43830), .B(n43833), .Z(n43621) );
  NAND U44876 ( .A(b[1]), .B(a[34]), .Z(n43833) );
  IV U44877 ( .A(n43827), .Z(n43830) );
  NANDN U44878 ( .A(n145), .B(n146), .Z(n43827) );
  XOR U44879 ( .A(n43834), .B(n43835), .Z(n146) );
  NAND U44880 ( .A(a[34]), .B(b[0]), .Z(n145) );
  XNOR U44881 ( .A(n43815), .B(n43819), .Z(n43836) );
  XNOR U44882 ( .A(n43810), .B(n43814), .Z(n43837) );
  XNOR U44883 ( .A(n43805), .B(n43809), .Z(n43838) );
  XNOR U44884 ( .A(n43800), .B(n43804), .Z(n43839) );
  XNOR U44885 ( .A(n43795), .B(n43799), .Z(n43840) );
  XNOR U44886 ( .A(n43790), .B(n43794), .Z(n43841) );
  XNOR U44887 ( .A(n43785), .B(n43789), .Z(n43842) );
  XNOR U44888 ( .A(n43780), .B(n43784), .Z(n43843) );
  XNOR U44889 ( .A(n43775), .B(n43779), .Z(n43844) );
  XNOR U44890 ( .A(n43770), .B(n43774), .Z(n43845) );
  XNOR U44891 ( .A(n43765), .B(n43769), .Z(n43846) );
  XNOR U44892 ( .A(n43760), .B(n43764), .Z(n43847) );
  XNOR U44893 ( .A(n43755), .B(n43759), .Z(n43848) );
  XNOR U44894 ( .A(n43750), .B(n43754), .Z(n43849) );
  XNOR U44895 ( .A(n43745), .B(n43749), .Z(n43850) );
  XNOR U44896 ( .A(n43740), .B(n43744), .Z(n43851) );
  XNOR U44897 ( .A(n43735), .B(n43739), .Z(n43852) );
  XNOR U44898 ( .A(n43730), .B(n43734), .Z(n43853) );
  XNOR U44899 ( .A(n43725), .B(n43729), .Z(n43854) );
  XNOR U44900 ( .A(n43720), .B(n43724), .Z(n43855) );
  XNOR U44901 ( .A(n43715), .B(n43719), .Z(n43856) );
  XNOR U44902 ( .A(n43710), .B(n43714), .Z(n43857) );
  XNOR U44903 ( .A(n43705), .B(n43709), .Z(n43858) );
  XNOR U44904 ( .A(n43700), .B(n43704), .Z(n43859) );
  XNOR U44905 ( .A(n43695), .B(n43699), .Z(n43860) );
  XNOR U44906 ( .A(n43690), .B(n43694), .Z(n43861) );
  XNOR U44907 ( .A(n43685), .B(n43689), .Z(n43862) );
  XNOR U44908 ( .A(n43680), .B(n43684), .Z(n43863) );
  XNOR U44909 ( .A(n43675), .B(n43679), .Z(n43864) );
  XNOR U44910 ( .A(n43670), .B(n43674), .Z(n43865) );
  XNOR U44911 ( .A(n43665), .B(n43669), .Z(n43866) );
  XNOR U44912 ( .A(n43660), .B(n43664), .Z(n43867) );
  XOR U44913 ( .A(n43868), .B(n43659), .Z(n43660) );
  AND U44914 ( .A(a[0]), .B(b[36]), .Z(n43868) );
  XNOR U44915 ( .A(n43869), .B(n43659), .Z(n43661) );
  XNOR U44916 ( .A(n43870), .B(n43871), .Z(n43659) );
  ANDN U44917 ( .B(n43872), .A(n43873), .Z(n43870) );
  AND U44918 ( .A(a[1]), .B(b[35]), .Z(n43869) );
  XOR U44919 ( .A(n43875), .B(n43876), .Z(n43664) );
  ANDN U44920 ( .B(n43877), .A(n43878), .Z(n43875) );
  AND U44921 ( .A(a[2]), .B(b[34]), .Z(n43874) );
  XOR U44922 ( .A(n43880), .B(n43881), .Z(n43669) );
  ANDN U44923 ( .B(n43882), .A(n43883), .Z(n43880) );
  AND U44924 ( .A(a[3]), .B(b[33]), .Z(n43879) );
  XOR U44925 ( .A(n43885), .B(n43886), .Z(n43674) );
  ANDN U44926 ( .B(n43887), .A(n43888), .Z(n43885) );
  AND U44927 ( .A(a[4]), .B(b[32]), .Z(n43884) );
  XOR U44928 ( .A(n43890), .B(n43891), .Z(n43679) );
  ANDN U44929 ( .B(n43892), .A(n43893), .Z(n43890) );
  AND U44930 ( .A(a[5]), .B(b[31]), .Z(n43889) );
  XOR U44931 ( .A(n43895), .B(n43896), .Z(n43684) );
  ANDN U44932 ( .B(n43897), .A(n43898), .Z(n43895) );
  AND U44933 ( .A(a[6]), .B(b[30]), .Z(n43894) );
  XOR U44934 ( .A(n43900), .B(n43901), .Z(n43689) );
  ANDN U44935 ( .B(n43902), .A(n43903), .Z(n43900) );
  AND U44936 ( .A(a[7]), .B(b[29]), .Z(n43899) );
  XOR U44937 ( .A(n43905), .B(n43906), .Z(n43694) );
  ANDN U44938 ( .B(n43907), .A(n43908), .Z(n43905) );
  AND U44939 ( .A(a[8]), .B(b[28]), .Z(n43904) );
  XOR U44940 ( .A(n43910), .B(n43911), .Z(n43699) );
  ANDN U44941 ( .B(n43912), .A(n43913), .Z(n43910) );
  AND U44942 ( .A(a[9]), .B(b[27]), .Z(n43909) );
  XOR U44943 ( .A(n43915), .B(n43916), .Z(n43704) );
  ANDN U44944 ( .B(n43917), .A(n43918), .Z(n43915) );
  AND U44945 ( .A(a[10]), .B(b[26]), .Z(n43914) );
  XOR U44946 ( .A(n43920), .B(n43921), .Z(n43709) );
  ANDN U44947 ( .B(n43922), .A(n43923), .Z(n43920) );
  AND U44948 ( .A(a[11]), .B(b[25]), .Z(n43919) );
  XOR U44949 ( .A(n43925), .B(n43926), .Z(n43714) );
  ANDN U44950 ( .B(n43927), .A(n43928), .Z(n43925) );
  AND U44951 ( .A(a[12]), .B(b[24]), .Z(n43924) );
  XOR U44952 ( .A(n43930), .B(n43931), .Z(n43719) );
  ANDN U44953 ( .B(n43932), .A(n43933), .Z(n43930) );
  AND U44954 ( .A(a[13]), .B(b[23]), .Z(n43929) );
  XOR U44955 ( .A(n43935), .B(n43936), .Z(n43724) );
  ANDN U44956 ( .B(n43937), .A(n43938), .Z(n43935) );
  AND U44957 ( .A(a[14]), .B(b[22]), .Z(n43934) );
  XOR U44958 ( .A(n43940), .B(n43941), .Z(n43729) );
  ANDN U44959 ( .B(n43942), .A(n43943), .Z(n43940) );
  AND U44960 ( .A(a[15]), .B(b[21]), .Z(n43939) );
  XOR U44961 ( .A(n43945), .B(n43946), .Z(n43734) );
  ANDN U44962 ( .B(n43947), .A(n43948), .Z(n43945) );
  AND U44963 ( .A(a[16]), .B(b[20]), .Z(n43944) );
  XOR U44964 ( .A(n43950), .B(n43951), .Z(n43739) );
  ANDN U44965 ( .B(n43952), .A(n43953), .Z(n43950) );
  AND U44966 ( .A(a[17]), .B(b[19]), .Z(n43949) );
  XOR U44967 ( .A(n43955), .B(n43956), .Z(n43744) );
  ANDN U44968 ( .B(n43957), .A(n43958), .Z(n43955) );
  AND U44969 ( .A(a[18]), .B(b[18]), .Z(n43954) );
  XOR U44970 ( .A(n43960), .B(n43961), .Z(n43749) );
  ANDN U44971 ( .B(n43962), .A(n43963), .Z(n43960) );
  AND U44972 ( .A(a[19]), .B(b[17]), .Z(n43959) );
  XOR U44973 ( .A(n43965), .B(n43966), .Z(n43754) );
  ANDN U44974 ( .B(n43967), .A(n43968), .Z(n43965) );
  AND U44975 ( .A(a[20]), .B(b[16]), .Z(n43964) );
  XOR U44976 ( .A(n43970), .B(n43971), .Z(n43759) );
  ANDN U44977 ( .B(n43972), .A(n43973), .Z(n43970) );
  AND U44978 ( .A(a[21]), .B(b[15]), .Z(n43969) );
  XOR U44979 ( .A(n43975), .B(n43976), .Z(n43764) );
  ANDN U44980 ( .B(n43977), .A(n43978), .Z(n43975) );
  AND U44981 ( .A(a[22]), .B(b[14]), .Z(n43974) );
  XOR U44982 ( .A(n43980), .B(n43981), .Z(n43769) );
  ANDN U44983 ( .B(n43982), .A(n43983), .Z(n43980) );
  AND U44984 ( .A(a[23]), .B(b[13]), .Z(n43979) );
  XOR U44985 ( .A(n43985), .B(n43986), .Z(n43774) );
  ANDN U44986 ( .B(n43987), .A(n43988), .Z(n43985) );
  AND U44987 ( .A(a[24]), .B(b[12]), .Z(n43984) );
  XOR U44988 ( .A(n43990), .B(n43991), .Z(n43779) );
  ANDN U44989 ( .B(n43992), .A(n43993), .Z(n43990) );
  AND U44990 ( .A(a[25]), .B(b[11]), .Z(n43989) );
  XOR U44991 ( .A(n43995), .B(n43996), .Z(n43784) );
  ANDN U44992 ( .B(n43997), .A(n43998), .Z(n43995) );
  AND U44993 ( .A(a[26]), .B(b[10]), .Z(n43994) );
  XOR U44994 ( .A(n44000), .B(n44001), .Z(n43789) );
  ANDN U44995 ( .B(n44002), .A(n44003), .Z(n44000) );
  AND U44996 ( .A(b[9]), .B(a[27]), .Z(n43999) );
  XOR U44997 ( .A(n44005), .B(n44006), .Z(n43794) );
  ANDN U44998 ( .B(n44007), .A(n44008), .Z(n44005) );
  AND U44999 ( .A(b[8]), .B(a[28]), .Z(n44004) );
  XOR U45000 ( .A(n44010), .B(n44011), .Z(n43799) );
  ANDN U45001 ( .B(n44012), .A(n44013), .Z(n44010) );
  AND U45002 ( .A(b[7]), .B(a[29]), .Z(n44009) );
  XOR U45003 ( .A(n44015), .B(n44016), .Z(n43804) );
  ANDN U45004 ( .B(n44017), .A(n44018), .Z(n44015) );
  AND U45005 ( .A(b[6]), .B(a[30]), .Z(n44014) );
  XOR U45006 ( .A(n44020), .B(n44021), .Z(n43809) );
  ANDN U45007 ( .B(n44022), .A(n44023), .Z(n44020) );
  AND U45008 ( .A(b[5]), .B(a[31]), .Z(n44019) );
  XOR U45009 ( .A(n44025), .B(n44026), .Z(n43814) );
  ANDN U45010 ( .B(n44027), .A(n44028), .Z(n44025) );
  AND U45011 ( .A(b[4]), .B(a[32]), .Z(n44024) );
  XOR U45012 ( .A(n44030), .B(n44031), .Z(n43819) );
  ANDN U45013 ( .B(n43831), .A(n43832), .Z(n44030) );
  AND U45014 ( .A(b[2]), .B(a[33]), .Z(n44032) );
  XNOR U45015 ( .A(n44027), .B(n44031), .Z(n44033) );
  XOR U45016 ( .A(n44034), .B(n44035), .Z(n44031) );
  OR U45017 ( .A(n43834), .B(n43835), .Z(n44035) );
  XNOR U45018 ( .A(n44037), .B(n44038), .Z(n44036) );
  XOR U45019 ( .A(n44037), .B(n44040), .Z(n43834) );
  NAND U45020 ( .A(b[1]), .B(a[33]), .Z(n44040) );
  IV U45021 ( .A(n44034), .Z(n44037) );
  NANDN U45022 ( .A(n147), .B(n148), .Z(n44034) );
  XOR U45023 ( .A(n44041), .B(n44042), .Z(n148) );
  NAND U45024 ( .A(a[33]), .B(b[0]), .Z(n147) );
  XNOR U45025 ( .A(n44022), .B(n44026), .Z(n44043) );
  XNOR U45026 ( .A(n44017), .B(n44021), .Z(n44044) );
  XNOR U45027 ( .A(n44012), .B(n44016), .Z(n44045) );
  XNOR U45028 ( .A(n44007), .B(n44011), .Z(n44046) );
  XNOR U45029 ( .A(n44002), .B(n44006), .Z(n44047) );
  XNOR U45030 ( .A(n43997), .B(n44001), .Z(n44048) );
  XNOR U45031 ( .A(n43992), .B(n43996), .Z(n44049) );
  XNOR U45032 ( .A(n43987), .B(n43991), .Z(n44050) );
  XNOR U45033 ( .A(n43982), .B(n43986), .Z(n44051) );
  XNOR U45034 ( .A(n43977), .B(n43981), .Z(n44052) );
  XNOR U45035 ( .A(n43972), .B(n43976), .Z(n44053) );
  XNOR U45036 ( .A(n43967), .B(n43971), .Z(n44054) );
  XNOR U45037 ( .A(n43962), .B(n43966), .Z(n44055) );
  XNOR U45038 ( .A(n43957), .B(n43961), .Z(n44056) );
  XNOR U45039 ( .A(n43952), .B(n43956), .Z(n44057) );
  XNOR U45040 ( .A(n43947), .B(n43951), .Z(n44058) );
  XNOR U45041 ( .A(n43942), .B(n43946), .Z(n44059) );
  XNOR U45042 ( .A(n43937), .B(n43941), .Z(n44060) );
  XNOR U45043 ( .A(n43932), .B(n43936), .Z(n44061) );
  XNOR U45044 ( .A(n43927), .B(n43931), .Z(n44062) );
  XNOR U45045 ( .A(n43922), .B(n43926), .Z(n44063) );
  XNOR U45046 ( .A(n43917), .B(n43921), .Z(n44064) );
  XNOR U45047 ( .A(n43912), .B(n43916), .Z(n44065) );
  XNOR U45048 ( .A(n43907), .B(n43911), .Z(n44066) );
  XNOR U45049 ( .A(n43902), .B(n43906), .Z(n44067) );
  XNOR U45050 ( .A(n43897), .B(n43901), .Z(n44068) );
  XNOR U45051 ( .A(n43892), .B(n43896), .Z(n44069) );
  XNOR U45052 ( .A(n43887), .B(n43891), .Z(n44070) );
  XNOR U45053 ( .A(n43882), .B(n43886), .Z(n44071) );
  XNOR U45054 ( .A(n43877), .B(n43881), .Z(n44072) );
  XNOR U45055 ( .A(n43872), .B(n43876), .Z(n44073) );
  XNOR U45056 ( .A(n44074), .B(n43871), .Z(n43872) );
  AND U45057 ( .A(a[0]), .B(b[35]), .Z(n44074) );
  XOR U45058 ( .A(n44075), .B(n43871), .Z(n43873) );
  XNOR U45059 ( .A(n44076), .B(n44077), .Z(n43871) );
  ANDN U45060 ( .B(n44078), .A(n44079), .Z(n44076) );
  AND U45061 ( .A(a[1]), .B(b[34]), .Z(n44075) );
  XOR U45062 ( .A(n44081), .B(n44082), .Z(n43876) );
  ANDN U45063 ( .B(n44083), .A(n44084), .Z(n44081) );
  AND U45064 ( .A(a[2]), .B(b[33]), .Z(n44080) );
  XOR U45065 ( .A(n44086), .B(n44087), .Z(n43881) );
  ANDN U45066 ( .B(n44088), .A(n44089), .Z(n44086) );
  AND U45067 ( .A(a[3]), .B(b[32]), .Z(n44085) );
  XOR U45068 ( .A(n44091), .B(n44092), .Z(n43886) );
  ANDN U45069 ( .B(n44093), .A(n44094), .Z(n44091) );
  AND U45070 ( .A(a[4]), .B(b[31]), .Z(n44090) );
  XOR U45071 ( .A(n44096), .B(n44097), .Z(n43891) );
  ANDN U45072 ( .B(n44098), .A(n44099), .Z(n44096) );
  AND U45073 ( .A(a[5]), .B(b[30]), .Z(n44095) );
  XOR U45074 ( .A(n44101), .B(n44102), .Z(n43896) );
  ANDN U45075 ( .B(n44103), .A(n44104), .Z(n44101) );
  AND U45076 ( .A(a[6]), .B(b[29]), .Z(n44100) );
  XOR U45077 ( .A(n44106), .B(n44107), .Z(n43901) );
  ANDN U45078 ( .B(n44108), .A(n44109), .Z(n44106) );
  AND U45079 ( .A(a[7]), .B(b[28]), .Z(n44105) );
  XOR U45080 ( .A(n44111), .B(n44112), .Z(n43906) );
  ANDN U45081 ( .B(n44113), .A(n44114), .Z(n44111) );
  AND U45082 ( .A(a[8]), .B(b[27]), .Z(n44110) );
  XOR U45083 ( .A(n44116), .B(n44117), .Z(n43911) );
  ANDN U45084 ( .B(n44118), .A(n44119), .Z(n44116) );
  AND U45085 ( .A(a[9]), .B(b[26]), .Z(n44115) );
  XOR U45086 ( .A(n44121), .B(n44122), .Z(n43916) );
  ANDN U45087 ( .B(n44123), .A(n44124), .Z(n44121) );
  AND U45088 ( .A(a[10]), .B(b[25]), .Z(n44120) );
  XOR U45089 ( .A(n44126), .B(n44127), .Z(n43921) );
  ANDN U45090 ( .B(n44128), .A(n44129), .Z(n44126) );
  AND U45091 ( .A(a[11]), .B(b[24]), .Z(n44125) );
  XOR U45092 ( .A(n44131), .B(n44132), .Z(n43926) );
  ANDN U45093 ( .B(n44133), .A(n44134), .Z(n44131) );
  AND U45094 ( .A(a[12]), .B(b[23]), .Z(n44130) );
  XOR U45095 ( .A(n44136), .B(n44137), .Z(n43931) );
  ANDN U45096 ( .B(n44138), .A(n44139), .Z(n44136) );
  AND U45097 ( .A(a[13]), .B(b[22]), .Z(n44135) );
  XOR U45098 ( .A(n44141), .B(n44142), .Z(n43936) );
  ANDN U45099 ( .B(n44143), .A(n44144), .Z(n44141) );
  AND U45100 ( .A(a[14]), .B(b[21]), .Z(n44140) );
  XOR U45101 ( .A(n44146), .B(n44147), .Z(n43941) );
  ANDN U45102 ( .B(n44148), .A(n44149), .Z(n44146) );
  AND U45103 ( .A(a[15]), .B(b[20]), .Z(n44145) );
  XOR U45104 ( .A(n44151), .B(n44152), .Z(n43946) );
  ANDN U45105 ( .B(n44153), .A(n44154), .Z(n44151) );
  AND U45106 ( .A(a[16]), .B(b[19]), .Z(n44150) );
  XOR U45107 ( .A(n44156), .B(n44157), .Z(n43951) );
  ANDN U45108 ( .B(n44158), .A(n44159), .Z(n44156) );
  AND U45109 ( .A(a[17]), .B(b[18]), .Z(n44155) );
  XOR U45110 ( .A(n44161), .B(n44162), .Z(n43956) );
  ANDN U45111 ( .B(n44163), .A(n44164), .Z(n44161) );
  AND U45112 ( .A(a[18]), .B(b[17]), .Z(n44160) );
  XOR U45113 ( .A(n44166), .B(n44167), .Z(n43961) );
  ANDN U45114 ( .B(n44168), .A(n44169), .Z(n44166) );
  AND U45115 ( .A(a[19]), .B(b[16]), .Z(n44165) );
  XOR U45116 ( .A(n44171), .B(n44172), .Z(n43966) );
  ANDN U45117 ( .B(n44173), .A(n44174), .Z(n44171) );
  AND U45118 ( .A(a[20]), .B(b[15]), .Z(n44170) );
  XOR U45119 ( .A(n44176), .B(n44177), .Z(n43971) );
  ANDN U45120 ( .B(n44178), .A(n44179), .Z(n44176) );
  AND U45121 ( .A(a[21]), .B(b[14]), .Z(n44175) );
  XOR U45122 ( .A(n44181), .B(n44182), .Z(n43976) );
  ANDN U45123 ( .B(n44183), .A(n44184), .Z(n44181) );
  AND U45124 ( .A(a[22]), .B(b[13]), .Z(n44180) );
  XOR U45125 ( .A(n44186), .B(n44187), .Z(n43981) );
  ANDN U45126 ( .B(n44188), .A(n44189), .Z(n44186) );
  AND U45127 ( .A(a[23]), .B(b[12]), .Z(n44185) );
  XOR U45128 ( .A(n44191), .B(n44192), .Z(n43986) );
  ANDN U45129 ( .B(n44193), .A(n44194), .Z(n44191) );
  AND U45130 ( .A(a[24]), .B(b[11]), .Z(n44190) );
  XOR U45131 ( .A(n44196), .B(n44197), .Z(n43991) );
  ANDN U45132 ( .B(n44198), .A(n44199), .Z(n44196) );
  AND U45133 ( .A(a[25]), .B(b[10]), .Z(n44195) );
  XOR U45134 ( .A(n44201), .B(n44202), .Z(n43996) );
  ANDN U45135 ( .B(n44203), .A(n44204), .Z(n44201) );
  AND U45136 ( .A(b[9]), .B(a[26]), .Z(n44200) );
  XOR U45137 ( .A(n44206), .B(n44207), .Z(n44001) );
  ANDN U45138 ( .B(n44208), .A(n44209), .Z(n44206) );
  AND U45139 ( .A(b[8]), .B(a[27]), .Z(n44205) );
  XOR U45140 ( .A(n44211), .B(n44212), .Z(n44006) );
  ANDN U45141 ( .B(n44213), .A(n44214), .Z(n44211) );
  AND U45142 ( .A(b[7]), .B(a[28]), .Z(n44210) );
  XOR U45143 ( .A(n44216), .B(n44217), .Z(n44011) );
  ANDN U45144 ( .B(n44218), .A(n44219), .Z(n44216) );
  AND U45145 ( .A(b[6]), .B(a[29]), .Z(n44215) );
  XOR U45146 ( .A(n44221), .B(n44222), .Z(n44016) );
  ANDN U45147 ( .B(n44223), .A(n44224), .Z(n44221) );
  AND U45148 ( .A(b[5]), .B(a[30]), .Z(n44220) );
  XOR U45149 ( .A(n44226), .B(n44227), .Z(n44021) );
  ANDN U45150 ( .B(n44228), .A(n44229), .Z(n44226) );
  AND U45151 ( .A(b[4]), .B(a[31]), .Z(n44225) );
  XOR U45152 ( .A(n44231), .B(n44232), .Z(n44026) );
  ANDN U45153 ( .B(n44038), .A(n44039), .Z(n44231) );
  AND U45154 ( .A(b[2]), .B(a[32]), .Z(n44233) );
  XNOR U45155 ( .A(n44228), .B(n44232), .Z(n44234) );
  XOR U45156 ( .A(n44235), .B(n44236), .Z(n44232) );
  OR U45157 ( .A(n44041), .B(n44042), .Z(n44236) );
  XNOR U45158 ( .A(n44238), .B(n44239), .Z(n44237) );
  XOR U45159 ( .A(n44238), .B(n44241), .Z(n44041) );
  NAND U45160 ( .A(b[1]), .B(a[32]), .Z(n44241) );
  IV U45161 ( .A(n44235), .Z(n44238) );
  NANDN U45162 ( .A(n149), .B(n150), .Z(n44235) );
  XOR U45163 ( .A(n44242), .B(n44243), .Z(n150) );
  NAND U45164 ( .A(a[32]), .B(b[0]), .Z(n149) );
  XNOR U45165 ( .A(n44223), .B(n44227), .Z(n44244) );
  XNOR U45166 ( .A(n44218), .B(n44222), .Z(n44245) );
  XNOR U45167 ( .A(n44213), .B(n44217), .Z(n44246) );
  XNOR U45168 ( .A(n44208), .B(n44212), .Z(n44247) );
  XNOR U45169 ( .A(n44203), .B(n44207), .Z(n44248) );
  XNOR U45170 ( .A(n44198), .B(n44202), .Z(n44249) );
  XNOR U45171 ( .A(n44193), .B(n44197), .Z(n44250) );
  XNOR U45172 ( .A(n44188), .B(n44192), .Z(n44251) );
  XNOR U45173 ( .A(n44183), .B(n44187), .Z(n44252) );
  XNOR U45174 ( .A(n44178), .B(n44182), .Z(n44253) );
  XNOR U45175 ( .A(n44173), .B(n44177), .Z(n44254) );
  XNOR U45176 ( .A(n44168), .B(n44172), .Z(n44255) );
  XNOR U45177 ( .A(n44163), .B(n44167), .Z(n44256) );
  XNOR U45178 ( .A(n44158), .B(n44162), .Z(n44257) );
  XNOR U45179 ( .A(n44153), .B(n44157), .Z(n44258) );
  XNOR U45180 ( .A(n44148), .B(n44152), .Z(n44259) );
  XNOR U45181 ( .A(n44143), .B(n44147), .Z(n44260) );
  XNOR U45182 ( .A(n44138), .B(n44142), .Z(n44261) );
  XNOR U45183 ( .A(n44133), .B(n44137), .Z(n44262) );
  XNOR U45184 ( .A(n44128), .B(n44132), .Z(n44263) );
  XNOR U45185 ( .A(n44123), .B(n44127), .Z(n44264) );
  XNOR U45186 ( .A(n44118), .B(n44122), .Z(n44265) );
  XNOR U45187 ( .A(n44113), .B(n44117), .Z(n44266) );
  XNOR U45188 ( .A(n44108), .B(n44112), .Z(n44267) );
  XNOR U45189 ( .A(n44103), .B(n44107), .Z(n44268) );
  XNOR U45190 ( .A(n44098), .B(n44102), .Z(n44269) );
  XNOR U45191 ( .A(n44093), .B(n44097), .Z(n44270) );
  XNOR U45192 ( .A(n44088), .B(n44092), .Z(n44271) );
  XNOR U45193 ( .A(n44083), .B(n44087), .Z(n44272) );
  XNOR U45194 ( .A(n44078), .B(n44082), .Z(n44273) );
  XOR U45195 ( .A(n44274), .B(n44077), .Z(n44078) );
  AND U45196 ( .A(a[0]), .B(b[34]), .Z(n44274) );
  XNOR U45197 ( .A(n44275), .B(n44077), .Z(n44079) );
  XNOR U45198 ( .A(n44276), .B(n44277), .Z(n44077) );
  ANDN U45199 ( .B(n44278), .A(n44279), .Z(n44276) );
  AND U45200 ( .A(a[1]), .B(b[33]), .Z(n44275) );
  XOR U45201 ( .A(n44281), .B(n44282), .Z(n44082) );
  ANDN U45202 ( .B(n44283), .A(n44284), .Z(n44281) );
  AND U45203 ( .A(a[2]), .B(b[32]), .Z(n44280) );
  XOR U45204 ( .A(n44286), .B(n44287), .Z(n44087) );
  ANDN U45205 ( .B(n44288), .A(n44289), .Z(n44286) );
  AND U45206 ( .A(a[3]), .B(b[31]), .Z(n44285) );
  XOR U45207 ( .A(n44291), .B(n44292), .Z(n44092) );
  ANDN U45208 ( .B(n44293), .A(n44294), .Z(n44291) );
  AND U45209 ( .A(a[4]), .B(b[30]), .Z(n44290) );
  XOR U45210 ( .A(n44296), .B(n44297), .Z(n44097) );
  ANDN U45211 ( .B(n44298), .A(n44299), .Z(n44296) );
  AND U45212 ( .A(a[5]), .B(b[29]), .Z(n44295) );
  XOR U45213 ( .A(n44301), .B(n44302), .Z(n44102) );
  ANDN U45214 ( .B(n44303), .A(n44304), .Z(n44301) );
  AND U45215 ( .A(a[6]), .B(b[28]), .Z(n44300) );
  XOR U45216 ( .A(n44306), .B(n44307), .Z(n44107) );
  ANDN U45217 ( .B(n44308), .A(n44309), .Z(n44306) );
  AND U45218 ( .A(a[7]), .B(b[27]), .Z(n44305) );
  XOR U45219 ( .A(n44311), .B(n44312), .Z(n44112) );
  ANDN U45220 ( .B(n44313), .A(n44314), .Z(n44311) );
  AND U45221 ( .A(a[8]), .B(b[26]), .Z(n44310) );
  XOR U45222 ( .A(n44316), .B(n44317), .Z(n44117) );
  ANDN U45223 ( .B(n44318), .A(n44319), .Z(n44316) );
  AND U45224 ( .A(a[9]), .B(b[25]), .Z(n44315) );
  XOR U45225 ( .A(n44321), .B(n44322), .Z(n44122) );
  ANDN U45226 ( .B(n44323), .A(n44324), .Z(n44321) );
  AND U45227 ( .A(a[10]), .B(b[24]), .Z(n44320) );
  XOR U45228 ( .A(n44326), .B(n44327), .Z(n44127) );
  ANDN U45229 ( .B(n44328), .A(n44329), .Z(n44326) );
  AND U45230 ( .A(a[11]), .B(b[23]), .Z(n44325) );
  XOR U45231 ( .A(n44331), .B(n44332), .Z(n44132) );
  ANDN U45232 ( .B(n44333), .A(n44334), .Z(n44331) );
  AND U45233 ( .A(a[12]), .B(b[22]), .Z(n44330) );
  XOR U45234 ( .A(n44336), .B(n44337), .Z(n44137) );
  ANDN U45235 ( .B(n44338), .A(n44339), .Z(n44336) );
  AND U45236 ( .A(a[13]), .B(b[21]), .Z(n44335) );
  XOR U45237 ( .A(n44341), .B(n44342), .Z(n44142) );
  ANDN U45238 ( .B(n44343), .A(n44344), .Z(n44341) );
  AND U45239 ( .A(a[14]), .B(b[20]), .Z(n44340) );
  XOR U45240 ( .A(n44346), .B(n44347), .Z(n44147) );
  ANDN U45241 ( .B(n44348), .A(n44349), .Z(n44346) );
  AND U45242 ( .A(a[15]), .B(b[19]), .Z(n44345) );
  XOR U45243 ( .A(n44351), .B(n44352), .Z(n44152) );
  ANDN U45244 ( .B(n44353), .A(n44354), .Z(n44351) );
  AND U45245 ( .A(a[16]), .B(b[18]), .Z(n44350) );
  XOR U45246 ( .A(n44356), .B(n44357), .Z(n44157) );
  ANDN U45247 ( .B(n44358), .A(n44359), .Z(n44356) );
  AND U45248 ( .A(a[17]), .B(b[17]), .Z(n44355) );
  XOR U45249 ( .A(n44361), .B(n44362), .Z(n44162) );
  ANDN U45250 ( .B(n44363), .A(n44364), .Z(n44361) );
  AND U45251 ( .A(a[18]), .B(b[16]), .Z(n44360) );
  XOR U45252 ( .A(n44366), .B(n44367), .Z(n44167) );
  ANDN U45253 ( .B(n44368), .A(n44369), .Z(n44366) );
  AND U45254 ( .A(a[19]), .B(b[15]), .Z(n44365) );
  XOR U45255 ( .A(n44371), .B(n44372), .Z(n44172) );
  ANDN U45256 ( .B(n44373), .A(n44374), .Z(n44371) );
  AND U45257 ( .A(a[20]), .B(b[14]), .Z(n44370) );
  XOR U45258 ( .A(n44376), .B(n44377), .Z(n44177) );
  ANDN U45259 ( .B(n44378), .A(n44379), .Z(n44376) );
  AND U45260 ( .A(a[21]), .B(b[13]), .Z(n44375) );
  XOR U45261 ( .A(n44381), .B(n44382), .Z(n44182) );
  ANDN U45262 ( .B(n44383), .A(n44384), .Z(n44381) );
  AND U45263 ( .A(a[22]), .B(b[12]), .Z(n44380) );
  XOR U45264 ( .A(n44386), .B(n44387), .Z(n44187) );
  ANDN U45265 ( .B(n44388), .A(n44389), .Z(n44386) );
  AND U45266 ( .A(a[23]), .B(b[11]), .Z(n44385) );
  XOR U45267 ( .A(n44391), .B(n44392), .Z(n44192) );
  ANDN U45268 ( .B(n44393), .A(n44394), .Z(n44391) );
  AND U45269 ( .A(a[24]), .B(b[10]), .Z(n44390) );
  XOR U45270 ( .A(n44396), .B(n44397), .Z(n44197) );
  ANDN U45271 ( .B(n44398), .A(n44399), .Z(n44396) );
  AND U45272 ( .A(b[9]), .B(a[25]), .Z(n44395) );
  XOR U45273 ( .A(n44401), .B(n44402), .Z(n44202) );
  ANDN U45274 ( .B(n44403), .A(n44404), .Z(n44401) );
  AND U45275 ( .A(b[8]), .B(a[26]), .Z(n44400) );
  XOR U45276 ( .A(n44406), .B(n44407), .Z(n44207) );
  ANDN U45277 ( .B(n44408), .A(n44409), .Z(n44406) );
  AND U45278 ( .A(b[7]), .B(a[27]), .Z(n44405) );
  XOR U45279 ( .A(n44411), .B(n44412), .Z(n44212) );
  ANDN U45280 ( .B(n44413), .A(n44414), .Z(n44411) );
  AND U45281 ( .A(b[6]), .B(a[28]), .Z(n44410) );
  XOR U45282 ( .A(n44416), .B(n44417), .Z(n44217) );
  ANDN U45283 ( .B(n44418), .A(n44419), .Z(n44416) );
  AND U45284 ( .A(b[5]), .B(a[29]), .Z(n44415) );
  XOR U45285 ( .A(n44421), .B(n44422), .Z(n44222) );
  ANDN U45286 ( .B(n44423), .A(n44424), .Z(n44421) );
  AND U45287 ( .A(b[4]), .B(a[30]), .Z(n44420) );
  XOR U45288 ( .A(n44426), .B(n44427), .Z(n44227) );
  ANDN U45289 ( .B(n44239), .A(n44240), .Z(n44426) );
  AND U45290 ( .A(b[2]), .B(a[31]), .Z(n44428) );
  XNOR U45291 ( .A(n44423), .B(n44427), .Z(n44429) );
  XOR U45292 ( .A(n44430), .B(n44431), .Z(n44427) );
  OR U45293 ( .A(n44242), .B(n44243), .Z(n44431) );
  XNOR U45294 ( .A(n44433), .B(n44434), .Z(n44432) );
  XOR U45295 ( .A(n44433), .B(n44436), .Z(n44242) );
  NAND U45296 ( .A(b[1]), .B(a[31]), .Z(n44436) );
  IV U45297 ( .A(n44430), .Z(n44433) );
  NANDN U45298 ( .A(n151), .B(n152), .Z(n44430) );
  XOR U45299 ( .A(n44437), .B(n44438), .Z(n152) );
  NAND U45300 ( .A(a[31]), .B(b[0]), .Z(n151) );
  XNOR U45301 ( .A(n44418), .B(n44422), .Z(n44439) );
  XNOR U45302 ( .A(n44413), .B(n44417), .Z(n44440) );
  XNOR U45303 ( .A(n44408), .B(n44412), .Z(n44441) );
  XNOR U45304 ( .A(n44403), .B(n44407), .Z(n44442) );
  XNOR U45305 ( .A(n44398), .B(n44402), .Z(n44443) );
  XNOR U45306 ( .A(n44393), .B(n44397), .Z(n44444) );
  XNOR U45307 ( .A(n44388), .B(n44392), .Z(n44445) );
  XNOR U45308 ( .A(n44383), .B(n44387), .Z(n44446) );
  XNOR U45309 ( .A(n44378), .B(n44382), .Z(n44447) );
  XNOR U45310 ( .A(n44373), .B(n44377), .Z(n44448) );
  XNOR U45311 ( .A(n44368), .B(n44372), .Z(n44449) );
  XNOR U45312 ( .A(n44363), .B(n44367), .Z(n44450) );
  XNOR U45313 ( .A(n44358), .B(n44362), .Z(n44451) );
  XNOR U45314 ( .A(n44353), .B(n44357), .Z(n44452) );
  XNOR U45315 ( .A(n44348), .B(n44352), .Z(n44453) );
  XNOR U45316 ( .A(n44343), .B(n44347), .Z(n44454) );
  XNOR U45317 ( .A(n44338), .B(n44342), .Z(n44455) );
  XNOR U45318 ( .A(n44333), .B(n44337), .Z(n44456) );
  XNOR U45319 ( .A(n44328), .B(n44332), .Z(n44457) );
  XNOR U45320 ( .A(n44323), .B(n44327), .Z(n44458) );
  XNOR U45321 ( .A(n44318), .B(n44322), .Z(n44459) );
  XNOR U45322 ( .A(n44313), .B(n44317), .Z(n44460) );
  XNOR U45323 ( .A(n44308), .B(n44312), .Z(n44461) );
  XNOR U45324 ( .A(n44303), .B(n44307), .Z(n44462) );
  XNOR U45325 ( .A(n44298), .B(n44302), .Z(n44463) );
  XNOR U45326 ( .A(n44293), .B(n44297), .Z(n44464) );
  XNOR U45327 ( .A(n44288), .B(n44292), .Z(n44465) );
  XNOR U45328 ( .A(n44283), .B(n44287), .Z(n44466) );
  XNOR U45329 ( .A(n44278), .B(n44282), .Z(n44467) );
  XNOR U45330 ( .A(n44468), .B(n44277), .Z(n44278) );
  AND U45331 ( .A(a[0]), .B(b[33]), .Z(n44468) );
  XOR U45332 ( .A(n44469), .B(n44277), .Z(n44279) );
  XNOR U45333 ( .A(n44470), .B(n44471), .Z(n44277) );
  ANDN U45334 ( .B(n44472), .A(n44473), .Z(n44470) );
  AND U45335 ( .A(a[1]), .B(b[32]), .Z(n44469) );
  XOR U45336 ( .A(n44475), .B(n44476), .Z(n44282) );
  ANDN U45337 ( .B(n44477), .A(n44478), .Z(n44475) );
  AND U45338 ( .A(a[2]), .B(b[31]), .Z(n44474) );
  XOR U45339 ( .A(n44480), .B(n44481), .Z(n44287) );
  ANDN U45340 ( .B(n44482), .A(n44483), .Z(n44480) );
  AND U45341 ( .A(a[3]), .B(b[30]), .Z(n44479) );
  XOR U45342 ( .A(n44485), .B(n44486), .Z(n44292) );
  ANDN U45343 ( .B(n44487), .A(n44488), .Z(n44485) );
  AND U45344 ( .A(a[4]), .B(b[29]), .Z(n44484) );
  XOR U45345 ( .A(n44490), .B(n44491), .Z(n44297) );
  ANDN U45346 ( .B(n44492), .A(n44493), .Z(n44490) );
  AND U45347 ( .A(a[5]), .B(b[28]), .Z(n44489) );
  XOR U45348 ( .A(n44495), .B(n44496), .Z(n44302) );
  ANDN U45349 ( .B(n44497), .A(n44498), .Z(n44495) );
  AND U45350 ( .A(a[6]), .B(b[27]), .Z(n44494) );
  XOR U45351 ( .A(n44500), .B(n44501), .Z(n44307) );
  ANDN U45352 ( .B(n44502), .A(n44503), .Z(n44500) );
  AND U45353 ( .A(a[7]), .B(b[26]), .Z(n44499) );
  XOR U45354 ( .A(n44505), .B(n44506), .Z(n44312) );
  ANDN U45355 ( .B(n44507), .A(n44508), .Z(n44505) );
  AND U45356 ( .A(a[8]), .B(b[25]), .Z(n44504) );
  XOR U45357 ( .A(n44510), .B(n44511), .Z(n44317) );
  ANDN U45358 ( .B(n44512), .A(n44513), .Z(n44510) );
  AND U45359 ( .A(a[9]), .B(b[24]), .Z(n44509) );
  XOR U45360 ( .A(n44515), .B(n44516), .Z(n44322) );
  ANDN U45361 ( .B(n44517), .A(n44518), .Z(n44515) );
  AND U45362 ( .A(a[10]), .B(b[23]), .Z(n44514) );
  XOR U45363 ( .A(n44520), .B(n44521), .Z(n44327) );
  ANDN U45364 ( .B(n44522), .A(n44523), .Z(n44520) );
  AND U45365 ( .A(a[11]), .B(b[22]), .Z(n44519) );
  XOR U45366 ( .A(n44525), .B(n44526), .Z(n44332) );
  ANDN U45367 ( .B(n44527), .A(n44528), .Z(n44525) );
  AND U45368 ( .A(a[12]), .B(b[21]), .Z(n44524) );
  XOR U45369 ( .A(n44530), .B(n44531), .Z(n44337) );
  ANDN U45370 ( .B(n44532), .A(n44533), .Z(n44530) );
  AND U45371 ( .A(a[13]), .B(b[20]), .Z(n44529) );
  XOR U45372 ( .A(n44535), .B(n44536), .Z(n44342) );
  ANDN U45373 ( .B(n44537), .A(n44538), .Z(n44535) );
  AND U45374 ( .A(a[14]), .B(b[19]), .Z(n44534) );
  XOR U45375 ( .A(n44540), .B(n44541), .Z(n44347) );
  ANDN U45376 ( .B(n44542), .A(n44543), .Z(n44540) );
  AND U45377 ( .A(a[15]), .B(b[18]), .Z(n44539) );
  XOR U45378 ( .A(n44545), .B(n44546), .Z(n44352) );
  ANDN U45379 ( .B(n44547), .A(n44548), .Z(n44545) );
  AND U45380 ( .A(a[16]), .B(b[17]), .Z(n44544) );
  XOR U45381 ( .A(n44550), .B(n44551), .Z(n44357) );
  ANDN U45382 ( .B(n44552), .A(n44553), .Z(n44550) );
  AND U45383 ( .A(a[17]), .B(b[16]), .Z(n44549) );
  XOR U45384 ( .A(n44555), .B(n44556), .Z(n44362) );
  ANDN U45385 ( .B(n44557), .A(n44558), .Z(n44555) );
  AND U45386 ( .A(a[18]), .B(b[15]), .Z(n44554) );
  XOR U45387 ( .A(n44560), .B(n44561), .Z(n44367) );
  ANDN U45388 ( .B(n44562), .A(n44563), .Z(n44560) );
  AND U45389 ( .A(a[19]), .B(b[14]), .Z(n44559) );
  XOR U45390 ( .A(n44565), .B(n44566), .Z(n44372) );
  ANDN U45391 ( .B(n44567), .A(n44568), .Z(n44565) );
  AND U45392 ( .A(a[20]), .B(b[13]), .Z(n44564) );
  XOR U45393 ( .A(n44570), .B(n44571), .Z(n44377) );
  ANDN U45394 ( .B(n44572), .A(n44573), .Z(n44570) );
  AND U45395 ( .A(a[21]), .B(b[12]), .Z(n44569) );
  XOR U45396 ( .A(n44575), .B(n44576), .Z(n44382) );
  ANDN U45397 ( .B(n44577), .A(n44578), .Z(n44575) );
  AND U45398 ( .A(a[22]), .B(b[11]), .Z(n44574) );
  XOR U45399 ( .A(n44580), .B(n44581), .Z(n44387) );
  ANDN U45400 ( .B(n44582), .A(n44583), .Z(n44580) );
  AND U45401 ( .A(a[23]), .B(b[10]), .Z(n44579) );
  XOR U45402 ( .A(n44585), .B(n44586), .Z(n44392) );
  ANDN U45403 ( .B(n44587), .A(n44588), .Z(n44585) );
  AND U45404 ( .A(b[9]), .B(a[24]), .Z(n44584) );
  XOR U45405 ( .A(n44590), .B(n44591), .Z(n44397) );
  ANDN U45406 ( .B(n44592), .A(n44593), .Z(n44590) );
  AND U45407 ( .A(b[8]), .B(a[25]), .Z(n44589) );
  XOR U45408 ( .A(n44595), .B(n44596), .Z(n44402) );
  ANDN U45409 ( .B(n44597), .A(n44598), .Z(n44595) );
  AND U45410 ( .A(b[7]), .B(a[26]), .Z(n44594) );
  XOR U45411 ( .A(n44600), .B(n44601), .Z(n44407) );
  ANDN U45412 ( .B(n44602), .A(n44603), .Z(n44600) );
  AND U45413 ( .A(b[6]), .B(a[27]), .Z(n44599) );
  XOR U45414 ( .A(n44605), .B(n44606), .Z(n44412) );
  ANDN U45415 ( .B(n44607), .A(n44608), .Z(n44605) );
  AND U45416 ( .A(b[5]), .B(a[28]), .Z(n44604) );
  XOR U45417 ( .A(n44610), .B(n44611), .Z(n44417) );
  ANDN U45418 ( .B(n44612), .A(n44613), .Z(n44610) );
  AND U45419 ( .A(b[4]), .B(a[29]), .Z(n44609) );
  XOR U45420 ( .A(n44615), .B(n44616), .Z(n44422) );
  ANDN U45421 ( .B(n44434), .A(n44435), .Z(n44615) );
  AND U45422 ( .A(b[2]), .B(a[30]), .Z(n44617) );
  XNOR U45423 ( .A(n44612), .B(n44616), .Z(n44618) );
  XOR U45424 ( .A(n44619), .B(n44620), .Z(n44616) );
  OR U45425 ( .A(n44437), .B(n44438), .Z(n44620) );
  XNOR U45426 ( .A(n44622), .B(n44623), .Z(n44621) );
  XOR U45427 ( .A(n44622), .B(n44625), .Z(n44437) );
  NAND U45428 ( .A(b[1]), .B(a[30]), .Z(n44625) );
  IV U45429 ( .A(n44619), .Z(n44622) );
  NANDN U45430 ( .A(n153), .B(n154), .Z(n44619) );
  XOR U45431 ( .A(n44626), .B(n44627), .Z(n154) );
  NAND U45432 ( .A(a[30]), .B(b[0]), .Z(n153) );
  XNOR U45433 ( .A(n44607), .B(n44611), .Z(n44628) );
  XNOR U45434 ( .A(n44602), .B(n44606), .Z(n44629) );
  XNOR U45435 ( .A(n44597), .B(n44601), .Z(n44630) );
  XNOR U45436 ( .A(n44592), .B(n44596), .Z(n44631) );
  XNOR U45437 ( .A(n44587), .B(n44591), .Z(n44632) );
  XNOR U45438 ( .A(n44582), .B(n44586), .Z(n44633) );
  XNOR U45439 ( .A(n44577), .B(n44581), .Z(n44634) );
  XNOR U45440 ( .A(n44572), .B(n44576), .Z(n44635) );
  XNOR U45441 ( .A(n44567), .B(n44571), .Z(n44636) );
  XNOR U45442 ( .A(n44562), .B(n44566), .Z(n44637) );
  XNOR U45443 ( .A(n44557), .B(n44561), .Z(n44638) );
  XNOR U45444 ( .A(n44552), .B(n44556), .Z(n44639) );
  XNOR U45445 ( .A(n44547), .B(n44551), .Z(n44640) );
  XNOR U45446 ( .A(n44542), .B(n44546), .Z(n44641) );
  XNOR U45447 ( .A(n44537), .B(n44541), .Z(n44642) );
  XNOR U45448 ( .A(n44532), .B(n44536), .Z(n44643) );
  XNOR U45449 ( .A(n44527), .B(n44531), .Z(n44644) );
  XNOR U45450 ( .A(n44522), .B(n44526), .Z(n44645) );
  XNOR U45451 ( .A(n44517), .B(n44521), .Z(n44646) );
  XNOR U45452 ( .A(n44512), .B(n44516), .Z(n44647) );
  XNOR U45453 ( .A(n44507), .B(n44511), .Z(n44648) );
  XNOR U45454 ( .A(n44502), .B(n44506), .Z(n44649) );
  XNOR U45455 ( .A(n44497), .B(n44501), .Z(n44650) );
  XNOR U45456 ( .A(n44492), .B(n44496), .Z(n44651) );
  XNOR U45457 ( .A(n44487), .B(n44491), .Z(n44652) );
  XNOR U45458 ( .A(n44482), .B(n44486), .Z(n44653) );
  XNOR U45459 ( .A(n44477), .B(n44481), .Z(n44654) );
  XNOR U45460 ( .A(n44472), .B(n44476), .Z(n44655) );
  XOR U45461 ( .A(n44656), .B(n44471), .Z(n44472) );
  AND U45462 ( .A(a[0]), .B(b[32]), .Z(n44656) );
  XNOR U45463 ( .A(n44657), .B(n44471), .Z(n44473) );
  XNOR U45464 ( .A(n44658), .B(n44659), .Z(n44471) );
  ANDN U45465 ( .B(n44660), .A(n44661), .Z(n44658) );
  AND U45466 ( .A(a[1]), .B(b[31]), .Z(n44657) );
  XOR U45467 ( .A(n44663), .B(n44664), .Z(n44476) );
  ANDN U45468 ( .B(n44665), .A(n44666), .Z(n44663) );
  AND U45469 ( .A(a[2]), .B(b[30]), .Z(n44662) );
  XOR U45470 ( .A(n44668), .B(n44669), .Z(n44481) );
  ANDN U45471 ( .B(n44670), .A(n44671), .Z(n44668) );
  AND U45472 ( .A(a[3]), .B(b[29]), .Z(n44667) );
  XOR U45473 ( .A(n44673), .B(n44674), .Z(n44486) );
  ANDN U45474 ( .B(n44675), .A(n44676), .Z(n44673) );
  AND U45475 ( .A(a[4]), .B(b[28]), .Z(n44672) );
  XOR U45476 ( .A(n44678), .B(n44679), .Z(n44491) );
  ANDN U45477 ( .B(n44680), .A(n44681), .Z(n44678) );
  AND U45478 ( .A(a[5]), .B(b[27]), .Z(n44677) );
  XOR U45479 ( .A(n44683), .B(n44684), .Z(n44496) );
  ANDN U45480 ( .B(n44685), .A(n44686), .Z(n44683) );
  AND U45481 ( .A(a[6]), .B(b[26]), .Z(n44682) );
  XOR U45482 ( .A(n44688), .B(n44689), .Z(n44501) );
  ANDN U45483 ( .B(n44690), .A(n44691), .Z(n44688) );
  AND U45484 ( .A(a[7]), .B(b[25]), .Z(n44687) );
  XOR U45485 ( .A(n44693), .B(n44694), .Z(n44506) );
  ANDN U45486 ( .B(n44695), .A(n44696), .Z(n44693) );
  AND U45487 ( .A(a[8]), .B(b[24]), .Z(n44692) );
  XOR U45488 ( .A(n44698), .B(n44699), .Z(n44511) );
  ANDN U45489 ( .B(n44700), .A(n44701), .Z(n44698) );
  AND U45490 ( .A(a[9]), .B(b[23]), .Z(n44697) );
  XOR U45491 ( .A(n44703), .B(n44704), .Z(n44516) );
  ANDN U45492 ( .B(n44705), .A(n44706), .Z(n44703) );
  AND U45493 ( .A(a[10]), .B(b[22]), .Z(n44702) );
  XOR U45494 ( .A(n44708), .B(n44709), .Z(n44521) );
  ANDN U45495 ( .B(n44710), .A(n44711), .Z(n44708) );
  AND U45496 ( .A(a[11]), .B(b[21]), .Z(n44707) );
  XOR U45497 ( .A(n44713), .B(n44714), .Z(n44526) );
  ANDN U45498 ( .B(n44715), .A(n44716), .Z(n44713) );
  AND U45499 ( .A(a[12]), .B(b[20]), .Z(n44712) );
  XOR U45500 ( .A(n44718), .B(n44719), .Z(n44531) );
  ANDN U45501 ( .B(n44720), .A(n44721), .Z(n44718) );
  AND U45502 ( .A(a[13]), .B(b[19]), .Z(n44717) );
  XOR U45503 ( .A(n44723), .B(n44724), .Z(n44536) );
  ANDN U45504 ( .B(n44725), .A(n44726), .Z(n44723) );
  AND U45505 ( .A(a[14]), .B(b[18]), .Z(n44722) );
  XOR U45506 ( .A(n44728), .B(n44729), .Z(n44541) );
  ANDN U45507 ( .B(n44730), .A(n44731), .Z(n44728) );
  AND U45508 ( .A(a[15]), .B(b[17]), .Z(n44727) );
  XOR U45509 ( .A(n44733), .B(n44734), .Z(n44546) );
  ANDN U45510 ( .B(n44735), .A(n44736), .Z(n44733) );
  AND U45511 ( .A(a[16]), .B(b[16]), .Z(n44732) );
  XOR U45512 ( .A(n44738), .B(n44739), .Z(n44551) );
  ANDN U45513 ( .B(n44740), .A(n44741), .Z(n44738) );
  AND U45514 ( .A(a[17]), .B(b[15]), .Z(n44737) );
  XOR U45515 ( .A(n44743), .B(n44744), .Z(n44556) );
  ANDN U45516 ( .B(n44745), .A(n44746), .Z(n44743) );
  AND U45517 ( .A(a[18]), .B(b[14]), .Z(n44742) );
  XOR U45518 ( .A(n44748), .B(n44749), .Z(n44561) );
  ANDN U45519 ( .B(n44750), .A(n44751), .Z(n44748) );
  AND U45520 ( .A(a[19]), .B(b[13]), .Z(n44747) );
  XOR U45521 ( .A(n44753), .B(n44754), .Z(n44566) );
  ANDN U45522 ( .B(n44755), .A(n44756), .Z(n44753) );
  AND U45523 ( .A(a[20]), .B(b[12]), .Z(n44752) );
  XOR U45524 ( .A(n44758), .B(n44759), .Z(n44571) );
  ANDN U45525 ( .B(n44760), .A(n44761), .Z(n44758) );
  AND U45526 ( .A(a[21]), .B(b[11]), .Z(n44757) );
  XOR U45527 ( .A(n44763), .B(n44764), .Z(n44576) );
  ANDN U45528 ( .B(n44765), .A(n44766), .Z(n44763) );
  AND U45529 ( .A(a[22]), .B(b[10]), .Z(n44762) );
  XOR U45530 ( .A(n44768), .B(n44769), .Z(n44581) );
  ANDN U45531 ( .B(n44770), .A(n44771), .Z(n44768) );
  AND U45532 ( .A(b[9]), .B(a[23]), .Z(n44767) );
  XOR U45533 ( .A(n44773), .B(n44774), .Z(n44586) );
  ANDN U45534 ( .B(n44775), .A(n44776), .Z(n44773) );
  AND U45535 ( .A(b[8]), .B(a[24]), .Z(n44772) );
  XOR U45536 ( .A(n44778), .B(n44779), .Z(n44591) );
  ANDN U45537 ( .B(n44780), .A(n44781), .Z(n44778) );
  AND U45538 ( .A(b[7]), .B(a[25]), .Z(n44777) );
  XOR U45539 ( .A(n44783), .B(n44784), .Z(n44596) );
  ANDN U45540 ( .B(n44785), .A(n44786), .Z(n44783) );
  AND U45541 ( .A(b[6]), .B(a[26]), .Z(n44782) );
  XOR U45542 ( .A(n44788), .B(n44789), .Z(n44601) );
  ANDN U45543 ( .B(n44790), .A(n44791), .Z(n44788) );
  AND U45544 ( .A(b[5]), .B(a[27]), .Z(n44787) );
  XOR U45545 ( .A(n44793), .B(n44794), .Z(n44606) );
  ANDN U45546 ( .B(n44795), .A(n44796), .Z(n44793) );
  AND U45547 ( .A(b[4]), .B(a[28]), .Z(n44792) );
  XOR U45548 ( .A(n44798), .B(n44799), .Z(n44611) );
  ANDN U45549 ( .B(n44623), .A(n44624), .Z(n44798) );
  AND U45550 ( .A(b[2]), .B(a[29]), .Z(n44800) );
  XNOR U45551 ( .A(n44795), .B(n44799), .Z(n44801) );
  XOR U45552 ( .A(n44802), .B(n44803), .Z(n44799) );
  OR U45553 ( .A(n44626), .B(n44627), .Z(n44803) );
  XNOR U45554 ( .A(n44805), .B(n44806), .Z(n44804) );
  XOR U45555 ( .A(n44805), .B(n44808), .Z(n44626) );
  NAND U45556 ( .A(b[1]), .B(a[29]), .Z(n44808) );
  IV U45557 ( .A(n44802), .Z(n44805) );
  NANDN U45558 ( .A(n157), .B(n158), .Z(n44802) );
  XOR U45559 ( .A(n44809), .B(n44810), .Z(n158) );
  NAND U45560 ( .A(a[29]), .B(b[0]), .Z(n157) );
  XNOR U45561 ( .A(n44790), .B(n44794), .Z(n44811) );
  XNOR U45562 ( .A(n44785), .B(n44789), .Z(n44812) );
  XNOR U45563 ( .A(n44780), .B(n44784), .Z(n44813) );
  XNOR U45564 ( .A(n44775), .B(n44779), .Z(n44814) );
  XNOR U45565 ( .A(n44770), .B(n44774), .Z(n44815) );
  XNOR U45566 ( .A(n44765), .B(n44769), .Z(n44816) );
  XNOR U45567 ( .A(n44760), .B(n44764), .Z(n44817) );
  XNOR U45568 ( .A(n44755), .B(n44759), .Z(n44818) );
  XNOR U45569 ( .A(n44750), .B(n44754), .Z(n44819) );
  XNOR U45570 ( .A(n44745), .B(n44749), .Z(n44820) );
  XNOR U45571 ( .A(n44740), .B(n44744), .Z(n44821) );
  XNOR U45572 ( .A(n44735), .B(n44739), .Z(n44822) );
  XNOR U45573 ( .A(n44730), .B(n44734), .Z(n44823) );
  XNOR U45574 ( .A(n44725), .B(n44729), .Z(n44824) );
  XNOR U45575 ( .A(n44720), .B(n44724), .Z(n44825) );
  XNOR U45576 ( .A(n44715), .B(n44719), .Z(n44826) );
  XNOR U45577 ( .A(n44710), .B(n44714), .Z(n44827) );
  XNOR U45578 ( .A(n44705), .B(n44709), .Z(n44828) );
  XNOR U45579 ( .A(n44700), .B(n44704), .Z(n44829) );
  XNOR U45580 ( .A(n44695), .B(n44699), .Z(n44830) );
  XNOR U45581 ( .A(n44690), .B(n44694), .Z(n44831) );
  XNOR U45582 ( .A(n44685), .B(n44689), .Z(n44832) );
  XNOR U45583 ( .A(n44680), .B(n44684), .Z(n44833) );
  XNOR U45584 ( .A(n44675), .B(n44679), .Z(n44834) );
  XNOR U45585 ( .A(n44670), .B(n44674), .Z(n44835) );
  XNOR U45586 ( .A(n44665), .B(n44669), .Z(n44836) );
  XNOR U45587 ( .A(n44660), .B(n44664), .Z(n44837) );
  XNOR U45588 ( .A(n44838), .B(n44659), .Z(n44660) );
  AND U45589 ( .A(a[0]), .B(b[31]), .Z(n44838) );
  XOR U45590 ( .A(n44839), .B(n44659), .Z(n44661) );
  XNOR U45591 ( .A(n44840), .B(n44841), .Z(n44659) );
  ANDN U45592 ( .B(n44842), .A(n44843), .Z(n44840) );
  AND U45593 ( .A(a[1]), .B(b[30]), .Z(n44839) );
  XOR U45594 ( .A(n44845), .B(n44846), .Z(n44664) );
  ANDN U45595 ( .B(n44847), .A(n44848), .Z(n44845) );
  AND U45596 ( .A(a[2]), .B(b[29]), .Z(n44844) );
  XOR U45597 ( .A(n44850), .B(n44851), .Z(n44669) );
  ANDN U45598 ( .B(n44852), .A(n44853), .Z(n44850) );
  AND U45599 ( .A(a[3]), .B(b[28]), .Z(n44849) );
  XOR U45600 ( .A(n44855), .B(n44856), .Z(n44674) );
  ANDN U45601 ( .B(n44857), .A(n44858), .Z(n44855) );
  AND U45602 ( .A(a[4]), .B(b[27]), .Z(n44854) );
  XOR U45603 ( .A(n44860), .B(n44861), .Z(n44679) );
  ANDN U45604 ( .B(n44862), .A(n44863), .Z(n44860) );
  AND U45605 ( .A(a[5]), .B(b[26]), .Z(n44859) );
  XOR U45606 ( .A(n44865), .B(n44866), .Z(n44684) );
  ANDN U45607 ( .B(n44867), .A(n44868), .Z(n44865) );
  AND U45608 ( .A(a[6]), .B(b[25]), .Z(n44864) );
  XOR U45609 ( .A(n44870), .B(n44871), .Z(n44689) );
  ANDN U45610 ( .B(n44872), .A(n44873), .Z(n44870) );
  AND U45611 ( .A(a[7]), .B(b[24]), .Z(n44869) );
  XOR U45612 ( .A(n44875), .B(n44876), .Z(n44694) );
  ANDN U45613 ( .B(n44877), .A(n44878), .Z(n44875) );
  AND U45614 ( .A(a[8]), .B(b[23]), .Z(n44874) );
  XOR U45615 ( .A(n44880), .B(n44881), .Z(n44699) );
  ANDN U45616 ( .B(n44882), .A(n44883), .Z(n44880) );
  AND U45617 ( .A(a[9]), .B(b[22]), .Z(n44879) );
  XOR U45618 ( .A(n44885), .B(n44886), .Z(n44704) );
  ANDN U45619 ( .B(n44887), .A(n44888), .Z(n44885) );
  AND U45620 ( .A(a[10]), .B(b[21]), .Z(n44884) );
  XOR U45621 ( .A(n44890), .B(n44891), .Z(n44709) );
  ANDN U45622 ( .B(n44892), .A(n44893), .Z(n44890) );
  AND U45623 ( .A(a[11]), .B(b[20]), .Z(n44889) );
  XOR U45624 ( .A(n44895), .B(n44896), .Z(n44714) );
  ANDN U45625 ( .B(n44897), .A(n44898), .Z(n44895) );
  AND U45626 ( .A(a[12]), .B(b[19]), .Z(n44894) );
  XOR U45627 ( .A(n44900), .B(n44901), .Z(n44719) );
  ANDN U45628 ( .B(n44902), .A(n44903), .Z(n44900) );
  AND U45629 ( .A(a[13]), .B(b[18]), .Z(n44899) );
  XOR U45630 ( .A(n44905), .B(n44906), .Z(n44724) );
  ANDN U45631 ( .B(n44907), .A(n44908), .Z(n44905) );
  AND U45632 ( .A(a[14]), .B(b[17]), .Z(n44904) );
  XOR U45633 ( .A(n44910), .B(n44911), .Z(n44729) );
  ANDN U45634 ( .B(n44912), .A(n44913), .Z(n44910) );
  AND U45635 ( .A(a[15]), .B(b[16]), .Z(n44909) );
  XOR U45636 ( .A(n44915), .B(n44916), .Z(n44734) );
  ANDN U45637 ( .B(n44917), .A(n44918), .Z(n44915) );
  AND U45638 ( .A(a[16]), .B(b[15]), .Z(n44914) );
  XOR U45639 ( .A(n44920), .B(n44921), .Z(n44739) );
  ANDN U45640 ( .B(n44922), .A(n44923), .Z(n44920) );
  AND U45641 ( .A(a[17]), .B(b[14]), .Z(n44919) );
  XOR U45642 ( .A(n44925), .B(n44926), .Z(n44744) );
  ANDN U45643 ( .B(n44927), .A(n44928), .Z(n44925) );
  AND U45644 ( .A(a[18]), .B(b[13]), .Z(n44924) );
  XOR U45645 ( .A(n44930), .B(n44931), .Z(n44749) );
  ANDN U45646 ( .B(n44932), .A(n44933), .Z(n44930) );
  AND U45647 ( .A(a[19]), .B(b[12]), .Z(n44929) );
  XOR U45648 ( .A(n44935), .B(n44936), .Z(n44754) );
  ANDN U45649 ( .B(n44937), .A(n44938), .Z(n44935) );
  AND U45650 ( .A(a[20]), .B(b[11]), .Z(n44934) );
  XOR U45651 ( .A(n44940), .B(n44941), .Z(n44759) );
  ANDN U45652 ( .B(n44942), .A(n44943), .Z(n44940) );
  AND U45653 ( .A(a[21]), .B(b[10]), .Z(n44939) );
  XOR U45654 ( .A(n44945), .B(n44946), .Z(n44764) );
  ANDN U45655 ( .B(n44947), .A(n44948), .Z(n44945) );
  AND U45656 ( .A(b[9]), .B(a[22]), .Z(n44944) );
  XOR U45657 ( .A(n44950), .B(n44951), .Z(n44769) );
  ANDN U45658 ( .B(n44952), .A(n44953), .Z(n44950) );
  AND U45659 ( .A(b[8]), .B(a[23]), .Z(n44949) );
  XOR U45660 ( .A(n44955), .B(n44956), .Z(n44774) );
  ANDN U45661 ( .B(n44957), .A(n44958), .Z(n44955) );
  AND U45662 ( .A(b[7]), .B(a[24]), .Z(n44954) );
  XOR U45663 ( .A(n44960), .B(n44961), .Z(n44779) );
  ANDN U45664 ( .B(n44962), .A(n44963), .Z(n44960) );
  AND U45665 ( .A(b[6]), .B(a[25]), .Z(n44959) );
  XOR U45666 ( .A(n44965), .B(n44966), .Z(n44784) );
  ANDN U45667 ( .B(n44967), .A(n44968), .Z(n44965) );
  AND U45668 ( .A(b[5]), .B(a[26]), .Z(n44964) );
  XOR U45669 ( .A(n44970), .B(n44971), .Z(n44789) );
  ANDN U45670 ( .B(n44972), .A(n44973), .Z(n44970) );
  AND U45671 ( .A(b[4]), .B(a[27]), .Z(n44969) );
  XOR U45672 ( .A(n44975), .B(n44976), .Z(n44794) );
  ANDN U45673 ( .B(n44806), .A(n44807), .Z(n44975) );
  AND U45674 ( .A(b[2]), .B(a[28]), .Z(n44977) );
  XNOR U45675 ( .A(n44972), .B(n44976), .Z(n44978) );
  XOR U45676 ( .A(n44979), .B(n44980), .Z(n44976) );
  OR U45677 ( .A(n44809), .B(n44810), .Z(n44980) );
  XNOR U45678 ( .A(n44982), .B(n44983), .Z(n44981) );
  XOR U45679 ( .A(n44982), .B(n44985), .Z(n44809) );
  NAND U45680 ( .A(b[1]), .B(a[28]), .Z(n44985) );
  IV U45681 ( .A(n44979), .Z(n44982) );
  NANDN U45682 ( .A(n159), .B(n160), .Z(n44979) );
  XOR U45683 ( .A(n44986), .B(n44987), .Z(n160) );
  NAND U45684 ( .A(a[28]), .B(b[0]), .Z(n159) );
  XNOR U45685 ( .A(n44967), .B(n44971), .Z(n44988) );
  XNOR U45686 ( .A(n44962), .B(n44966), .Z(n44989) );
  XNOR U45687 ( .A(n44957), .B(n44961), .Z(n44990) );
  XNOR U45688 ( .A(n44952), .B(n44956), .Z(n44991) );
  XNOR U45689 ( .A(n44947), .B(n44951), .Z(n44992) );
  XNOR U45690 ( .A(n44942), .B(n44946), .Z(n44993) );
  XNOR U45691 ( .A(n44937), .B(n44941), .Z(n44994) );
  XNOR U45692 ( .A(n44932), .B(n44936), .Z(n44995) );
  XNOR U45693 ( .A(n44927), .B(n44931), .Z(n44996) );
  XNOR U45694 ( .A(n44922), .B(n44926), .Z(n44997) );
  XNOR U45695 ( .A(n44917), .B(n44921), .Z(n44998) );
  XNOR U45696 ( .A(n44912), .B(n44916), .Z(n44999) );
  XNOR U45697 ( .A(n44907), .B(n44911), .Z(n45000) );
  XNOR U45698 ( .A(n44902), .B(n44906), .Z(n45001) );
  XNOR U45699 ( .A(n44897), .B(n44901), .Z(n45002) );
  XNOR U45700 ( .A(n44892), .B(n44896), .Z(n45003) );
  XNOR U45701 ( .A(n44887), .B(n44891), .Z(n45004) );
  XNOR U45702 ( .A(n44882), .B(n44886), .Z(n45005) );
  XNOR U45703 ( .A(n44877), .B(n44881), .Z(n45006) );
  XNOR U45704 ( .A(n44872), .B(n44876), .Z(n45007) );
  XNOR U45705 ( .A(n44867), .B(n44871), .Z(n45008) );
  XNOR U45706 ( .A(n44862), .B(n44866), .Z(n45009) );
  XNOR U45707 ( .A(n44857), .B(n44861), .Z(n45010) );
  XNOR U45708 ( .A(n44852), .B(n44856), .Z(n45011) );
  XNOR U45709 ( .A(n44847), .B(n44851), .Z(n45012) );
  XNOR U45710 ( .A(n44842), .B(n44846), .Z(n45013) );
  XOR U45711 ( .A(n45014), .B(n44841), .Z(n44842) );
  AND U45712 ( .A(a[0]), .B(b[30]), .Z(n45014) );
  XNOR U45713 ( .A(n45015), .B(n44841), .Z(n44843) );
  XNOR U45714 ( .A(n45016), .B(n45017), .Z(n44841) );
  ANDN U45715 ( .B(n45018), .A(n45019), .Z(n45016) );
  AND U45716 ( .A(a[1]), .B(b[29]), .Z(n45015) );
  XOR U45717 ( .A(n45021), .B(n45022), .Z(n44846) );
  ANDN U45718 ( .B(n45023), .A(n45024), .Z(n45021) );
  AND U45719 ( .A(a[2]), .B(b[28]), .Z(n45020) );
  XOR U45720 ( .A(n45026), .B(n45027), .Z(n44851) );
  ANDN U45721 ( .B(n45028), .A(n45029), .Z(n45026) );
  AND U45722 ( .A(a[3]), .B(b[27]), .Z(n45025) );
  XOR U45723 ( .A(n45031), .B(n45032), .Z(n44856) );
  ANDN U45724 ( .B(n45033), .A(n45034), .Z(n45031) );
  AND U45725 ( .A(a[4]), .B(b[26]), .Z(n45030) );
  XOR U45726 ( .A(n45036), .B(n45037), .Z(n44861) );
  ANDN U45727 ( .B(n45038), .A(n45039), .Z(n45036) );
  AND U45728 ( .A(a[5]), .B(b[25]), .Z(n45035) );
  XOR U45729 ( .A(n45041), .B(n45042), .Z(n44866) );
  ANDN U45730 ( .B(n45043), .A(n45044), .Z(n45041) );
  AND U45731 ( .A(a[6]), .B(b[24]), .Z(n45040) );
  XOR U45732 ( .A(n45046), .B(n45047), .Z(n44871) );
  ANDN U45733 ( .B(n45048), .A(n45049), .Z(n45046) );
  AND U45734 ( .A(a[7]), .B(b[23]), .Z(n45045) );
  XOR U45735 ( .A(n45051), .B(n45052), .Z(n44876) );
  ANDN U45736 ( .B(n45053), .A(n45054), .Z(n45051) );
  AND U45737 ( .A(a[8]), .B(b[22]), .Z(n45050) );
  XOR U45738 ( .A(n45056), .B(n45057), .Z(n44881) );
  ANDN U45739 ( .B(n45058), .A(n45059), .Z(n45056) );
  AND U45740 ( .A(a[9]), .B(b[21]), .Z(n45055) );
  XOR U45741 ( .A(n45061), .B(n45062), .Z(n44886) );
  ANDN U45742 ( .B(n45063), .A(n45064), .Z(n45061) );
  AND U45743 ( .A(a[10]), .B(b[20]), .Z(n45060) );
  XOR U45744 ( .A(n45066), .B(n45067), .Z(n44891) );
  ANDN U45745 ( .B(n45068), .A(n45069), .Z(n45066) );
  AND U45746 ( .A(a[11]), .B(b[19]), .Z(n45065) );
  XOR U45747 ( .A(n45071), .B(n45072), .Z(n44896) );
  ANDN U45748 ( .B(n45073), .A(n45074), .Z(n45071) );
  AND U45749 ( .A(a[12]), .B(b[18]), .Z(n45070) );
  XOR U45750 ( .A(n45076), .B(n45077), .Z(n44901) );
  ANDN U45751 ( .B(n45078), .A(n45079), .Z(n45076) );
  AND U45752 ( .A(a[13]), .B(b[17]), .Z(n45075) );
  XOR U45753 ( .A(n45081), .B(n45082), .Z(n44906) );
  ANDN U45754 ( .B(n45083), .A(n45084), .Z(n45081) );
  AND U45755 ( .A(a[14]), .B(b[16]), .Z(n45080) );
  XOR U45756 ( .A(n45086), .B(n45087), .Z(n44911) );
  ANDN U45757 ( .B(n45088), .A(n45089), .Z(n45086) );
  AND U45758 ( .A(a[15]), .B(b[15]), .Z(n45085) );
  XOR U45759 ( .A(n45091), .B(n45092), .Z(n44916) );
  ANDN U45760 ( .B(n45093), .A(n45094), .Z(n45091) );
  AND U45761 ( .A(a[16]), .B(b[14]), .Z(n45090) );
  XOR U45762 ( .A(n45096), .B(n45097), .Z(n44921) );
  ANDN U45763 ( .B(n45098), .A(n45099), .Z(n45096) );
  AND U45764 ( .A(a[17]), .B(b[13]), .Z(n45095) );
  XOR U45765 ( .A(n45101), .B(n45102), .Z(n44926) );
  ANDN U45766 ( .B(n45103), .A(n45104), .Z(n45101) );
  AND U45767 ( .A(a[18]), .B(b[12]), .Z(n45100) );
  XOR U45768 ( .A(n45106), .B(n45107), .Z(n44931) );
  ANDN U45769 ( .B(n45108), .A(n45109), .Z(n45106) );
  AND U45770 ( .A(a[19]), .B(b[11]), .Z(n45105) );
  XOR U45771 ( .A(n45111), .B(n45112), .Z(n44936) );
  ANDN U45772 ( .B(n45113), .A(n45114), .Z(n45111) );
  AND U45773 ( .A(a[20]), .B(b[10]), .Z(n45110) );
  XOR U45774 ( .A(n45116), .B(n45117), .Z(n44941) );
  ANDN U45775 ( .B(n45118), .A(n45119), .Z(n45116) );
  AND U45776 ( .A(b[9]), .B(a[21]), .Z(n45115) );
  XOR U45777 ( .A(n45121), .B(n45122), .Z(n44946) );
  ANDN U45778 ( .B(n45123), .A(n45124), .Z(n45121) );
  AND U45779 ( .A(b[8]), .B(a[22]), .Z(n45120) );
  XOR U45780 ( .A(n45126), .B(n45127), .Z(n44951) );
  ANDN U45781 ( .B(n45128), .A(n45129), .Z(n45126) );
  AND U45782 ( .A(b[7]), .B(a[23]), .Z(n45125) );
  XOR U45783 ( .A(n45131), .B(n45132), .Z(n44956) );
  ANDN U45784 ( .B(n45133), .A(n45134), .Z(n45131) );
  AND U45785 ( .A(b[6]), .B(a[24]), .Z(n45130) );
  XOR U45786 ( .A(n45136), .B(n45137), .Z(n44961) );
  ANDN U45787 ( .B(n45138), .A(n45139), .Z(n45136) );
  AND U45788 ( .A(b[5]), .B(a[25]), .Z(n45135) );
  XOR U45789 ( .A(n45141), .B(n45142), .Z(n44966) );
  ANDN U45790 ( .B(n45143), .A(n45144), .Z(n45141) );
  AND U45791 ( .A(b[4]), .B(a[26]), .Z(n45140) );
  XOR U45792 ( .A(n45146), .B(n45147), .Z(n44971) );
  ANDN U45793 ( .B(n44983), .A(n44984), .Z(n45146) );
  AND U45794 ( .A(b[2]), .B(a[27]), .Z(n45148) );
  XNOR U45795 ( .A(n45143), .B(n45147), .Z(n45149) );
  XOR U45796 ( .A(n45150), .B(n45151), .Z(n45147) );
  OR U45797 ( .A(n44986), .B(n44987), .Z(n45151) );
  XNOR U45798 ( .A(n45153), .B(n45154), .Z(n45152) );
  XOR U45799 ( .A(n45153), .B(n45156), .Z(n44986) );
  NAND U45800 ( .A(b[1]), .B(a[27]), .Z(n45156) );
  IV U45801 ( .A(n45150), .Z(n45153) );
  NANDN U45802 ( .A(n161), .B(n162), .Z(n45150) );
  XOR U45803 ( .A(n45157), .B(n45158), .Z(n162) );
  NAND U45804 ( .A(a[27]), .B(b[0]), .Z(n161) );
  XNOR U45805 ( .A(n45138), .B(n45142), .Z(n45159) );
  XNOR U45806 ( .A(n45133), .B(n45137), .Z(n45160) );
  XNOR U45807 ( .A(n45128), .B(n45132), .Z(n45161) );
  XNOR U45808 ( .A(n45123), .B(n45127), .Z(n45162) );
  XNOR U45809 ( .A(n45118), .B(n45122), .Z(n45163) );
  XNOR U45810 ( .A(n45113), .B(n45117), .Z(n45164) );
  XNOR U45811 ( .A(n45108), .B(n45112), .Z(n45165) );
  XNOR U45812 ( .A(n45103), .B(n45107), .Z(n45166) );
  XNOR U45813 ( .A(n45098), .B(n45102), .Z(n45167) );
  XNOR U45814 ( .A(n45093), .B(n45097), .Z(n45168) );
  XNOR U45815 ( .A(n45088), .B(n45092), .Z(n45169) );
  XNOR U45816 ( .A(n45083), .B(n45087), .Z(n45170) );
  XNOR U45817 ( .A(n45078), .B(n45082), .Z(n45171) );
  XNOR U45818 ( .A(n45073), .B(n45077), .Z(n45172) );
  XNOR U45819 ( .A(n45068), .B(n45072), .Z(n45173) );
  XNOR U45820 ( .A(n45063), .B(n45067), .Z(n45174) );
  XNOR U45821 ( .A(n45058), .B(n45062), .Z(n45175) );
  XNOR U45822 ( .A(n45053), .B(n45057), .Z(n45176) );
  XNOR U45823 ( .A(n45048), .B(n45052), .Z(n45177) );
  XNOR U45824 ( .A(n45043), .B(n45047), .Z(n45178) );
  XNOR U45825 ( .A(n45038), .B(n45042), .Z(n45179) );
  XNOR U45826 ( .A(n45033), .B(n45037), .Z(n45180) );
  XNOR U45827 ( .A(n45028), .B(n45032), .Z(n45181) );
  XNOR U45828 ( .A(n45023), .B(n45027), .Z(n45182) );
  XNOR U45829 ( .A(n45018), .B(n45022), .Z(n45183) );
  XNOR U45830 ( .A(n45184), .B(n45017), .Z(n45018) );
  AND U45831 ( .A(a[0]), .B(b[29]), .Z(n45184) );
  XOR U45832 ( .A(n45185), .B(n45017), .Z(n45019) );
  XNOR U45833 ( .A(n45186), .B(n45187), .Z(n45017) );
  ANDN U45834 ( .B(n45188), .A(n45189), .Z(n45186) );
  AND U45835 ( .A(a[1]), .B(b[28]), .Z(n45185) );
  XOR U45836 ( .A(n45191), .B(n45192), .Z(n45022) );
  ANDN U45837 ( .B(n45193), .A(n45194), .Z(n45191) );
  AND U45838 ( .A(a[2]), .B(b[27]), .Z(n45190) );
  XOR U45839 ( .A(n45196), .B(n45197), .Z(n45027) );
  ANDN U45840 ( .B(n45198), .A(n45199), .Z(n45196) );
  AND U45841 ( .A(a[3]), .B(b[26]), .Z(n45195) );
  XOR U45842 ( .A(n45201), .B(n45202), .Z(n45032) );
  ANDN U45843 ( .B(n45203), .A(n45204), .Z(n45201) );
  AND U45844 ( .A(a[4]), .B(b[25]), .Z(n45200) );
  XOR U45845 ( .A(n45206), .B(n45207), .Z(n45037) );
  ANDN U45846 ( .B(n45208), .A(n45209), .Z(n45206) );
  AND U45847 ( .A(a[5]), .B(b[24]), .Z(n45205) );
  XOR U45848 ( .A(n45211), .B(n45212), .Z(n45042) );
  ANDN U45849 ( .B(n45213), .A(n45214), .Z(n45211) );
  AND U45850 ( .A(a[6]), .B(b[23]), .Z(n45210) );
  XOR U45851 ( .A(n45216), .B(n45217), .Z(n45047) );
  ANDN U45852 ( .B(n45218), .A(n45219), .Z(n45216) );
  AND U45853 ( .A(a[7]), .B(b[22]), .Z(n45215) );
  XOR U45854 ( .A(n45221), .B(n45222), .Z(n45052) );
  ANDN U45855 ( .B(n45223), .A(n45224), .Z(n45221) );
  AND U45856 ( .A(a[8]), .B(b[21]), .Z(n45220) );
  XOR U45857 ( .A(n45226), .B(n45227), .Z(n45057) );
  ANDN U45858 ( .B(n45228), .A(n45229), .Z(n45226) );
  AND U45859 ( .A(a[9]), .B(b[20]), .Z(n45225) );
  XOR U45860 ( .A(n45231), .B(n45232), .Z(n45062) );
  ANDN U45861 ( .B(n45233), .A(n45234), .Z(n45231) );
  AND U45862 ( .A(a[10]), .B(b[19]), .Z(n45230) );
  XOR U45863 ( .A(n45236), .B(n45237), .Z(n45067) );
  ANDN U45864 ( .B(n45238), .A(n45239), .Z(n45236) );
  AND U45865 ( .A(a[11]), .B(b[18]), .Z(n45235) );
  XOR U45866 ( .A(n45241), .B(n45242), .Z(n45072) );
  ANDN U45867 ( .B(n45243), .A(n45244), .Z(n45241) );
  AND U45868 ( .A(a[12]), .B(b[17]), .Z(n45240) );
  XOR U45869 ( .A(n45246), .B(n45247), .Z(n45077) );
  ANDN U45870 ( .B(n45248), .A(n45249), .Z(n45246) );
  AND U45871 ( .A(a[13]), .B(b[16]), .Z(n45245) );
  XOR U45872 ( .A(n45251), .B(n45252), .Z(n45082) );
  ANDN U45873 ( .B(n45253), .A(n45254), .Z(n45251) );
  AND U45874 ( .A(a[14]), .B(b[15]), .Z(n45250) );
  XOR U45875 ( .A(n45256), .B(n45257), .Z(n45087) );
  ANDN U45876 ( .B(n45258), .A(n45259), .Z(n45256) );
  AND U45877 ( .A(a[15]), .B(b[14]), .Z(n45255) );
  XOR U45878 ( .A(n45261), .B(n45262), .Z(n45092) );
  ANDN U45879 ( .B(n45263), .A(n45264), .Z(n45261) );
  AND U45880 ( .A(a[16]), .B(b[13]), .Z(n45260) );
  XOR U45881 ( .A(n45266), .B(n45267), .Z(n45097) );
  ANDN U45882 ( .B(n45268), .A(n45269), .Z(n45266) );
  AND U45883 ( .A(a[17]), .B(b[12]), .Z(n45265) );
  XOR U45884 ( .A(n45271), .B(n45272), .Z(n45102) );
  ANDN U45885 ( .B(n45273), .A(n45274), .Z(n45271) );
  AND U45886 ( .A(a[18]), .B(b[11]), .Z(n45270) );
  XOR U45887 ( .A(n45276), .B(n45277), .Z(n45107) );
  ANDN U45888 ( .B(n45278), .A(n45279), .Z(n45276) );
  AND U45889 ( .A(a[19]), .B(b[10]), .Z(n45275) );
  XOR U45890 ( .A(n45281), .B(n45282), .Z(n45112) );
  ANDN U45891 ( .B(n45283), .A(n45284), .Z(n45281) );
  AND U45892 ( .A(b[9]), .B(a[20]), .Z(n45280) );
  XOR U45893 ( .A(n45286), .B(n45287), .Z(n45117) );
  ANDN U45894 ( .B(n45288), .A(n45289), .Z(n45286) );
  AND U45895 ( .A(b[8]), .B(a[21]), .Z(n45285) );
  XOR U45896 ( .A(n45291), .B(n45292), .Z(n45122) );
  ANDN U45897 ( .B(n45293), .A(n45294), .Z(n45291) );
  AND U45898 ( .A(b[7]), .B(a[22]), .Z(n45290) );
  XOR U45899 ( .A(n45296), .B(n45297), .Z(n45127) );
  ANDN U45900 ( .B(n45298), .A(n45299), .Z(n45296) );
  AND U45901 ( .A(b[6]), .B(a[23]), .Z(n45295) );
  XOR U45902 ( .A(n45301), .B(n45302), .Z(n45132) );
  ANDN U45903 ( .B(n45303), .A(n45304), .Z(n45301) );
  AND U45904 ( .A(b[5]), .B(a[24]), .Z(n45300) );
  XOR U45905 ( .A(n45306), .B(n45307), .Z(n45137) );
  ANDN U45906 ( .B(n45308), .A(n45309), .Z(n45306) );
  AND U45907 ( .A(b[4]), .B(a[25]), .Z(n45305) );
  XOR U45908 ( .A(n45311), .B(n45312), .Z(n45142) );
  ANDN U45909 ( .B(n45154), .A(n45155), .Z(n45311) );
  AND U45910 ( .A(b[2]), .B(a[26]), .Z(n45313) );
  XNOR U45911 ( .A(n45308), .B(n45312), .Z(n45314) );
  XOR U45912 ( .A(n45315), .B(n45316), .Z(n45312) );
  OR U45913 ( .A(n45157), .B(n45158), .Z(n45316) );
  XNOR U45914 ( .A(n45318), .B(n45319), .Z(n45317) );
  XOR U45915 ( .A(n45318), .B(n45321), .Z(n45157) );
  NAND U45916 ( .A(b[1]), .B(a[26]), .Z(n45321) );
  IV U45917 ( .A(n45315), .Z(n45318) );
  NANDN U45918 ( .A(n163), .B(n164), .Z(n45315) );
  XOR U45919 ( .A(n45322), .B(n45323), .Z(n164) );
  NAND U45920 ( .A(a[26]), .B(b[0]), .Z(n163) );
  XNOR U45921 ( .A(n45303), .B(n45307), .Z(n45324) );
  XNOR U45922 ( .A(n45298), .B(n45302), .Z(n45325) );
  XNOR U45923 ( .A(n45293), .B(n45297), .Z(n45326) );
  XNOR U45924 ( .A(n45288), .B(n45292), .Z(n45327) );
  XNOR U45925 ( .A(n45283), .B(n45287), .Z(n45328) );
  XNOR U45926 ( .A(n45278), .B(n45282), .Z(n45329) );
  XNOR U45927 ( .A(n45273), .B(n45277), .Z(n45330) );
  XNOR U45928 ( .A(n45268), .B(n45272), .Z(n45331) );
  XNOR U45929 ( .A(n45263), .B(n45267), .Z(n45332) );
  XNOR U45930 ( .A(n45258), .B(n45262), .Z(n45333) );
  XNOR U45931 ( .A(n45253), .B(n45257), .Z(n45334) );
  XNOR U45932 ( .A(n45248), .B(n45252), .Z(n45335) );
  XNOR U45933 ( .A(n45243), .B(n45247), .Z(n45336) );
  XNOR U45934 ( .A(n45238), .B(n45242), .Z(n45337) );
  XNOR U45935 ( .A(n45233), .B(n45237), .Z(n45338) );
  XNOR U45936 ( .A(n45228), .B(n45232), .Z(n45339) );
  XNOR U45937 ( .A(n45223), .B(n45227), .Z(n45340) );
  XNOR U45938 ( .A(n45218), .B(n45222), .Z(n45341) );
  XNOR U45939 ( .A(n45213), .B(n45217), .Z(n45342) );
  XNOR U45940 ( .A(n45208), .B(n45212), .Z(n45343) );
  XNOR U45941 ( .A(n45203), .B(n45207), .Z(n45344) );
  XNOR U45942 ( .A(n45198), .B(n45202), .Z(n45345) );
  XNOR U45943 ( .A(n45193), .B(n45197), .Z(n45346) );
  XNOR U45944 ( .A(n45188), .B(n45192), .Z(n45347) );
  XOR U45945 ( .A(n45348), .B(n45187), .Z(n45188) );
  AND U45946 ( .A(a[0]), .B(b[28]), .Z(n45348) );
  XNOR U45947 ( .A(n45349), .B(n45187), .Z(n45189) );
  XNOR U45948 ( .A(n45350), .B(n45351), .Z(n45187) );
  ANDN U45949 ( .B(n45352), .A(n45353), .Z(n45350) );
  AND U45950 ( .A(a[1]), .B(b[27]), .Z(n45349) );
  XOR U45951 ( .A(n45355), .B(n45356), .Z(n45192) );
  ANDN U45952 ( .B(n45357), .A(n45358), .Z(n45355) );
  AND U45953 ( .A(a[2]), .B(b[26]), .Z(n45354) );
  XOR U45954 ( .A(n45360), .B(n45361), .Z(n45197) );
  ANDN U45955 ( .B(n45362), .A(n45363), .Z(n45360) );
  AND U45956 ( .A(a[3]), .B(b[25]), .Z(n45359) );
  XOR U45957 ( .A(n45365), .B(n45366), .Z(n45202) );
  ANDN U45958 ( .B(n45367), .A(n45368), .Z(n45365) );
  AND U45959 ( .A(a[4]), .B(b[24]), .Z(n45364) );
  XOR U45960 ( .A(n45370), .B(n45371), .Z(n45207) );
  ANDN U45961 ( .B(n45372), .A(n45373), .Z(n45370) );
  AND U45962 ( .A(a[5]), .B(b[23]), .Z(n45369) );
  XOR U45963 ( .A(n45375), .B(n45376), .Z(n45212) );
  ANDN U45964 ( .B(n45377), .A(n45378), .Z(n45375) );
  AND U45965 ( .A(a[6]), .B(b[22]), .Z(n45374) );
  XOR U45966 ( .A(n45380), .B(n45381), .Z(n45217) );
  ANDN U45967 ( .B(n45382), .A(n45383), .Z(n45380) );
  AND U45968 ( .A(a[7]), .B(b[21]), .Z(n45379) );
  XOR U45969 ( .A(n45385), .B(n45386), .Z(n45222) );
  ANDN U45970 ( .B(n45387), .A(n45388), .Z(n45385) );
  AND U45971 ( .A(a[8]), .B(b[20]), .Z(n45384) );
  XOR U45972 ( .A(n45390), .B(n45391), .Z(n45227) );
  ANDN U45973 ( .B(n45392), .A(n45393), .Z(n45390) );
  AND U45974 ( .A(a[9]), .B(b[19]), .Z(n45389) );
  XOR U45975 ( .A(n45395), .B(n45396), .Z(n45232) );
  ANDN U45976 ( .B(n45397), .A(n45398), .Z(n45395) );
  AND U45977 ( .A(a[10]), .B(b[18]), .Z(n45394) );
  XOR U45978 ( .A(n45400), .B(n45401), .Z(n45237) );
  ANDN U45979 ( .B(n45402), .A(n45403), .Z(n45400) );
  AND U45980 ( .A(a[11]), .B(b[17]), .Z(n45399) );
  XOR U45981 ( .A(n45405), .B(n45406), .Z(n45242) );
  ANDN U45982 ( .B(n45407), .A(n45408), .Z(n45405) );
  AND U45983 ( .A(a[12]), .B(b[16]), .Z(n45404) );
  XOR U45984 ( .A(n45410), .B(n45411), .Z(n45247) );
  ANDN U45985 ( .B(n45412), .A(n45413), .Z(n45410) );
  AND U45986 ( .A(a[13]), .B(b[15]), .Z(n45409) );
  XOR U45987 ( .A(n45415), .B(n45416), .Z(n45252) );
  ANDN U45988 ( .B(n45417), .A(n45418), .Z(n45415) );
  AND U45989 ( .A(a[14]), .B(b[14]), .Z(n45414) );
  XOR U45990 ( .A(n45420), .B(n45421), .Z(n45257) );
  ANDN U45991 ( .B(n45422), .A(n45423), .Z(n45420) );
  AND U45992 ( .A(a[15]), .B(b[13]), .Z(n45419) );
  XOR U45993 ( .A(n45425), .B(n45426), .Z(n45262) );
  ANDN U45994 ( .B(n45427), .A(n45428), .Z(n45425) );
  AND U45995 ( .A(a[16]), .B(b[12]), .Z(n45424) );
  XOR U45996 ( .A(n45430), .B(n45431), .Z(n45267) );
  ANDN U45997 ( .B(n45432), .A(n45433), .Z(n45430) );
  AND U45998 ( .A(a[17]), .B(b[11]), .Z(n45429) );
  XOR U45999 ( .A(n45435), .B(n45436), .Z(n45272) );
  ANDN U46000 ( .B(n45437), .A(n45438), .Z(n45435) );
  AND U46001 ( .A(a[18]), .B(b[10]), .Z(n45434) );
  XOR U46002 ( .A(n45440), .B(n45441), .Z(n45277) );
  ANDN U46003 ( .B(n45442), .A(n45443), .Z(n45440) );
  AND U46004 ( .A(b[9]), .B(a[19]), .Z(n45439) );
  XOR U46005 ( .A(n45445), .B(n45446), .Z(n45282) );
  ANDN U46006 ( .B(n45447), .A(n45448), .Z(n45445) );
  AND U46007 ( .A(b[8]), .B(a[20]), .Z(n45444) );
  XOR U46008 ( .A(n45450), .B(n45451), .Z(n45287) );
  ANDN U46009 ( .B(n45452), .A(n45453), .Z(n45450) );
  AND U46010 ( .A(b[7]), .B(a[21]), .Z(n45449) );
  XOR U46011 ( .A(n45455), .B(n45456), .Z(n45292) );
  ANDN U46012 ( .B(n45457), .A(n45458), .Z(n45455) );
  AND U46013 ( .A(b[6]), .B(a[22]), .Z(n45454) );
  XOR U46014 ( .A(n45460), .B(n45461), .Z(n45297) );
  ANDN U46015 ( .B(n45462), .A(n45463), .Z(n45460) );
  AND U46016 ( .A(b[5]), .B(a[23]), .Z(n45459) );
  XOR U46017 ( .A(n45465), .B(n45466), .Z(n45302) );
  ANDN U46018 ( .B(n45467), .A(n45468), .Z(n45465) );
  AND U46019 ( .A(b[4]), .B(a[24]), .Z(n45464) );
  XOR U46020 ( .A(n45470), .B(n45471), .Z(n45307) );
  ANDN U46021 ( .B(n45319), .A(n45320), .Z(n45470) );
  AND U46022 ( .A(b[2]), .B(a[25]), .Z(n45472) );
  XNOR U46023 ( .A(n45467), .B(n45471), .Z(n45473) );
  XOR U46024 ( .A(n45474), .B(n45475), .Z(n45471) );
  OR U46025 ( .A(n45322), .B(n45323), .Z(n45475) );
  XNOR U46026 ( .A(n45477), .B(n45478), .Z(n45476) );
  XOR U46027 ( .A(n45477), .B(n45480), .Z(n45322) );
  NAND U46028 ( .A(b[1]), .B(a[25]), .Z(n45480) );
  IV U46029 ( .A(n45474), .Z(n45477) );
  NANDN U46030 ( .A(n165), .B(n166), .Z(n45474) );
  XOR U46031 ( .A(n45481), .B(n45482), .Z(n166) );
  NAND U46032 ( .A(a[25]), .B(b[0]), .Z(n165) );
  XNOR U46033 ( .A(n45462), .B(n45466), .Z(n45483) );
  XNOR U46034 ( .A(n45457), .B(n45461), .Z(n45484) );
  XNOR U46035 ( .A(n45452), .B(n45456), .Z(n45485) );
  XNOR U46036 ( .A(n45447), .B(n45451), .Z(n45486) );
  XNOR U46037 ( .A(n45442), .B(n45446), .Z(n45487) );
  XNOR U46038 ( .A(n45437), .B(n45441), .Z(n45488) );
  XNOR U46039 ( .A(n45432), .B(n45436), .Z(n45489) );
  XNOR U46040 ( .A(n45427), .B(n45431), .Z(n45490) );
  XNOR U46041 ( .A(n45422), .B(n45426), .Z(n45491) );
  XNOR U46042 ( .A(n45417), .B(n45421), .Z(n45492) );
  XNOR U46043 ( .A(n45412), .B(n45416), .Z(n45493) );
  XNOR U46044 ( .A(n45407), .B(n45411), .Z(n45494) );
  XNOR U46045 ( .A(n45402), .B(n45406), .Z(n45495) );
  XNOR U46046 ( .A(n45397), .B(n45401), .Z(n45496) );
  XNOR U46047 ( .A(n45392), .B(n45396), .Z(n45497) );
  XNOR U46048 ( .A(n45387), .B(n45391), .Z(n45498) );
  XNOR U46049 ( .A(n45382), .B(n45386), .Z(n45499) );
  XNOR U46050 ( .A(n45377), .B(n45381), .Z(n45500) );
  XNOR U46051 ( .A(n45372), .B(n45376), .Z(n45501) );
  XNOR U46052 ( .A(n45367), .B(n45371), .Z(n45502) );
  XNOR U46053 ( .A(n45362), .B(n45366), .Z(n45503) );
  XNOR U46054 ( .A(n45357), .B(n45361), .Z(n45504) );
  XNOR U46055 ( .A(n45352), .B(n45356), .Z(n45505) );
  XNOR U46056 ( .A(n45506), .B(n45351), .Z(n45352) );
  AND U46057 ( .A(a[0]), .B(b[27]), .Z(n45506) );
  XOR U46058 ( .A(n45507), .B(n45351), .Z(n45353) );
  XNOR U46059 ( .A(n45508), .B(n45509), .Z(n45351) );
  ANDN U46060 ( .B(n45510), .A(n45511), .Z(n45508) );
  AND U46061 ( .A(a[1]), .B(b[26]), .Z(n45507) );
  XOR U46062 ( .A(n45513), .B(n45514), .Z(n45356) );
  ANDN U46063 ( .B(n45515), .A(n45516), .Z(n45513) );
  AND U46064 ( .A(a[2]), .B(b[25]), .Z(n45512) );
  XOR U46065 ( .A(n45518), .B(n45519), .Z(n45361) );
  ANDN U46066 ( .B(n45520), .A(n45521), .Z(n45518) );
  AND U46067 ( .A(a[3]), .B(b[24]), .Z(n45517) );
  XOR U46068 ( .A(n45523), .B(n45524), .Z(n45366) );
  ANDN U46069 ( .B(n45525), .A(n45526), .Z(n45523) );
  AND U46070 ( .A(a[4]), .B(b[23]), .Z(n45522) );
  XOR U46071 ( .A(n45528), .B(n45529), .Z(n45371) );
  ANDN U46072 ( .B(n45530), .A(n45531), .Z(n45528) );
  AND U46073 ( .A(a[5]), .B(b[22]), .Z(n45527) );
  XOR U46074 ( .A(n45533), .B(n45534), .Z(n45376) );
  ANDN U46075 ( .B(n45535), .A(n45536), .Z(n45533) );
  AND U46076 ( .A(a[6]), .B(b[21]), .Z(n45532) );
  XOR U46077 ( .A(n45538), .B(n45539), .Z(n45381) );
  ANDN U46078 ( .B(n45540), .A(n45541), .Z(n45538) );
  AND U46079 ( .A(a[7]), .B(b[20]), .Z(n45537) );
  XOR U46080 ( .A(n45543), .B(n45544), .Z(n45386) );
  ANDN U46081 ( .B(n45545), .A(n45546), .Z(n45543) );
  AND U46082 ( .A(a[8]), .B(b[19]), .Z(n45542) );
  XOR U46083 ( .A(n45548), .B(n45549), .Z(n45391) );
  ANDN U46084 ( .B(n45550), .A(n45551), .Z(n45548) );
  AND U46085 ( .A(a[9]), .B(b[18]), .Z(n45547) );
  XOR U46086 ( .A(n45553), .B(n45554), .Z(n45396) );
  ANDN U46087 ( .B(n45555), .A(n45556), .Z(n45553) );
  AND U46088 ( .A(a[10]), .B(b[17]), .Z(n45552) );
  XOR U46089 ( .A(n45558), .B(n45559), .Z(n45401) );
  ANDN U46090 ( .B(n45560), .A(n45561), .Z(n45558) );
  AND U46091 ( .A(a[11]), .B(b[16]), .Z(n45557) );
  XOR U46092 ( .A(n45563), .B(n45564), .Z(n45406) );
  ANDN U46093 ( .B(n45565), .A(n45566), .Z(n45563) );
  AND U46094 ( .A(a[12]), .B(b[15]), .Z(n45562) );
  XOR U46095 ( .A(n45568), .B(n45569), .Z(n45411) );
  ANDN U46096 ( .B(n45570), .A(n45571), .Z(n45568) );
  AND U46097 ( .A(a[13]), .B(b[14]), .Z(n45567) );
  XOR U46098 ( .A(n45573), .B(n45574), .Z(n45416) );
  ANDN U46099 ( .B(n45575), .A(n45576), .Z(n45573) );
  AND U46100 ( .A(a[14]), .B(b[13]), .Z(n45572) );
  XOR U46101 ( .A(n45578), .B(n45579), .Z(n45421) );
  ANDN U46102 ( .B(n45580), .A(n45581), .Z(n45578) );
  AND U46103 ( .A(a[15]), .B(b[12]), .Z(n45577) );
  XOR U46104 ( .A(n45583), .B(n45584), .Z(n45426) );
  ANDN U46105 ( .B(n45585), .A(n45586), .Z(n45583) );
  AND U46106 ( .A(a[16]), .B(b[11]), .Z(n45582) );
  XOR U46107 ( .A(n45588), .B(n45589), .Z(n45431) );
  ANDN U46108 ( .B(n45590), .A(n45591), .Z(n45588) );
  AND U46109 ( .A(a[17]), .B(b[10]), .Z(n45587) );
  XOR U46110 ( .A(n45593), .B(n45594), .Z(n45436) );
  ANDN U46111 ( .B(n45595), .A(n45596), .Z(n45593) );
  AND U46112 ( .A(b[9]), .B(a[18]), .Z(n45592) );
  XOR U46113 ( .A(n45598), .B(n45599), .Z(n45441) );
  ANDN U46114 ( .B(n45600), .A(n45601), .Z(n45598) );
  AND U46115 ( .A(b[8]), .B(a[19]), .Z(n45597) );
  XOR U46116 ( .A(n45603), .B(n45604), .Z(n45446) );
  ANDN U46117 ( .B(n45605), .A(n45606), .Z(n45603) );
  AND U46118 ( .A(b[7]), .B(a[20]), .Z(n45602) );
  XOR U46119 ( .A(n45608), .B(n45609), .Z(n45451) );
  ANDN U46120 ( .B(n45610), .A(n45611), .Z(n45608) );
  AND U46121 ( .A(b[6]), .B(a[21]), .Z(n45607) );
  XOR U46122 ( .A(n45613), .B(n45614), .Z(n45456) );
  ANDN U46123 ( .B(n45615), .A(n45616), .Z(n45613) );
  AND U46124 ( .A(b[5]), .B(a[22]), .Z(n45612) );
  XOR U46125 ( .A(n45618), .B(n45619), .Z(n45461) );
  ANDN U46126 ( .B(n45620), .A(n45621), .Z(n45618) );
  AND U46127 ( .A(b[4]), .B(a[23]), .Z(n45617) );
  XOR U46128 ( .A(n45623), .B(n45624), .Z(n45466) );
  ANDN U46129 ( .B(n45478), .A(n45479), .Z(n45623) );
  AND U46130 ( .A(b[2]), .B(a[24]), .Z(n45625) );
  XNOR U46131 ( .A(n45620), .B(n45624), .Z(n45626) );
  XOR U46132 ( .A(n45627), .B(n45628), .Z(n45624) );
  OR U46133 ( .A(n45481), .B(n45482), .Z(n45628) );
  XNOR U46134 ( .A(n45630), .B(n45631), .Z(n45629) );
  XOR U46135 ( .A(n45630), .B(n45633), .Z(n45481) );
  NAND U46136 ( .A(b[1]), .B(a[24]), .Z(n45633) );
  IV U46137 ( .A(n45627), .Z(n45630) );
  NANDN U46138 ( .A(n167), .B(n168), .Z(n45627) );
  XOR U46139 ( .A(n45634), .B(n45635), .Z(n168) );
  NAND U46140 ( .A(a[24]), .B(b[0]), .Z(n167) );
  XNOR U46141 ( .A(n45615), .B(n45619), .Z(n45636) );
  XNOR U46142 ( .A(n45610), .B(n45614), .Z(n45637) );
  XNOR U46143 ( .A(n45605), .B(n45609), .Z(n45638) );
  XNOR U46144 ( .A(n45600), .B(n45604), .Z(n45639) );
  XNOR U46145 ( .A(n45595), .B(n45599), .Z(n45640) );
  XNOR U46146 ( .A(n45590), .B(n45594), .Z(n45641) );
  XNOR U46147 ( .A(n45585), .B(n45589), .Z(n45642) );
  XNOR U46148 ( .A(n45580), .B(n45584), .Z(n45643) );
  XNOR U46149 ( .A(n45575), .B(n45579), .Z(n45644) );
  XNOR U46150 ( .A(n45570), .B(n45574), .Z(n45645) );
  XNOR U46151 ( .A(n45565), .B(n45569), .Z(n45646) );
  XNOR U46152 ( .A(n45560), .B(n45564), .Z(n45647) );
  XNOR U46153 ( .A(n45555), .B(n45559), .Z(n45648) );
  XNOR U46154 ( .A(n45550), .B(n45554), .Z(n45649) );
  XNOR U46155 ( .A(n45545), .B(n45549), .Z(n45650) );
  XNOR U46156 ( .A(n45540), .B(n45544), .Z(n45651) );
  XNOR U46157 ( .A(n45535), .B(n45539), .Z(n45652) );
  XNOR U46158 ( .A(n45530), .B(n45534), .Z(n45653) );
  XNOR U46159 ( .A(n45525), .B(n45529), .Z(n45654) );
  XNOR U46160 ( .A(n45520), .B(n45524), .Z(n45655) );
  XNOR U46161 ( .A(n45515), .B(n45519), .Z(n45656) );
  XNOR U46162 ( .A(n45510), .B(n45514), .Z(n45657) );
  XOR U46163 ( .A(n45658), .B(n45509), .Z(n45510) );
  AND U46164 ( .A(a[0]), .B(b[26]), .Z(n45658) );
  XNOR U46165 ( .A(n45659), .B(n45509), .Z(n45511) );
  XNOR U46166 ( .A(n45660), .B(n45661), .Z(n45509) );
  ANDN U46167 ( .B(n45662), .A(n45663), .Z(n45660) );
  AND U46168 ( .A(a[1]), .B(b[25]), .Z(n45659) );
  XOR U46169 ( .A(n45665), .B(n45666), .Z(n45514) );
  ANDN U46170 ( .B(n45667), .A(n45668), .Z(n45665) );
  AND U46171 ( .A(a[2]), .B(b[24]), .Z(n45664) );
  XOR U46172 ( .A(n45670), .B(n45671), .Z(n45519) );
  ANDN U46173 ( .B(n45672), .A(n45673), .Z(n45670) );
  AND U46174 ( .A(a[3]), .B(b[23]), .Z(n45669) );
  XOR U46175 ( .A(n45675), .B(n45676), .Z(n45524) );
  ANDN U46176 ( .B(n45677), .A(n45678), .Z(n45675) );
  AND U46177 ( .A(a[4]), .B(b[22]), .Z(n45674) );
  XOR U46178 ( .A(n45680), .B(n45681), .Z(n45529) );
  ANDN U46179 ( .B(n45682), .A(n45683), .Z(n45680) );
  AND U46180 ( .A(a[5]), .B(b[21]), .Z(n45679) );
  XOR U46181 ( .A(n45685), .B(n45686), .Z(n45534) );
  ANDN U46182 ( .B(n45687), .A(n45688), .Z(n45685) );
  AND U46183 ( .A(a[6]), .B(b[20]), .Z(n45684) );
  XOR U46184 ( .A(n45690), .B(n45691), .Z(n45539) );
  ANDN U46185 ( .B(n45692), .A(n45693), .Z(n45690) );
  AND U46186 ( .A(a[7]), .B(b[19]), .Z(n45689) );
  XOR U46187 ( .A(n45695), .B(n45696), .Z(n45544) );
  ANDN U46188 ( .B(n45697), .A(n45698), .Z(n45695) );
  AND U46189 ( .A(a[8]), .B(b[18]), .Z(n45694) );
  XOR U46190 ( .A(n45700), .B(n45701), .Z(n45549) );
  ANDN U46191 ( .B(n45702), .A(n45703), .Z(n45700) );
  AND U46192 ( .A(a[9]), .B(b[17]), .Z(n45699) );
  XOR U46193 ( .A(n45705), .B(n45706), .Z(n45554) );
  ANDN U46194 ( .B(n45707), .A(n45708), .Z(n45705) );
  AND U46195 ( .A(a[10]), .B(b[16]), .Z(n45704) );
  XOR U46196 ( .A(n45710), .B(n45711), .Z(n45559) );
  ANDN U46197 ( .B(n45712), .A(n45713), .Z(n45710) );
  AND U46198 ( .A(a[11]), .B(b[15]), .Z(n45709) );
  XOR U46199 ( .A(n45715), .B(n45716), .Z(n45564) );
  ANDN U46200 ( .B(n45717), .A(n45718), .Z(n45715) );
  AND U46201 ( .A(a[12]), .B(b[14]), .Z(n45714) );
  XOR U46202 ( .A(n45720), .B(n45721), .Z(n45569) );
  ANDN U46203 ( .B(n45722), .A(n45723), .Z(n45720) );
  AND U46204 ( .A(a[13]), .B(b[13]), .Z(n45719) );
  XOR U46205 ( .A(n45725), .B(n45726), .Z(n45574) );
  ANDN U46206 ( .B(n45727), .A(n45728), .Z(n45725) );
  AND U46207 ( .A(a[14]), .B(b[12]), .Z(n45724) );
  XOR U46208 ( .A(n45730), .B(n45731), .Z(n45579) );
  ANDN U46209 ( .B(n45732), .A(n45733), .Z(n45730) );
  AND U46210 ( .A(a[15]), .B(b[11]), .Z(n45729) );
  XOR U46211 ( .A(n45735), .B(n45736), .Z(n45584) );
  ANDN U46212 ( .B(n45737), .A(n45738), .Z(n45735) );
  AND U46213 ( .A(a[16]), .B(b[10]), .Z(n45734) );
  XOR U46214 ( .A(n45740), .B(n45741), .Z(n45589) );
  ANDN U46215 ( .B(n45742), .A(n45743), .Z(n45740) );
  AND U46216 ( .A(b[9]), .B(a[17]), .Z(n45739) );
  XOR U46217 ( .A(n45745), .B(n45746), .Z(n45594) );
  ANDN U46218 ( .B(n45747), .A(n45748), .Z(n45745) );
  AND U46219 ( .A(b[8]), .B(a[18]), .Z(n45744) );
  XOR U46220 ( .A(n45750), .B(n45751), .Z(n45599) );
  ANDN U46221 ( .B(n45752), .A(n45753), .Z(n45750) );
  AND U46222 ( .A(b[7]), .B(a[19]), .Z(n45749) );
  XOR U46223 ( .A(n45755), .B(n45756), .Z(n45604) );
  ANDN U46224 ( .B(n45757), .A(n45758), .Z(n45755) );
  AND U46225 ( .A(b[6]), .B(a[20]), .Z(n45754) );
  XOR U46226 ( .A(n45760), .B(n45761), .Z(n45609) );
  ANDN U46227 ( .B(n45762), .A(n45763), .Z(n45760) );
  AND U46228 ( .A(b[5]), .B(a[21]), .Z(n45759) );
  XOR U46229 ( .A(n45765), .B(n45766), .Z(n45614) );
  ANDN U46230 ( .B(n45767), .A(n45768), .Z(n45765) );
  AND U46231 ( .A(b[4]), .B(a[22]), .Z(n45764) );
  XOR U46232 ( .A(n45770), .B(n45771), .Z(n45619) );
  ANDN U46233 ( .B(n45631), .A(n45632), .Z(n45770) );
  AND U46234 ( .A(b[2]), .B(a[23]), .Z(n45772) );
  XNOR U46235 ( .A(n45767), .B(n45771), .Z(n45773) );
  XOR U46236 ( .A(n45774), .B(n45775), .Z(n45771) );
  OR U46237 ( .A(n45634), .B(n45635), .Z(n45775) );
  XNOR U46238 ( .A(n45777), .B(n45778), .Z(n45776) );
  XOR U46239 ( .A(n45777), .B(n45780), .Z(n45634) );
  NAND U46240 ( .A(b[1]), .B(a[23]), .Z(n45780) );
  IV U46241 ( .A(n45774), .Z(n45777) );
  NANDN U46242 ( .A(n169), .B(n170), .Z(n45774) );
  XOR U46243 ( .A(n45781), .B(n45782), .Z(n170) );
  NAND U46244 ( .A(a[23]), .B(b[0]), .Z(n169) );
  XNOR U46245 ( .A(n45762), .B(n45766), .Z(n45783) );
  XNOR U46246 ( .A(n45757), .B(n45761), .Z(n45784) );
  XNOR U46247 ( .A(n45752), .B(n45756), .Z(n45785) );
  XNOR U46248 ( .A(n45747), .B(n45751), .Z(n45786) );
  XNOR U46249 ( .A(n45742), .B(n45746), .Z(n45787) );
  XNOR U46250 ( .A(n45737), .B(n45741), .Z(n45788) );
  XNOR U46251 ( .A(n45732), .B(n45736), .Z(n45789) );
  XNOR U46252 ( .A(n45727), .B(n45731), .Z(n45790) );
  XNOR U46253 ( .A(n45722), .B(n45726), .Z(n45791) );
  XNOR U46254 ( .A(n45717), .B(n45721), .Z(n45792) );
  XNOR U46255 ( .A(n45712), .B(n45716), .Z(n45793) );
  XNOR U46256 ( .A(n45707), .B(n45711), .Z(n45794) );
  XNOR U46257 ( .A(n45702), .B(n45706), .Z(n45795) );
  XNOR U46258 ( .A(n45697), .B(n45701), .Z(n45796) );
  XNOR U46259 ( .A(n45692), .B(n45696), .Z(n45797) );
  XNOR U46260 ( .A(n45687), .B(n45691), .Z(n45798) );
  XNOR U46261 ( .A(n45682), .B(n45686), .Z(n45799) );
  XNOR U46262 ( .A(n45677), .B(n45681), .Z(n45800) );
  XNOR U46263 ( .A(n45672), .B(n45676), .Z(n45801) );
  XNOR U46264 ( .A(n45667), .B(n45671), .Z(n45802) );
  XNOR U46265 ( .A(n45662), .B(n45666), .Z(n45803) );
  XNOR U46266 ( .A(n45804), .B(n45661), .Z(n45662) );
  AND U46267 ( .A(a[0]), .B(b[25]), .Z(n45804) );
  XOR U46268 ( .A(n45805), .B(n45661), .Z(n45663) );
  XNOR U46269 ( .A(n45806), .B(n45807), .Z(n45661) );
  ANDN U46270 ( .B(n45808), .A(n45809), .Z(n45806) );
  AND U46271 ( .A(a[1]), .B(b[24]), .Z(n45805) );
  XOR U46272 ( .A(n45811), .B(n45812), .Z(n45666) );
  ANDN U46273 ( .B(n45813), .A(n45814), .Z(n45811) );
  AND U46274 ( .A(a[2]), .B(b[23]), .Z(n45810) );
  XOR U46275 ( .A(n45816), .B(n45817), .Z(n45671) );
  ANDN U46276 ( .B(n45818), .A(n45819), .Z(n45816) );
  AND U46277 ( .A(a[3]), .B(b[22]), .Z(n45815) );
  XOR U46278 ( .A(n45821), .B(n45822), .Z(n45676) );
  ANDN U46279 ( .B(n45823), .A(n45824), .Z(n45821) );
  AND U46280 ( .A(a[4]), .B(b[21]), .Z(n45820) );
  XOR U46281 ( .A(n45826), .B(n45827), .Z(n45681) );
  ANDN U46282 ( .B(n45828), .A(n45829), .Z(n45826) );
  AND U46283 ( .A(a[5]), .B(b[20]), .Z(n45825) );
  XOR U46284 ( .A(n45831), .B(n45832), .Z(n45686) );
  ANDN U46285 ( .B(n45833), .A(n45834), .Z(n45831) );
  AND U46286 ( .A(a[6]), .B(b[19]), .Z(n45830) );
  XOR U46287 ( .A(n45836), .B(n45837), .Z(n45691) );
  ANDN U46288 ( .B(n45838), .A(n45839), .Z(n45836) );
  AND U46289 ( .A(a[7]), .B(b[18]), .Z(n45835) );
  XOR U46290 ( .A(n45841), .B(n45842), .Z(n45696) );
  ANDN U46291 ( .B(n45843), .A(n45844), .Z(n45841) );
  AND U46292 ( .A(a[8]), .B(b[17]), .Z(n45840) );
  XOR U46293 ( .A(n45846), .B(n45847), .Z(n45701) );
  ANDN U46294 ( .B(n45848), .A(n45849), .Z(n45846) );
  AND U46295 ( .A(a[9]), .B(b[16]), .Z(n45845) );
  XOR U46296 ( .A(n45851), .B(n45852), .Z(n45706) );
  ANDN U46297 ( .B(n45853), .A(n45854), .Z(n45851) );
  AND U46298 ( .A(a[10]), .B(b[15]), .Z(n45850) );
  XOR U46299 ( .A(n45856), .B(n45857), .Z(n45711) );
  ANDN U46300 ( .B(n45858), .A(n45859), .Z(n45856) );
  AND U46301 ( .A(a[11]), .B(b[14]), .Z(n45855) );
  XOR U46302 ( .A(n45861), .B(n45862), .Z(n45716) );
  ANDN U46303 ( .B(n45863), .A(n45864), .Z(n45861) );
  AND U46304 ( .A(a[12]), .B(b[13]), .Z(n45860) );
  XOR U46305 ( .A(n45866), .B(n45867), .Z(n45721) );
  ANDN U46306 ( .B(n45868), .A(n45869), .Z(n45866) );
  AND U46307 ( .A(a[13]), .B(b[12]), .Z(n45865) );
  XOR U46308 ( .A(n45871), .B(n45872), .Z(n45726) );
  ANDN U46309 ( .B(n45873), .A(n45874), .Z(n45871) );
  AND U46310 ( .A(a[14]), .B(b[11]), .Z(n45870) );
  XOR U46311 ( .A(n45876), .B(n45877), .Z(n45731) );
  ANDN U46312 ( .B(n45878), .A(n45879), .Z(n45876) );
  AND U46313 ( .A(a[15]), .B(b[10]), .Z(n45875) );
  XOR U46314 ( .A(n45881), .B(n45882), .Z(n45736) );
  ANDN U46315 ( .B(n45883), .A(n45884), .Z(n45881) );
  AND U46316 ( .A(b[9]), .B(a[16]), .Z(n45880) );
  XOR U46317 ( .A(n45886), .B(n45887), .Z(n45741) );
  ANDN U46318 ( .B(n45888), .A(n45889), .Z(n45886) );
  AND U46319 ( .A(b[8]), .B(a[17]), .Z(n45885) );
  XOR U46320 ( .A(n45891), .B(n45892), .Z(n45746) );
  ANDN U46321 ( .B(n45893), .A(n45894), .Z(n45891) );
  AND U46322 ( .A(b[7]), .B(a[18]), .Z(n45890) );
  XOR U46323 ( .A(n45896), .B(n45897), .Z(n45751) );
  ANDN U46324 ( .B(n45898), .A(n45899), .Z(n45896) );
  AND U46325 ( .A(b[6]), .B(a[19]), .Z(n45895) );
  XOR U46326 ( .A(n45901), .B(n45902), .Z(n45756) );
  ANDN U46327 ( .B(n45903), .A(n45904), .Z(n45901) );
  AND U46328 ( .A(b[5]), .B(a[20]), .Z(n45900) );
  XOR U46329 ( .A(n45906), .B(n45907), .Z(n45761) );
  ANDN U46330 ( .B(n45908), .A(n45909), .Z(n45906) );
  AND U46331 ( .A(b[4]), .B(a[21]), .Z(n45905) );
  XOR U46332 ( .A(n45911), .B(n45912), .Z(n45766) );
  ANDN U46333 ( .B(n45778), .A(n45779), .Z(n45911) );
  AND U46334 ( .A(b[2]), .B(a[22]), .Z(n45913) );
  XNOR U46335 ( .A(n45908), .B(n45912), .Z(n45914) );
  XOR U46336 ( .A(n45915), .B(n45916), .Z(n45912) );
  OR U46337 ( .A(n45781), .B(n45782), .Z(n45916) );
  XNOR U46338 ( .A(n45918), .B(n45919), .Z(n45917) );
  XOR U46339 ( .A(n45918), .B(n45921), .Z(n45781) );
  NAND U46340 ( .A(b[1]), .B(a[22]), .Z(n45921) );
  IV U46341 ( .A(n45915), .Z(n45918) );
  NANDN U46342 ( .A(n171), .B(n172), .Z(n45915) );
  XOR U46343 ( .A(n45922), .B(n45923), .Z(n172) );
  NAND U46344 ( .A(a[22]), .B(b[0]), .Z(n171) );
  XNOR U46345 ( .A(n45903), .B(n45907), .Z(n45924) );
  XNOR U46346 ( .A(n45898), .B(n45902), .Z(n45925) );
  XNOR U46347 ( .A(n45893), .B(n45897), .Z(n45926) );
  XNOR U46348 ( .A(n45888), .B(n45892), .Z(n45927) );
  XNOR U46349 ( .A(n45883), .B(n45887), .Z(n45928) );
  XNOR U46350 ( .A(n45878), .B(n45882), .Z(n45929) );
  XNOR U46351 ( .A(n45873), .B(n45877), .Z(n45930) );
  XNOR U46352 ( .A(n45868), .B(n45872), .Z(n45931) );
  XNOR U46353 ( .A(n45863), .B(n45867), .Z(n45932) );
  XNOR U46354 ( .A(n45858), .B(n45862), .Z(n45933) );
  XNOR U46355 ( .A(n45853), .B(n45857), .Z(n45934) );
  XNOR U46356 ( .A(n45848), .B(n45852), .Z(n45935) );
  XNOR U46357 ( .A(n45843), .B(n45847), .Z(n45936) );
  XNOR U46358 ( .A(n45838), .B(n45842), .Z(n45937) );
  XNOR U46359 ( .A(n45833), .B(n45837), .Z(n45938) );
  XNOR U46360 ( .A(n45828), .B(n45832), .Z(n45939) );
  XNOR U46361 ( .A(n45823), .B(n45827), .Z(n45940) );
  XNOR U46362 ( .A(n45818), .B(n45822), .Z(n45941) );
  XNOR U46363 ( .A(n45813), .B(n45817), .Z(n45942) );
  XNOR U46364 ( .A(n45808), .B(n45812), .Z(n45943) );
  XOR U46365 ( .A(n45944), .B(n45807), .Z(n45808) );
  AND U46366 ( .A(a[0]), .B(b[24]), .Z(n45944) );
  XNOR U46367 ( .A(n45945), .B(n45807), .Z(n45809) );
  XNOR U46368 ( .A(n45946), .B(n45947), .Z(n45807) );
  ANDN U46369 ( .B(n45948), .A(n45949), .Z(n45946) );
  AND U46370 ( .A(a[1]), .B(b[23]), .Z(n45945) );
  XOR U46371 ( .A(n45951), .B(n45952), .Z(n45812) );
  ANDN U46372 ( .B(n45953), .A(n45954), .Z(n45951) );
  AND U46373 ( .A(a[2]), .B(b[22]), .Z(n45950) );
  XOR U46374 ( .A(n45956), .B(n45957), .Z(n45817) );
  ANDN U46375 ( .B(n45958), .A(n45959), .Z(n45956) );
  AND U46376 ( .A(a[3]), .B(b[21]), .Z(n45955) );
  XOR U46377 ( .A(n45961), .B(n45962), .Z(n45822) );
  ANDN U46378 ( .B(n45963), .A(n45964), .Z(n45961) );
  AND U46379 ( .A(a[4]), .B(b[20]), .Z(n45960) );
  XOR U46380 ( .A(n45966), .B(n45967), .Z(n45827) );
  ANDN U46381 ( .B(n45968), .A(n45969), .Z(n45966) );
  AND U46382 ( .A(a[5]), .B(b[19]), .Z(n45965) );
  XOR U46383 ( .A(n45971), .B(n45972), .Z(n45832) );
  ANDN U46384 ( .B(n45973), .A(n45974), .Z(n45971) );
  AND U46385 ( .A(a[6]), .B(b[18]), .Z(n45970) );
  XOR U46386 ( .A(n45976), .B(n45977), .Z(n45837) );
  ANDN U46387 ( .B(n45978), .A(n45979), .Z(n45976) );
  AND U46388 ( .A(a[7]), .B(b[17]), .Z(n45975) );
  XOR U46389 ( .A(n45981), .B(n45982), .Z(n45842) );
  ANDN U46390 ( .B(n45983), .A(n45984), .Z(n45981) );
  AND U46391 ( .A(a[8]), .B(b[16]), .Z(n45980) );
  XOR U46392 ( .A(n45986), .B(n45987), .Z(n45847) );
  ANDN U46393 ( .B(n45988), .A(n45989), .Z(n45986) );
  AND U46394 ( .A(a[9]), .B(b[15]), .Z(n45985) );
  XOR U46395 ( .A(n45991), .B(n45992), .Z(n45852) );
  ANDN U46396 ( .B(n45993), .A(n45994), .Z(n45991) );
  AND U46397 ( .A(a[10]), .B(b[14]), .Z(n45990) );
  XOR U46398 ( .A(n45996), .B(n45997), .Z(n45857) );
  ANDN U46399 ( .B(n45998), .A(n45999), .Z(n45996) );
  AND U46400 ( .A(a[11]), .B(b[13]), .Z(n45995) );
  XOR U46401 ( .A(n46001), .B(n46002), .Z(n45862) );
  ANDN U46402 ( .B(n46003), .A(n46004), .Z(n46001) );
  AND U46403 ( .A(a[12]), .B(b[12]), .Z(n46000) );
  XOR U46404 ( .A(n46006), .B(n46007), .Z(n45867) );
  ANDN U46405 ( .B(n46008), .A(n46009), .Z(n46006) );
  AND U46406 ( .A(a[13]), .B(b[11]), .Z(n46005) );
  XOR U46407 ( .A(n46011), .B(n46012), .Z(n45872) );
  ANDN U46408 ( .B(n46013), .A(n46014), .Z(n46011) );
  AND U46409 ( .A(a[14]), .B(b[10]), .Z(n46010) );
  XOR U46410 ( .A(n46016), .B(n46017), .Z(n45877) );
  ANDN U46411 ( .B(n46018), .A(n46019), .Z(n46016) );
  AND U46412 ( .A(b[9]), .B(a[15]), .Z(n46015) );
  XOR U46413 ( .A(n46021), .B(n46022), .Z(n45882) );
  ANDN U46414 ( .B(n46023), .A(n46024), .Z(n46021) );
  AND U46415 ( .A(b[8]), .B(a[16]), .Z(n46020) );
  XOR U46416 ( .A(n46026), .B(n46027), .Z(n45887) );
  ANDN U46417 ( .B(n46028), .A(n46029), .Z(n46026) );
  AND U46418 ( .A(b[7]), .B(a[17]), .Z(n46025) );
  XOR U46419 ( .A(n46031), .B(n46032), .Z(n45892) );
  ANDN U46420 ( .B(n46033), .A(n46034), .Z(n46031) );
  AND U46421 ( .A(b[6]), .B(a[18]), .Z(n46030) );
  XOR U46422 ( .A(n46036), .B(n46037), .Z(n45897) );
  ANDN U46423 ( .B(n46038), .A(n46039), .Z(n46036) );
  AND U46424 ( .A(b[5]), .B(a[19]), .Z(n46035) );
  XOR U46425 ( .A(n46041), .B(n46042), .Z(n45902) );
  ANDN U46426 ( .B(n46043), .A(n46044), .Z(n46041) );
  AND U46427 ( .A(b[4]), .B(a[20]), .Z(n46040) );
  XOR U46428 ( .A(n46046), .B(n46047), .Z(n45907) );
  ANDN U46429 ( .B(n45919), .A(n45920), .Z(n46046) );
  AND U46430 ( .A(b[2]), .B(a[21]), .Z(n46048) );
  XNOR U46431 ( .A(n46043), .B(n46047), .Z(n46049) );
  XOR U46432 ( .A(n46050), .B(n46051), .Z(n46047) );
  OR U46433 ( .A(n45922), .B(n45923), .Z(n46051) );
  XNOR U46434 ( .A(n46053), .B(n46054), .Z(n46052) );
  XOR U46435 ( .A(n46053), .B(n46056), .Z(n45922) );
  NAND U46436 ( .A(b[1]), .B(a[21]), .Z(n46056) );
  IV U46437 ( .A(n46050), .Z(n46053) );
  NANDN U46438 ( .A(n173), .B(n174), .Z(n46050) );
  XOR U46439 ( .A(n46057), .B(n46058), .Z(n174) );
  NAND U46440 ( .A(a[21]), .B(b[0]), .Z(n173) );
  XNOR U46441 ( .A(n46038), .B(n46042), .Z(n46059) );
  XNOR U46442 ( .A(n46033), .B(n46037), .Z(n46060) );
  XNOR U46443 ( .A(n46028), .B(n46032), .Z(n46061) );
  XNOR U46444 ( .A(n46023), .B(n46027), .Z(n46062) );
  XNOR U46445 ( .A(n46018), .B(n46022), .Z(n46063) );
  XNOR U46446 ( .A(n46013), .B(n46017), .Z(n46064) );
  XNOR U46447 ( .A(n46008), .B(n46012), .Z(n46065) );
  XNOR U46448 ( .A(n46003), .B(n46007), .Z(n46066) );
  XNOR U46449 ( .A(n45998), .B(n46002), .Z(n46067) );
  XNOR U46450 ( .A(n45993), .B(n45997), .Z(n46068) );
  XNOR U46451 ( .A(n45988), .B(n45992), .Z(n46069) );
  XNOR U46452 ( .A(n45983), .B(n45987), .Z(n46070) );
  XNOR U46453 ( .A(n45978), .B(n45982), .Z(n46071) );
  XNOR U46454 ( .A(n45973), .B(n45977), .Z(n46072) );
  XNOR U46455 ( .A(n45968), .B(n45972), .Z(n46073) );
  XNOR U46456 ( .A(n45963), .B(n45967), .Z(n46074) );
  XNOR U46457 ( .A(n45958), .B(n45962), .Z(n46075) );
  XNOR U46458 ( .A(n45953), .B(n45957), .Z(n46076) );
  XNOR U46459 ( .A(n45948), .B(n45952), .Z(n46077) );
  XNOR U46460 ( .A(n46078), .B(n45947), .Z(n45948) );
  AND U46461 ( .A(a[0]), .B(b[23]), .Z(n46078) );
  XOR U46462 ( .A(n46079), .B(n45947), .Z(n45949) );
  XNOR U46463 ( .A(n46080), .B(n46081), .Z(n45947) );
  ANDN U46464 ( .B(n46082), .A(n46083), .Z(n46080) );
  AND U46465 ( .A(a[1]), .B(b[22]), .Z(n46079) );
  XOR U46466 ( .A(n46085), .B(n46086), .Z(n45952) );
  ANDN U46467 ( .B(n46087), .A(n46088), .Z(n46085) );
  AND U46468 ( .A(a[2]), .B(b[21]), .Z(n46084) );
  XOR U46469 ( .A(n46090), .B(n46091), .Z(n45957) );
  ANDN U46470 ( .B(n46092), .A(n46093), .Z(n46090) );
  AND U46471 ( .A(a[3]), .B(b[20]), .Z(n46089) );
  XOR U46472 ( .A(n46095), .B(n46096), .Z(n45962) );
  ANDN U46473 ( .B(n46097), .A(n46098), .Z(n46095) );
  AND U46474 ( .A(a[4]), .B(b[19]), .Z(n46094) );
  XOR U46475 ( .A(n46100), .B(n46101), .Z(n45967) );
  ANDN U46476 ( .B(n46102), .A(n46103), .Z(n46100) );
  AND U46477 ( .A(a[5]), .B(b[18]), .Z(n46099) );
  XOR U46478 ( .A(n46105), .B(n46106), .Z(n45972) );
  ANDN U46479 ( .B(n46107), .A(n46108), .Z(n46105) );
  AND U46480 ( .A(a[6]), .B(b[17]), .Z(n46104) );
  XOR U46481 ( .A(n46110), .B(n46111), .Z(n45977) );
  ANDN U46482 ( .B(n46112), .A(n46113), .Z(n46110) );
  AND U46483 ( .A(a[7]), .B(b[16]), .Z(n46109) );
  XOR U46484 ( .A(n46115), .B(n46116), .Z(n45982) );
  ANDN U46485 ( .B(n46117), .A(n46118), .Z(n46115) );
  AND U46486 ( .A(a[8]), .B(b[15]), .Z(n46114) );
  XOR U46487 ( .A(n46120), .B(n46121), .Z(n45987) );
  ANDN U46488 ( .B(n46122), .A(n46123), .Z(n46120) );
  AND U46489 ( .A(a[9]), .B(b[14]), .Z(n46119) );
  XOR U46490 ( .A(n46125), .B(n46126), .Z(n45992) );
  ANDN U46491 ( .B(n46127), .A(n46128), .Z(n46125) );
  AND U46492 ( .A(a[10]), .B(b[13]), .Z(n46124) );
  XOR U46493 ( .A(n46130), .B(n46131), .Z(n45997) );
  ANDN U46494 ( .B(n46132), .A(n46133), .Z(n46130) );
  AND U46495 ( .A(a[11]), .B(b[12]), .Z(n46129) );
  XOR U46496 ( .A(n46135), .B(n46136), .Z(n46002) );
  ANDN U46497 ( .B(n46137), .A(n46138), .Z(n46135) );
  AND U46498 ( .A(a[12]), .B(b[11]), .Z(n46134) );
  XOR U46499 ( .A(n46140), .B(n46141), .Z(n46007) );
  ANDN U46500 ( .B(n46142), .A(n46143), .Z(n46140) );
  AND U46501 ( .A(a[13]), .B(b[10]), .Z(n46139) );
  XOR U46502 ( .A(n46145), .B(n46146), .Z(n46012) );
  ANDN U46503 ( .B(n46147), .A(n46148), .Z(n46145) );
  AND U46504 ( .A(b[9]), .B(a[14]), .Z(n46144) );
  XOR U46505 ( .A(n46150), .B(n46151), .Z(n46017) );
  ANDN U46506 ( .B(n46152), .A(n46153), .Z(n46150) );
  AND U46507 ( .A(b[8]), .B(a[15]), .Z(n46149) );
  XOR U46508 ( .A(n46155), .B(n46156), .Z(n46022) );
  ANDN U46509 ( .B(n46157), .A(n46158), .Z(n46155) );
  AND U46510 ( .A(b[7]), .B(a[16]), .Z(n46154) );
  XOR U46511 ( .A(n46160), .B(n46161), .Z(n46027) );
  ANDN U46512 ( .B(n46162), .A(n46163), .Z(n46160) );
  AND U46513 ( .A(b[6]), .B(a[17]), .Z(n46159) );
  XOR U46514 ( .A(n46165), .B(n46166), .Z(n46032) );
  ANDN U46515 ( .B(n46167), .A(n46168), .Z(n46165) );
  AND U46516 ( .A(b[5]), .B(a[18]), .Z(n46164) );
  XOR U46517 ( .A(n46170), .B(n46171), .Z(n46037) );
  ANDN U46518 ( .B(n46172), .A(n46173), .Z(n46170) );
  AND U46519 ( .A(b[4]), .B(a[19]), .Z(n46169) );
  XOR U46520 ( .A(n46175), .B(n46176), .Z(n46042) );
  ANDN U46521 ( .B(n46054), .A(n46055), .Z(n46175) );
  AND U46522 ( .A(b[2]), .B(a[20]), .Z(n46177) );
  XNOR U46523 ( .A(n46172), .B(n46176), .Z(n46178) );
  XOR U46524 ( .A(n46179), .B(n46180), .Z(n46176) );
  OR U46525 ( .A(n46057), .B(n46058), .Z(n46180) );
  XNOR U46526 ( .A(n46182), .B(n46183), .Z(n46181) );
  XOR U46527 ( .A(n46182), .B(n46185), .Z(n46057) );
  NAND U46528 ( .A(b[1]), .B(a[20]), .Z(n46185) );
  IV U46529 ( .A(n46179), .Z(n46182) );
  NANDN U46530 ( .A(n175), .B(n176), .Z(n46179) );
  XOR U46531 ( .A(n46186), .B(n46187), .Z(n176) );
  NAND U46532 ( .A(a[20]), .B(b[0]), .Z(n175) );
  XNOR U46533 ( .A(n46167), .B(n46171), .Z(n46188) );
  XNOR U46534 ( .A(n46162), .B(n46166), .Z(n46189) );
  XNOR U46535 ( .A(n46157), .B(n46161), .Z(n46190) );
  XNOR U46536 ( .A(n46152), .B(n46156), .Z(n46191) );
  XNOR U46537 ( .A(n46147), .B(n46151), .Z(n46192) );
  XNOR U46538 ( .A(n46142), .B(n46146), .Z(n46193) );
  XNOR U46539 ( .A(n46137), .B(n46141), .Z(n46194) );
  XNOR U46540 ( .A(n46132), .B(n46136), .Z(n46195) );
  XNOR U46541 ( .A(n46127), .B(n46131), .Z(n46196) );
  XNOR U46542 ( .A(n46122), .B(n46126), .Z(n46197) );
  XNOR U46543 ( .A(n46117), .B(n46121), .Z(n46198) );
  XNOR U46544 ( .A(n46112), .B(n46116), .Z(n46199) );
  XNOR U46545 ( .A(n46107), .B(n46111), .Z(n46200) );
  XNOR U46546 ( .A(n46102), .B(n46106), .Z(n46201) );
  XNOR U46547 ( .A(n46097), .B(n46101), .Z(n46202) );
  XNOR U46548 ( .A(n46092), .B(n46096), .Z(n46203) );
  XNOR U46549 ( .A(n46087), .B(n46091), .Z(n46204) );
  XNOR U46550 ( .A(n46082), .B(n46086), .Z(n46205) );
  XOR U46551 ( .A(n46206), .B(n46081), .Z(n46082) );
  AND U46552 ( .A(a[0]), .B(b[22]), .Z(n46206) );
  XNOR U46553 ( .A(n46207), .B(n46081), .Z(n46083) );
  XNOR U46554 ( .A(n46208), .B(n46209), .Z(n46081) );
  ANDN U46555 ( .B(n46210), .A(n46211), .Z(n46208) );
  AND U46556 ( .A(a[1]), .B(b[21]), .Z(n46207) );
  XOR U46557 ( .A(n46213), .B(n46214), .Z(n46086) );
  ANDN U46558 ( .B(n46215), .A(n46216), .Z(n46213) );
  AND U46559 ( .A(a[2]), .B(b[20]), .Z(n46212) );
  XOR U46560 ( .A(n46218), .B(n46219), .Z(n46091) );
  ANDN U46561 ( .B(n46220), .A(n46221), .Z(n46218) );
  AND U46562 ( .A(a[3]), .B(b[19]), .Z(n46217) );
  XOR U46563 ( .A(n46223), .B(n46224), .Z(n46096) );
  ANDN U46564 ( .B(n46225), .A(n46226), .Z(n46223) );
  AND U46565 ( .A(a[4]), .B(b[18]), .Z(n46222) );
  XOR U46566 ( .A(n46228), .B(n46229), .Z(n46101) );
  ANDN U46567 ( .B(n46230), .A(n46231), .Z(n46228) );
  AND U46568 ( .A(a[5]), .B(b[17]), .Z(n46227) );
  XOR U46569 ( .A(n46233), .B(n46234), .Z(n46106) );
  ANDN U46570 ( .B(n46235), .A(n46236), .Z(n46233) );
  AND U46571 ( .A(a[6]), .B(b[16]), .Z(n46232) );
  XOR U46572 ( .A(n46238), .B(n46239), .Z(n46111) );
  ANDN U46573 ( .B(n46240), .A(n46241), .Z(n46238) );
  AND U46574 ( .A(a[7]), .B(b[15]), .Z(n46237) );
  XOR U46575 ( .A(n46243), .B(n46244), .Z(n46116) );
  ANDN U46576 ( .B(n46245), .A(n46246), .Z(n46243) );
  AND U46577 ( .A(a[8]), .B(b[14]), .Z(n46242) );
  XOR U46578 ( .A(n46248), .B(n46249), .Z(n46121) );
  ANDN U46579 ( .B(n46250), .A(n46251), .Z(n46248) );
  AND U46580 ( .A(a[9]), .B(b[13]), .Z(n46247) );
  XOR U46581 ( .A(n46253), .B(n46254), .Z(n46126) );
  ANDN U46582 ( .B(n46255), .A(n46256), .Z(n46253) );
  AND U46583 ( .A(a[10]), .B(b[12]), .Z(n46252) );
  XOR U46584 ( .A(n46258), .B(n46259), .Z(n46131) );
  ANDN U46585 ( .B(n46260), .A(n46261), .Z(n46258) );
  AND U46586 ( .A(a[11]), .B(b[11]), .Z(n46257) );
  XOR U46587 ( .A(n46263), .B(n46264), .Z(n46136) );
  ANDN U46588 ( .B(n46265), .A(n46266), .Z(n46263) );
  AND U46589 ( .A(a[12]), .B(b[10]), .Z(n46262) );
  XOR U46590 ( .A(n46268), .B(n46269), .Z(n46141) );
  ANDN U46591 ( .B(n46270), .A(n46271), .Z(n46268) );
  AND U46592 ( .A(b[9]), .B(a[13]), .Z(n46267) );
  XOR U46593 ( .A(n46273), .B(n46274), .Z(n46146) );
  ANDN U46594 ( .B(n46275), .A(n46276), .Z(n46273) );
  AND U46595 ( .A(b[8]), .B(a[14]), .Z(n46272) );
  XOR U46596 ( .A(n46278), .B(n46279), .Z(n46151) );
  ANDN U46597 ( .B(n46280), .A(n46281), .Z(n46278) );
  AND U46598 ( .A(b[7]), .B(a[15]), .Z(n46277) );
  XOR U46599 ( .A(n46283), .B(n46284), .Z(n46156) );
  ANDN U46600 ( .B(n46285), .A(n46286), .Z(n46283) );
  AND U46601 ( .A(b[6]), .B(a[16]), .Z(n46282) );
  XOR U46602 ( .A(n46288), .B(n46289), .Z(n46161) );
  ANDN U46603 ( .B(n46290), .A(n46291), .Z(n46288) );
  AND U46604 ( .A(b[5]), .B(a[17]), .Z(n46287) );
  XOR U46605 ( .A(n46293), .B(n46294), .Z(n46166) );
  ANDN U46606 ( .B(n46295), .A(n46296), .Z(n46293) );
  AND U46607 ( .A(b[4]), .B(a[18]), .Z(n46292) );
  XOR U46608 ( .A(n46298), .B(n46299), .Z(n46171) );
  ANDN U46609 ( .B(n46183), .A(n46184), .Z(n46298) );
  AND U46610 ( .A(b[2]), .B(a[19]), .Z(n46300) );
  XNOR U46611 ( .A(n46295), .B(n46299), .Z(n46301) );
  XOR U46612 ( .A(n46302), .B(n46303), .Z(n46299) );
  OR U46613 ( .A(n46186), .B(n46187), .Z(n46303) );
  XNOR U46614 ( .A(n46305), .B(n46306), .Z(n46304) );
  XOR U46615 ( .A(n46305), .B(n46308), .Z(n46186) );
  NAND U46616 ( .A(b[1]), .B(a[19]), .Z(n46308) );
  IV U46617 ( .A(n46302), .Z(n46305) );
  NANDN U46618 ( .A(n179), .B(n180), .Z(n46302) );
  XOR U46619 ( .A(n46309), .B(n46310), .Z(n180) );
  NAND U46620 ( .A(a[19]), .B(b[0]), .Z(n179) );
  XNOR U46621 ( .A(n46290), .B(n46294), .Z(n46311) );
  XNOR U46622 ( .A(n46285), .B(n46289), .Z(n46312) );
  XNOR U46623 ( .A(n46280), .B(n46284), .Z(n46313) );
  XNOR U46624 ( .A(n46275), .B(n46279), .Z(n46314) );
  XNOR U46625 ( .A(n46270), .B(n46274), .Z(n46315) );
  XNOR U46626 ( .A(n46265), .B(n46269), .Z(n46316) );
  XNOR U46627 ( .A(n46260), .B(n46264), .Z(n46317) );
  XNOR U46628 ( .A(n46255), .B(n46259), .Z(n46318) );
  XNOR U46629 ( .A(n46250), .B(n46254), .Z(n46319) );
  XNOR U46630 ( .A(n46245), .B(n46249), .Z(n46320) );
  XNOR U46631 ( .A(n46240), .B(n46244), .Z(n46321) );
  XNOR U46632 ( .A(n46235), .B(n46239), .Z(n46322) );
  XNOR U46633 ( .A(n46230), .B(n46234), .Z(n46323) );
  XNOR U46634 ( .A(n46225), .B(n46229), .Z(n46324) );
  XNOR U46635 ( .A(n46220), .B(n46224), .Z(n46325) );
  XNOR U46636 ( .A(n46215), .B(n46219), .Z(n46326) );
  XNOR U46637 ( .A(n46210), .B(n46214), .Z(n46327) );
  XNOR U46638 ( .A(n46328), .B(n46209), .Z(n46210) );
  AND U46639 ( .A(a[0]), .B(b[21]), .Z(n46328) );
  XOR U46640 ( .A(n46329), .B(n46209), .Z(n46211) );
  XNOR U46641 ( .A(n46330), .B(n46331), .Z(n46209) );
  ANDN U46642 ( .B(n46332), .A(n46333), .Z(n46330) );
  AND U46643 ( .A(a[1]), .B(b[20]), .Z(n46329) );
  XOR U46644 ( .A(n46335), .B(n46336), .Z(n46214) );
  ANDN U46645 ( .B(n46337), .A(n46338), .Z(n46335) );
  AND U46646 ( .A(a[2]), .B(b[19]), .Z(n46334) );
  XOR U46647 ( .A(n46340), .B(n46341), .Z(n46219) );
  ANDN U46648 ( .B(n46342), .A(n46343), .Z(n46340) );
  AND U46649 ( .A(a[3]), .B(b[18]), .Z(n46339) );
  XOR U46650 ( .A(n46345), .B(n46346), .Z(n46224) );
  ANDN U46651 ( .B(n46347), .A(n46348), .Z(n46345) );
  AND U46652 ( .A(a[4]), .B(b[17]), .Z(n46344) );
  XOR U46653 ( .A(n46350), .B(n46351), .Z(n46229) );
  ANDN U46654 ( .B(n46352), .A(n46353), .Z(n46350) );
  AND U46655 ( .A(a[5]), .B(b[16]), .Z(n46349) );
  XOR U46656 ( .A(n46355), .B(n46356), .Z(n46234) );
  ANDN U46657 ( .B(n46357), .A(n46358), .Z(n46355) );
  AND U46658 ( .A(a[6]), .B(b[15]), .Z(n46354) );
  XOR U46659 ( .A(n46360), .B(n46361), .Z(n46239) );
  ANDN U46660 ( .B(n46362), .A(n46363), .Z(n46360) );
  AND U46661 ( .A(a[7]), .B(b[14]), .Z(n46359) );
  XOR U46662 ( .A(n46365), .B(n46366), .Z(n46244) );
  ANDN U46663 ( .B(n46367), .A(n46368), .Z(n46365) );
  AND U46664 ( .A(a[8]), .B(b[13]), .Z(n46364) );
  XOR U46665 ( .A(n46370), .B(n46371), .Z(n46249) );
  ANDN U46666 ( .B(n46372), .A(n46373), .Z(n46370) );
  AND U46667 ( .A(a[9]), .B(b[12]), .Z(n46369) );
  XOR U46668 ( .A(n46375), .B(n46376), .Z(n46254) );
  ANDN U46669 ( .B(n46377), .A(n46378), .Z(n46375) );
  AND U46670 ( .A(a[10]), .B(b[11]), .Z(n46374) );
  XOR U46671 ( .A(n46380), .B(n46381), .Z(n46259) );
  ANDN U46672 ( .B(n46382), .A(n46383), .Z(n46380) );
  AND U46673 ( .A(a[11]), .B(b[10]), .Z(n46379) );
  XOR U46674 ( .A(n46385), .B(n46386), .Z(n46264) );
  ANDN U46675 ( .B(n46387), .A(n46388), .Z(n46385) );
  AND U46676 ( .A(b[9]), .B(a[12]), .Z(n46384) );
  XOR U46677 ( .A(n46390), .B(n46391), .Z(n46269) );
  ANDN U46678 ( .B(n46392), .A(n46393), .Z(n46390) );
  AND U46679 ( .A(b[8]), .B(a[13]), .Z(n46389) );
  XOR U46680 ( .A(n46395), .B(n46396), .Z(n46274) );
  ANDN U46681 ( .B(n46397), .A(n46398), .Z(n46395) );
  AND U46682 ( .A(b[7]), .B(a[14]), .Z(n46394) );
  XOR U46683 ( .A(n46400), .B(n46401), .Z(n46279) );
  ANDN U46684 ( .B(n46402), .A(n46403), .Z(n46400) );
  AND U46685 ( .A(b[6]), .B(a[15]), .Z(n46399) );
  XOR U46686 ( .A(n46405), .B(n46406), .Z(n46284) );
  ANDN U46687 ( .B(n46407), .A(n46408), .Z(n46405) );
  AND U46688 ( .A(b[5]), .B(a[16]), .Z(n46404) );
  XOR U46689 ( .A(n46410), .B(n46411), .Z(n46289) );
  ANDN U46690 ( .B(n46412), .A(n46413), .Z(n46410) );
  AND U46691 ( .A(b[4]), .B(a[17]), .Z(n46409) );
  XOR U46692 ( .A(n46415), .B(n46416), .Z(n46294) );
  ANDN U46693 ( .B(n46306), .A(n46307), .Z(n46415) );
  AND U46694 ( .A(b[2]), .B(a[18]), .Z(n46417) );
  XNOR U46695 ( .A(n46412), .B(n46416), .Z(n46418) );
  XOR U46696 ( .A(n46419), .B(n46420), .Z(n46416) );
  OR U46697 ( .A(n46309), .B(n46310), .Z(n46420) );
  XNOR U46698 ( .A(n46422), .B(n46423), .Z(n46421) );
  XOR U46699 ( .A(n46422), .B(n46425), .Z(n46309) );
  NAND U46700 ( .A(b[1]), .B(a[18]), .Z(n46425) );
  IV U46701 ( .A(n46419), .Z(n46422) );
  NANDN U46702 ( .A(n181), .B(n182), .Z(n46419) );
  XOR U46703 ( .A(n46426), .B(n46427), .Z(n182) );
  NAND U46704 ( .A(a[18]), .B(b[0]), .Z(n181) );
  XNOR U46705 ( .A(n46407), .B(n46411), .Z(n46428) );
  XNOR U46706 ( .A(n46402), .B(n46406), .Z(n46429) );
  XNOR U46707 ( .A(n46397), .B(n46401), .Z(n46430) );
  XNOR U46708 ( .A(n46392), .B(n46396), .Z(n46431) );
  XNOR U46709 ( .A(n46387), .B(n46391), .Z(n46432) );
  XNOR U46710 ( .A(n46382), .B(n46386), .Z(n46433) );
  XNOR U46711 ( .A(n46377), .B(n46381), .Z(n46434) );
  XNOR U46712 ( .A(n46372), .B(n46376), .Z(n46435) );
  XNOR U46713 ( .A(n46367), .B(n46371), .Z(n46436) );
  XNOR U46714 ( .A(n46362), .B(n46366), .Z(n46437) );
  XNOR U46715 ( .A(n46357), .B(n46361), .Z(n46438) );
  XNOR U46716 ( .A(n46352), .B(n46356), .Z(n46439) );
  XNOR U46717 ( .A(n46347), .B(n46351), .Z(n46440) );
  XNOR U46718 ( .A(n46342), .B(n46346), .Z(n46441) );
  XNOR U46719 ( .A(n46337), .B(n46341), .Z(n46442) );
  XNOR U46720 ( .A(n46332), .B(n46336), .Z(n46443) );
  XOR U46721 ( .A(n46444), .B(n46331), .Z(n46332) );
  AND U46722 ( .A(a[0]), .B(b[20]), .Z(n46444) );
  XNOR U46723 ( .A(n46445), .B(n46331), .Z(n46333) );
  XNOR U46724 ( .A(n46446), .B(n46447), .Z(n46331) );
  ANDN U46725 ( .B(n46448), .A(n46449), .Z(n46446) );
  AND U46726 ( .A(a[1]), .B(b[19]), .Z(n46445) );
  XOR U46727 ( .A(n46451), .B(n46452), .Z(n46336) );
  ANDN U46728 ( .B(n46453), .A(n46454), .Z(n46451) );
  AND U46729 ( .A(a[2]), .B(b[18]), .Z(n46450) );
  XOR U46730 ( .A(n46456), .B(n46457), .Z(n46341) );
  ANDN U46731 ( .B(n46458), .A(n46459), .Z(n46456) );
  AND U46732 ( .A(a[3]), .B(b[17]), .Z(n46455) );
  XOR U46733 ( .A(n46461), .B(n46462), .Z(n46346) );
  ANDN U46734 ( .B(n46463), .A(n46464), .Z(n46461) );
  AND U46735 ( .A(a[4]), .B(b[16]), .Z(n46460) );
  XOR U46736 ( .A(n46466), .B(n46467), .Z(n46351) );
  ANDN U46737 ( .B(n46468), .A(n46469), .Z(n46466) );
  AND U46738 ( .A(a[5]), .B(b[15]), .Z(n46465) );
  XOR U46739 ( .A(n46471), .B(n46472), .Z(n46356) );
  ANDN U46740 ( .B(n46473), .A(n46474), .Z(n46471) );
  AND U46741 ( .A(a[6]), .B(b[14]), .Z(n46470) );
  XOR U46742 ( .A(n46476), .B(n46477), .Z(n46361) );
  ANDN U46743 ( .B(n46478), .A(n46479), .Z(n46476) );
  AND U46744 ( .A(a[7]), .B(b[13]), .Z(n46475) );
  XOR U46745 ( .A(n46481), .B(n46482), .Z(n46366) );
  ANDN U46746 ( .B(n46483), .A(n46484), .Z(n46481) );
  AND U46747 ( .A(a[8]), .B(b[12]), .Z(n46480) );
  XOR U46748 ( .A(n46486), .B(n46487), .Z(n46371) );
  ANDN U46749 ( .B(n46488), .A(n46489), .Z(n46486) );
  AND U46750 ( .A(a[9]), .B(b[11]), .Z(n46485) );
  XOR U46751 ( .A(n46491), .B(n46492), .Z(n46376) );
  ANDN U46752 ( .B(n46493), .A(n46494), .Z(n46491) );
  AND U46753 ( .A(a[10]), .B(b[10]), .Z(n46490) );
  XOR U46754 ( .A(n46496), .B(n46497), .Z(n46381) );
  ANDN U46755 ( .B(n46498), .A(n46499), .Z(n46496) );
  AND U46756 ( .A(b[9]), .B(a[11]), .Z(n46495) );
  XOR U46757 ( .A(n46501), .B(n46502), .Z(n46386) );
  ANDN U46758 ( .B(n46503), .A(n46504), .Z(n46501) );
  AND U46759 ( .A(b[8]), .B(a[12]), .Z(n46500) );
  XOR U46760 ( .A(n46506), .B(n46507), .Z(n46391) );
  ANDN U46761 ( .B(n46508), .A(n46509), .Z(n46506) );
  AND U46762 ( .A(b[7]), .B(a[13]), .Z(n46505) );
  XOR U46763 ( .A(n46511), .B(n46512), .Z(n46396) );
  ANDN U46764 ( .B(n46513), .A(n46514), .Z(n46511) );
  AND U46765 ( .A(b[6]), .B(a[14]), .Z(n46510) );
  XOR U46766 ( .A(n46516), .B(n46517), .Z(n46401) );
  ANDN U46767 ( .B(n46518), .A(n46519), .Z(n46516) );
  AND U46768 ( .A(b[5]), .B(a[15]), .Z(n46515) );
  XOR U46769 ( .A(n46521), .B(n46522), .Z(n46406) );
  ANDN U46770 ( .B(n46523), .A(n46524), .Z(n46521) );
  AND U46771 ( .A(b[4]), .B(a[16]), .Z(n46520) );
  XOR U46772 ( .A(n46526), .B(n46527), .Z(n46411) );
  ANDN U46773 ( .B(n46423), .A(n46424), .Z(n46526) );
  AND U46774 ( .A(b[2]), .B(a[17]), .Z(n46528) );
  XNOR U46775 ( .A(n46523), .B(n46527), .Z(n46529) );
  XOR U46776 ( .A(n46530), .B(n46531), .Z(n46527) );
  OR U46777 ( .A(n46426), .B(n46427), .Z(n46531) );
  XNOR U46778 ( .A(n46533), .B(n46534), .Z(n46532) );
  XOR U46779 ( .A(n46533), .B(n46536), .Z(n46426) );
  NAND U46780 ( .A(b[1]), .B(a[17]), .Z(n46536) );
  IV U46781 ( .A(n46530), .Z(n46533) );
  NANDN U46782 ( .A(n183), .B(n184), .Z(n46530) );
  XOR U46783 ( .A(n46537), .B(n46538), .Z(n184) );
  NAND U46784 ( .A(a[17]), .B(b[0]), .Z(n183) );
  XNOR U46785 ( .A(n46518), .B(n46522), .Z(n46539) );
  XNOR U46786 ( .A(n46513), .B(n46517), .Z(n46540) );
  XNOR U46787 ( .A(n46508), .B(n46512), .Z(n46541) );
  XNOR U46788 ( .A(n46503), .B(n46507), .Z(n46542) );
  XNOR U46789 ( .A(n46498), .B(n46502), .Z(n46543) );
  XNOR U46790 ( .A(n46493), .B(n46497), .Z(n46544) );
  XNOR U46791 ( .A(n46488), .B(n46492), .Z(n46545) );
  XNOR U46792 ( .A(n46483), .B(n46487), .Z(n46546) );
  XNOR U46793 ( .A(n46478), .B(n46482), .Z(n46547) );
  XNOR U46794 ( .A(n46473), .B(n46477), .Z(n46548) );
  XNOR U46795 ( .A(n46468), .B(n46472), .Z(n46549) );
  XNOR U46796 ( .A(n46463), .B(n46467), .Z(n46550) );
  XNOR U46797 ( .A(n46458), .B(n46462), .Z(n46551) );
  XNOR U46798 ( .A(n46453), .B(n46457), .Z(n46552) );
  XNOR U46799 ( .A(n46448), .B(n46452), .Z(n46553) );
  XNOR U46800 ( .A(n46554), .B(n46447), .Z(n46448) );
  AND U46801 ( .A(a[0]), .B(b[19]), .Z(n46554) );
  XOR U46802 ( .A(n46555), .B(n46447), .Z(n46449) );
  XNOR U46803 ( .A(n46556), .B(n46557), .Z(n46447) );
  ANDN U46804 ( .B(n46558), .A(n46559), .Z(n46556) );
  AND U46805 ( .A(a[1]), .B(b[18]), .Z(n46555) );
  XOR U46806 ( .A(n46561), .B(n46562), .Z(n46452) );
  ANDN U46807 ( .B(n46563), .A(n46564), .Z(n46561) );
  AND U46808 ( .A(a[2]), .B(b[17]), .Z(n46560) );
  XOR U46809 ( .A(n46566), .B(n46567), .Z(n46457) );
  ANDN U46810 ( .B(n46568), .A(n46569), .Z(n46566) );
  AND U46811 ( .A(a[3]), .B(b[16]), .Z(n46565) );
  XOR U46812 ( .A(n46571), .B(n46572), .Z(n46462) );
  ANDN U46813 ( .B(n46573), .A(n46574), .Z(n46571) );
  AND U46814 ( .A(a[4]), .B(b[15]), .Z(n46570) );
  XOR U46815 ( .A(n46576), .B(n46577), .Z(n46467) );
  ANDN U46816 ( .B(n46578), .A(n46579), .Z(n46576) );
  AND U46817 ( .A(a[5]), .B(b[14]), .Z(n46575) );
  XOR U46818 ( .A(n46581), .B(n46582), .Z(n46472) );
  ANDN U46819 ( .B(n46583), .A(n46584), .Z(n46581) );
  AND U46820 ( .A(a[6]), .B(b[13]), .Z(n46580) );
  XOR U46821 ( .A(n46586), .B(n46587), .Z(n46477) );
  ANDN U46822 ( .B(n46588), .A(n46589), .Z(n46586) );
  AND U46823 ( .A(a[7]), .B(b[12]), .Z(n46585) );
  XOR U46824 ( .A(n46591), .B(n46592), .Z(n46482) );
  ANDN U46825 ( .B(n46593), .A(n46594), .Z(n46591) );
  AND U46826 ( .A(a[8]), .B(b[11]), .Z(n46590) );
  XOR U46827 ( .A(n46596), .B(n46597), .Z(n46487) );
  ANDN U46828 ( .B(n46598), .A(n46599), .Z(n46596) );
  AND U46829 ( .A(a[9]), .B(b[10]), .Z(n46595) );
  XOR U46830 ( .A(n46601), .B(n46602), .Z(n46492) );
  ANDN U46831 ( .B(n46603), .A(n46604), .Z(n46601) );
  AND U46832 ( .A(b[9]), .B(a[10]), .Z(n46600) );
  XOR U46833 ( .A(n46606), .B(n46607), .Z(n46497) );
  ANDN U46834 ( .B(n46608), .A(n46609), .Z(n46606) );
  AND U46835 ( .A(b[8]), .B(a[11]), .Z(n46605) );
  XOR U46836 ( .A(n46611), .B(n46612), .Z(n46502) );
  ANDN U46837 ( .B(n46613), .A(n46614), .Z(n46611) );
  AND U46838 ( .A(b[7]), .B(a[12]), .Z(n46610) );
  XOR U46839 ( .A(n46616), .B(n46617), .Z(n46507) );
  ANDN U46840 ( .B(n46618), .A(n46619), .Z(n46616) );
  AND U46841 ( .A(b[6]), .B(a[13]), .Z(n46615) );
  XOR U46842 ( .A(n46621), .B(n46622), .Z(n46512) );
  ANDN U46843 ( .B(n46623), .A(n46624), .Z(n46621) );
  AND U46844 ( .A(b[5]), .B(a[14]), .Z(n46620) );
  XOR U46845 ( .A(n46626), .B(n46627), .Z(n46517) );
  ANDN U46846 ( .B(n46628), .A(n46629), .Z(n46626) );
  AND U46847 ( .A(b[4]), .B(a[15]), .Z(n46625) );
  XOR U46848 ( .A(n46631), .B(n46632), .Z(n46522) );
  ANDN U46849 ( .B(n46534), .A(n46535), .Z(n46631) );
  AND U46850 ( .A(b[2]), .B(a[16]), .Z(n46633) );
  XNOR U46851 ( .A(n46628), .B(n46632), .Z(n46634) );
  XOR U46852 ( .A(n46635), .B(n46636), .Z(n46632) );
  OR U46853 ( .A(n46537), .B(n46538), .Z(n46636) );
  XNOR U46854 ( .A(n46638), .B(n46639), .Z(n46637) );
  XOR U46855 ( .A(n46638), .B(n46641), .Z(n46537) );
  NAND U46856 ( .A(b[1]), .B(a[16]), .Z(n46641) );
  IV U46857 ( .A(n46635), .Z(n46638) );
  NANDN U46858 ( .A(n185), .B(n186), .Z(n46635) );
  XOR U46859 ( .A(n46642), .B(n46643), .Z(n186) );
  NAND U46860 ( .A(a[16]), .B(b[0]), .Z(n185) );
  XNOR U46861 ( .A(n46623), .B(n46627), .Z(n46644) );
  XNOR U46862 ( .A(n46618), .B(n46622), .Z(n46645) );
  XNOR U46863 ( .A(n46613), .B(n46617), .Z(n46646) );
  XNOR U46864 ( .A(n46608), .B(n46612), .Z(n46647) );
  XNOR U46865 ( .A(n46603), .B(n46607), .Z(n46648) );
  XNOR U46866 ( .A(n46598), .B(n46602), .Z(n46649) );
  XNOR U46867 ( .A(n46593), .B(n46597), .Z(n46650) );
  XNOR U46868 ( .A(n46588), .B(n46592), .Z(n46651) );
  XNOR U46869 ( .A(n46583), .B(n46587), .Z(n46652) );
  XNOR U46870 ( .A(n46578), .B(n46582), .Z(n46653) );
  XNOR U46871 ( .A(n46573), .B(n46577), .Z(n46654) );
  XNOR U46872 ( .A(n46568), .B(n46572), .Z(n46655) );
  XNOR U46873 ( .A(n46563), .B(n46567), .Z(n46656) );
  XNOR U46874 ( .A(n46558), .B(n46562), .Z(n46657) );
  XOR U46875 ( .A(n46658), .B(n46557), .Z(n46558) );
  AND U46876 ( .A(a[0]), .B(b[18]), .Z(n46658) );
  XNOR U46877 ( .A(n46659), .B(n46557), .Z(n46559) );
  XNOR U46878 ( .A(n46660), .B(n46661), .Z(n46557) );
  ANDN U46879 ( .B(n46662), .A(n46663), .Z(n46660) );
  AND U46880 ( .A(a[1]), .B(b[17]), .Z(n46659) );
  XOR U46881 ( .A(n46665), .B(n46666), .Z(n46562) );
  ANDN U46882 ( .B(n46667), .A(n46668), .Z(n46665) );
  AND U46883 ( .A(a[2]), .B(b[16]), .Z(n46664) );
  XOR U46884 ( .A(n46670), .B(n46671), .Z(n46567) );
  ANDN U46885 ( .B(n46672), .A(n46673), .Z(n46670) );
  AND U46886 ( .A(a[3]), .B(b[15]), .Z(n46669) );
  XOR U46887 ( .A(n46675), .B(n46676), .Z(n46572) );
  ANDN U46888 ( .B(n46677), .A(n46678), .Z(n46675) );
  AND U46889 ( .A(a[4]), .B(b[14]), .Z(n46674) );
  XOR U46890 ( .A(n46680), .B(n46681), .Z(n46577) );
  ANDN U46891 ( .B(n46682), .A(n46683), .Z(n46680) );
  AND U46892 ( .A(a[5]), .B(b[13]), .Z(n46679) );
  XOR U46893 ( .A(n46685), .B(n46686), .Z(n46582) );
  ANDN U46894 ( .B(n46687), .A(n46688), .Z(n46685) );
  AND U46895 ( .A(a[6]), .B(b[12]), .Z(n46684) );
  XOR U46896 ( .A(n46690), .B(n46691), .Z(n46587) );
  ANDN U46897 ( .B(n46692), .A(n46693), .Z(n46690) );
  AND U46898 ( .A(a[7]), .B(b[11]), .Z(n46689) );
  XOR U46899 ( .A(n46695), .B(n46696), .Z(n46592) );
  ANDN U46900 ( .B(n46697), .A(n46698), .Z(n46695) );
  AND U46901 ( .A(a[8]), .B(b[10]), .Z(n46694) );
  XOR U46902 ( .A(n46700), .B(n46701), .Z(n46597) );
  ANDN U46903 ( .B(n46702), .A(n46703), .Z(n46700) );
  AND U46904 ( .A(a[9]), .B(b[9]), .Z(n46699) );
  XOR U46905 ( .A(n46705), .B(n46706), .Z(n46602) );
  ANDN U46906 ( .B(n46707), .A(n46708), .Z(n46705) );
  AND U46907 ( .A(b[8]), .B(a[10]), .Z(n46704) );
  XOR U46908 ( .A(n46710), .B(n46711), .Z(n46607) );
  ANDN U46909 ( .B(n46712), .A(n46713), .Z(n46710) );
  AND U46910 ( .A(b[7]), .B(a[11]), .Z(n46709) );
  XOR U46911 ( .A(n46715), .B(n46716), .Z(n46612) );
  ANDN U46912 ( .B(n46717), .A(n46718), .Z(n46715) );
  AND U46913 ( .A(b[6]), .B(a[12]), .Z(n46714) );
  XOR U46914 ( .A(n46720), .B(n46721), .Z(n46617) );
  ANDN U46915 ( .B(n46722), .A(n46723), .Z(n46720) );
  AND U46916 ( .A(b[5]), .B(a[13]), .Z(n46719) );
  XOR U46917 ( .A(n46725), .B(n46726), .Z(n46622) );
  ANDN U46918 ( .B(n46727), .A(n46728), .Z(n46725) );
  AND U46919 ( .A(b[4]), .B(a[14]), .Z(n46724) );
  XOR U46920 ( .A(n46730), .B(n46731), .Z(n46627) );
  ANDN U46921 ( .B(n46639), .A(n46640), .Z(n46730) );
  AND U46922 ( .A(b[2]), .B(a[15]), .Z(n46732) );
  XNOR U46923 ( .A(n46727), .B(n46731), .Z(n46733) );
  XOR U46924 ( .A(n46734), .B(n46735), .Z(n46731) );
  OR U46925 ( .A(n46642), .B(n46643), .Z(n46735) );
  XNOR U46926 ( .A(n46737), .B(n46738), .Z(n46736) );
  XOR U46927 ( .A(n46737), .B(n46740), .Z(n46642) );
  NAND U46928 ( .A(b[1]), .B(a[15]), .Z(n46740) );
  IV U46929 ( .A(n46734), .Z(n46737) );
  NANDN U46930 ( .A(n187), .B(n188), .Z(n46734) );
  XOR U46931 ( .A(n46741), .B(n46742), .Z(n188) );
  NAND U46932 ( .A(a[15]), .B(b[0]), .Z(n187) );
  XNOR U46933 ( .A(n46722), .B(n46726), .Z(n46743) );
  XNOR U46934 ( .A(n46717), .B(n46721), .Z(n46744) );
  XNOR U46935 ( .A(n46712), .B(n46716), .Z(n46745) );
  XNOR U46936 ( .A(n46707), .B(n46711), .Z(n46746) );
  XNOR U46937 ( .A(n46702), .B(n46706), .Z(n46747) );
  XNOR U46938 ( .A(n46697), .B(n46701), .Z(n46748) );
  XNOR U46939 ( .A(n46692), .B(n46696), .Z(n46749) );
  XNOR U46940 ( .A(n46687), .B(n46691), .Z(n46750) );
  XNOR U46941 ( .A(n46682), .B(n46686), .Z(n46751) );
  XNOR U46942 ( .A(n46677), .B(n46681), .Z(n46752) );
  XNOR U46943 ( .A(n46672), .B(n46676), .Z(n46753) );
  XNOR U46944 ( .A(n46667), .B(n46671), .Z(n46754) );
  XNOR U46945 ( .A(n46662), .B(n46666), .Z(n46755) );
  XNOR U46946 ( .A(n46756), .B(n46661), .Z(n46662) );
  AND U46947 ( .A(a[0]), .B(b[17]), .Z(n46756) );
  XOR U46948 ( .A(n46757), .B(n46661), .Z(n46663) );
  XNOR U46949 ( .A(n46758), .B(n46759), .Z(n46661) );
  ANDN U46950 ( .B(n46760), .A(n46761), .Z(n46758) );
  AND U46951 ( .A(a[1]), .B(b[16]), .Z(n46757) );
  XOR U46952 ( .A(n46763), .B(n46764), .Z(n46666) );
  ANDN U46953 ( .B(n46765), .A(n46766), .Z(n46763) );
  AND U46954 ( .A(a[2]), .B(b[15]), .Z(n46762) );
  XOR U46955 ( .A(n46768), .B(n46769), .Z(n46671) );
  ANDN U46956 ( .B(n46770), .A(n46771), .Z(n46768) );
  AND U46957 ( .A(a[3]), .B(b[14]), .Z(n46767) );
  XOR U46958 ( .A(n46773), .B(n46774), .Z(n46676) );
  ANDN U46959 ( .B(n46775), .A(n46776), .Z(n46773) );
  AND U46960 ( .A(a[4]), .B(b[13]), .Z(n46772) );
  XOR U46961 ( .A(n46778), .B(n46779), .Z(n46681) );
  ANDN U46962 ( .B(n46780), .A(n46781), .Z(n46778) );
  AND U46963 ( .A(a[5]), .B(b[12]), .Z(n46777) );
  XOR U46964 ( .A(n46783), .B(n46784), .Z(n46686) );
  ANDN U46965 ( .B(n46785), .A(n46786), .Z(n46783) );
  AND U46966 ( .A(a[6]), .B(b[11]), .Z(n46782) );
  XOR U46967 ( .A(n46788), .B(n46789), .Z(n46691) );
  ANDN U46968 ( .B(n46790), .A(n46791), .Z(n46788) );
  AND U46969 ( .A(a[7]), .B(b[10]), .Z(n46787) );
  XOR U46970 ( .A(n46793), .B(n46794), .Z(n46696) );
  ANDN U46971 ( .B(n46795), .A(n46796), .Z(n46793) );
  AND U46972 ( .A(a[8]), .B(b[9]), .Z(n46792) );
  XOR U46973 ( .A(n46798), .B(n46799), .Z(n46701) );
  ANDN U46974 ( .B(n46800), .A(n46801), .Z(n46798) );
  AND U46975 ( .A(a[9]), .B(b[8]), .Z(n46797) );
  XOR U46976 ( .A(n46803), .B(n46804), .Z(n46706) );
  ANDN U46977 ( .B(n46805), .A(n46806), .Z(n46803) );
  AND U46978 ( .A(b[7]), .B(a[10]), .Z(n46802) );
  XOR U46979 ( .A(n46808), .B(n46809), .Z(n46711) );
  ANDN U46980 ( .B(n46810), .A(n46811), .Z(n46808) );
  AND U46981 ( .A(b[6]), .B(a[11]), .Z(n46807) );
  XOR U46982 ( .A(n46813), .B(n46814), .Z(n46716) );
  ANDN U46983 ( .B(n46815), .A(n46816), .Z(n46813) );
  AND U46984 ( .A(b[5]), .B(a[12]), .Z(n46812) );
  XOR U46985 ( .A(n46818), .B(n46819), .Z(n46721) );
  ANDN U46986 ( .B(n46820), .A(n46821), .Z(n46818) );
  AND U46987 ( .A(b[4]), .B(a[13]), .Z(n46817) );
  XOR U46988 ( .A(n46823), .B(n46824), .Z(n46726) );
  ANDN U46989 ( .B(n46738), .A(n46739), .Z(n46823) );
  AND U46990 ( .A(b[2]), .B(a[14]), .Z(n46825) );
  XNOR U46991 ( .A(n46820), .B(n46824), .Z(n46826) );
  XOR U46992 ( .A(n46827), .B(n46828), .Z(n46824) );
  OR U46993 ( .A(n46741), .B(n46742), .Z(n46828) );
  XNOR U46994 ( .A(n46830), .B(n46831), .Z(n46829) );
  XOR U46995 ( .A(n46830), .B(n46833), .Z(n46741) );
  NAND U46996 ( .A(b[1]), .B(a[14]), .Z(n46833) );
  IV U46997 ( .A(n46827), .Z(n46830) );
  NANDN U46998 ( .A(n189), .B(n190), .Z(n46827) );
  XOR U46999 ( .A(n46834), .B(n46835), .Z(n190) );
  NAND U47000 ( .A(a[14]), .B(b[0]), .Z(n189) );
  XNOR U47001 ( .A(n46815), .B(n46819), .Z(n46836) );
  XNOR U47002 ( .A(n46810), .B(n46814), .Z(n46837) );
  XNOR U47003 ( .A(n46805), .B(n46809), .Z(n46838) );
  XNOR U47004 ( .A(n46800), .B(n46804), .Z(n46839) );
  XNOR U47005 ( .A(n46795), .B(n46799), .Z(n46840) );
  XNOR U47006 ( .A(n46790), .B(n46794), .Z(n46841) );
  XNOR U47007 ( .A(n46785), .B(n46789), .Z(n46842) );
  XNOR U47008 ( .A(n46780), .B(n46784), .Z(n46843) );
  XNOR U47009 ( .A(n46775), .B(n46779), .Z(n46844) );
  XNOR U47010 ( .A(n46770), .B(n46774), .Z(n46845) );
  XNOR U47011 ( .A(n46765), .B(n46769), .Z(n46846) );
  XNOR U47012 ( .A(n46760), .B(n46764), .Z(n46847) );
  XOR U47013 ( .A(n46848), .B(n46759), .Z(n46760) );
  AND U47014 ( .A(a[0]), .B(b[16]), .Z(n46848) );
  XNOR U47015 ( .A(n46849), .B(n46759), .Z(n46761) );
  XNOR U47016 ( .A(n46850), .B(n46851), .Z(n46759) );
  ANDN U47017 ( .B(n46852), .A(n46853), .Z(n46850) );
  AND U47018 ( .A(a[1]), .B(b[15]), .Z(n46849) );
  XOR U47019 ( .A(n46855), .B(n46856), .Z(n46764) );
  ANDN U47020 ( .B(n46857), .A(n46858), .Z(n46855) );
  AND U47021 ( .A(a[2]), .B(b[14]), .Z(n46854) );
  XOR U47022 ( .A(n46860), .B(n46861), .Z(n46769) );
  ANDN U47023 ( .B(n46862), .A(n46863), .Z(n46860) );
  AND U47024 ( .A(a[3]), .B(b[13]), .Z(n46859) );
  XOR U47025 ( .A(n46865), .B(n46866), .Z(n46774) );
  ANDN U47026 ( .B(n46867), .A(n46868), .Z(n46865) );
  AND U47027 ( .A(a[4]), .B(b[12]), .Z(n46864) );
  XOR U47028 ( .A(n46870), .B(n46871), .Z(n46779) );
  ANDN U47029 ( .B(n46872), .A(n46873), .Z(n46870) );
  AND U47030 ( .A(a[5]), .B(b[11]), .Z(n46869) );
  XOR U47031 ( .A(n46875), .B(n46876), .Z(n46784) );
  ANDN U47032 ( .B(n46877), .A(n46878), .Z(n46875) );
  AND U47033 ( .A(a[6]), .B(b[10]), .Z(n46874) );
  XOR U47034 ( .A(n46880), .B(n46881), .Z(n46789) );
  ANDN U47035 ( .B(n46882), .A(n46883), .Z(n46880) );
  AND U47036 ( .A(a[7]), .B(b[9]), .Z(n46879) );
  XOR U47037 ( .A(n46885), .B(n46886), .Z(n46794) );
  ANDN U47038 ( .B(n46887), .A(n46888), .Z(n46885) );
  AND U47039 ( .A(a[8]), .B(b[8]), .Z(n46884) );
  XOR U47040 ( .A(n46890), .B(n46891), .Z(n46799) );
  ANDN U47041 ( .B(n46892), .A(n46893), .Z(n46890) );
  AND U47042 ( .A(a[9]), .B(b[7]), .Z(n46889) );
  XOR U47043 ( .A(n46895), .B(n46896), .Z(n46804) );
  ANDN U47044 ( .B(n46897), .A(n46898), .Z(n46895) );
  AND U47045 ( .A(b[6]), .B(a[10]), .Z(n46894) );
  XOR U47046 ( .A(n46900), .B(n46901), .Z(n46809) );
  ANDN U47047 ( .B(n46902), .A(n46903), .Z(n46900) );
  AND U47048 ( .A(b[5]), .B(a[11]), .Z(n46899) );
  XOR U47049 ( .A(n46905), .B(n46906), .Z(n46814) );
  ANDN U47050 ( .B(n46907), .A(n46908), .Z(n46905) );
  AND U47051 ( .A(b[4]), .B(a[12]), .Z(n46904) );
  XOR U47052 ( .A(n46910), .B(n46911), .Z(n46819) );
  ANDN U47053 ( .B(n46831), .A(n46832), .Z(n46910) );
  AND U47054 ( .A(b[2]), .B(a[13]), .Z(n46912) );
  XNOR U47055 ( .A(n46907), .B(n46911), .Z(n46913) );
  XOR U47056 ( .A(n46914), .B(n46915), .Z(n46911) );
  OR U47057 ( .A(n46834), .B(n46835), .Z(n46915) );
  XNOR U47058 ( .A(n46917), .B(n46918), .Z(n46916) );
  XOR U47059 ( .A(n46917), .B(n46920), .Z(n46834) );
  NAND U47060 ( .A(b[1]), .B(a[13]), .Z(n46920) );
  IV U47061 ( .A(n46914), .Z(n46917) );
  NANDN U47062 ( .A(n191), .B(n192), .Z(n46914) );
  XOR U47063 ( .A(n46921), .B(n46922), .Z(n192) );
  NAND U47064 ( .A(a[13]), .B(b[0]), .Z(n191) );
  XNOR U47065 ( .A(n46902), .B(n46906), .Z(n46923) );
  XNOR U47066 ( .A(n46897), .B(n46901), .Z(n46924) );
  XNOR U47067 ( .A(n46892), .B(n46896), .Z(n46925) );
  XNOR U47068 ( .A(n46887), .B(n46891), .Z(n46926) );
  XNOR U47069 ( .A(n46882), .B(n46886), .Z(n46927) );
  XNOR U47070 ( .A(n46877), .B(n46881), .Z(n46928) );
  XNOR U47071 ( .A(n46872), .B(n46876), .Z(n46929) );
  XNOR U47072 ( .A(n46867), .B(n46871), .Z(n46930) );
  XNOR U47073 ( .A(n46862), .B(n46866), .Z(n46931) );
  XNOR U47074 ( .A(n46857), .B(n46861), .Z(n46932) );
  XNOR U47075 ( .A(n46852), .B(n46856), .Z(n46933) );
  XNOR U47076 ( .A(n46934), .B(n46851), .Z(n46852) );
  AND U47077 ( .A(a[0]), .B(b[15]), .Z(n46934) );
  XOR U47078 ( .A(n46935), .B(n46851), .Z(n46853) );
  XNOR U47079 ( .A(n46936), .B(n46937), .Z(n46851) );
  ANDN U47080 ( .B(n46938), .A(n46939), .Z(n46936) );
  AND U47081 ( .A(a[1]), .B(b[14]), .Z(n46935) );
  XOR U47082 ( .A(n46941), .B(n46942), .Z(n46856) );
  ANDN U47083 ( .B(n46943), .A(n46944), .Z(n46941) );
  AND U47084 ( .A(a[2]), .B(b[13]), .Z(n46940) );
  XOR U47085 ( .A(n46946), .B(n46947), .Z(n46861) );
  ANDN U47086 ( .B(n46948), .A(n46949), .Z(n46946) );
  AND U47087 ( .A(a[3]), .B(b[12]), .Z(n46945) );
  XOR U47088 ( .A(n46951), .B(n46952), .Z(n46866) );
  ANDN U47089 ( .B(n46953), .A(n46954), .Z(n46951) );
  AND U47090 ( .A(a[4]), .B(b[11]), .Z(n46950) );
  XOR U47091 ( .A(n46956), .B(n46957), .Z(n46871) );
  ANDN U47092 ( .B(n46958), .A(n46959), .Z(n46956) );
  AND U47093 ( .A(a[5]), .B(b[10]), .Z(n46955) );
  XOR U47094 ( .A(n46961), .B(n46962), .Z(n46876) );
  ANDN U47095 ( .B(n46963), .A(n46964), .Z(n46961) );
  AND U47096 ( .A(a[6]), .B(b[9]), .Z(n46960) );
  XOR U47097 ( .A(n46966), .B(n46967), .Z(n46881) );
  ANDN U47098 ( .B(n46968), .A(n46969), .Z(n46966) );
  AND U47099 ( .A(a[7]), .B(b[8]), .Z(n46965) );
  XOR U47100 ( .A(n46971), .B(n46972), .Z(n46886) );
  ANDN U47101 ( .B(n46973), .A(n46974), .Z(n46971) );
  AND U47102 ( .A(a[8]), .B(b[7]), .Z(n46970) );
  XOR U47103 ( .A(n46976), .B(n46977), .Z(n46891) );
  ANDN U47104 ( .B(n46978), .A(n46979), .Z(n46976) );
  AND U47105 ( .A(a[9]), .B(b[6]), .Z(n46975) );
  XOR U47106 ( .A(n46981), .B(n46982), .Z(n46896) );
  ANDN U47107 ( .B(n46983), .A(n46984), .Z(n46981) );
  AND U47108 ( .A(b[5]), .B(a[10]), .Z(n46980) );
  XOR U47109 ( .A(n46986), .B(n46987), .Z(n46901) );
  ANDN U47110 ( .B(n46988), .A(n46989), .Z(n46986) );
  AND U47111 ( .A(b[4]), .B(a[11]), .Z(n46985) );
  XOR U47112 ( .A(n46991), .B(n46992), .Z(n46906) );
  ANDN U47113 ( .B(n46918), .A(n46919), .Z(n46991) );
  AND U47114 ( .A(b[2]), .B(a[12]), .Z(n46993) );
  XNOR U47115 ( .A(n46988), .B(n46992), .Z(n46994) );
  XOR U47116 ( .A(n46995), .B(n46996), .Z(n46992) );
  OR U47117 ( .A(n46921), .B(n46922), .Z(n46996) );
  XNOR U47118 ( .A(n46998), .B(n46999), .Z(n46997) );
  XOR U47119 ( .A(n46998), .B(n47001), .Z(n46921) );
  NAND U47120 ( .A(b[1]), .B(a[12]), .Z(n47001) );
  IV U47121 ( .A(n46995), .Z(n46998) );
  NANDN U47122 ( .A(n193), .B(n194), .Z(n46995) );
  XOR U47123 ( .A(n47002), .B(n47003), .Z(n194) );
  NAND U47124 ( .A(a[12]), .B(b[0]), .Z(n193) );
  XNOR U47125 ( .A(n46983), .B(n46987), .Z(n47004) );
  XNOR U47126 ( .A(n46978), .B(n46982), .Z(n47005) );
  XNOR U47127 ( .A(n46973), .B(n46977), .Z(n47006) );
  XNOR U47128 ( .A(n46968), .B(n46972), .Z(n47007) );
  XNOR U47129 ( .A(n46963), .B(n46967), .Z(n47008) );
  XNOR U47130 ( .A(n46958), .B(n46962), .Z(n47009) );
  XNOR U47131 ( .A(n46953), .B(n46957), .Z(n47010) );
  XNOR U47132 ( .A(n46948), .B(n46952), .Z(n47011) );
  XNOR U47133 ( .A(n46943), .B(n46947), .Z(n47012) );
  XNOR U47134 ( .A(n46938), .B(n46942), .Z(n47013) );
  XOR U47135 ( .A(n47014), .B(n46937), .Z(n46938) );
  AND U47136 ( .A(a[0]), .B(b[14]), .Z(n47014) );
  XNOR U47137 ( .A(n47015), .B(n46937), .Z(n46939) );
  XNOR U47138 ( .A(n47016), .B(n47017), .Z(n46937) );
  ANDN U47139 ( .B(n47018), .A(n47019), .Z(n47016) );
  AND U47140 ( .A(a[1]), .B(b[13]), .Z(n47015) );
  XOR U47141 ( .A(n47021), .B(n47022), .Z(n46942) );
  ANDN U47142 ( .B(n47023), .A(n47024), .Z(n47021) );
  AND U47143 ( .A(a[2]), .B(b[12]), .Z(n47020) );
  XOR U47144 ( .A(n47026), .B(n47027), .Z(n46947) );
  ANDN U47145 ( .B(n47028), .A(n47029), .Z(n47026) );
  AND U47146 ( .A(a[3]), .B(b[11]), .Z(n47025) );
  XOR U47147 ( .A(n47031), .B(n47032), .Z(n46952) );
  ANDN U47148 ( .B(n47033), .A(n47034), .Z(n47031) );
  AND U47149 ( .A(a[4]), .B(b[10]), .Z(n47030) );
  XOR U47150 ( .A(n47036), .B(n47037), .Z(n46957) );
  ANDN U47151 ( .B(n47038), .A(n47039), .Z(n47036) );
  AND U47152 ( .A(a[5]), .B(b[9]), .Z(n47035) );
  XOR U47153 ( .A(n47041), .B(n47042), .Z(n46962) );
  ANDN U47154 ( .B(n47043), .A(n47044), .Z(n47041) );
  AND U47155 ( .A(a[6]), .B(b[8]), .Z(n47040) );
  XOR U47156 ( .A(n47046), .B(n47047), .Z(n46967) );
  ANDN U47157 ( .B(n47048), .A(n47049), .Z(n47046) );
  AND U47158 ( .A(a[7]), .B(b[7]), .Z(n47045) );
  XOR U47159 ( .A(n47051), .B(n47052), .Z(n46972) );
  ANDN U47160 ( .B(n47053), .A(n47054), .Z(n47051) );
  AND U47161 ( .A(a[8]), .B(b[6]), .Z(n47050) );
  XOR U47162 ( .A(n47056), .B(n47057), .Z(n46977) );
  ANDN U47163 ( .B(n47058), .A(n47059), .Z(n47056) );
  AND U47164 ( .A(a[9]), .B(b[5]), .Z(n47055) );
  XOR U47165 ( .A(n47061), .B(n47062), .Z(n46982) );
  ANDN U47166 ( .B(n47063), .A(n47064), .Z(n47061) );
  AND U47167 ( .A(b[4]), .B(a[10]), .Z(n47060) );
  XOR U47168 ( .A(n47066), .B(n47067), .Z(n46987) );
  ANDN U47169 ( .B(n46999), .A(n47000), .Z(n47066) );
  AND U47170 ( .A(b[2]), .B(a[11]), .Z(n47068) );
  XNOR U47171 ( .A(n47063), .B(n47067), .Z(n47069) );
  XOR U47172 ( .A(n47070), .B(n47071), .Z(n47067) );
  OR U47173 ( .A(n47002), .B(n47003), .Z(n47071) );
  XNOR U47174 ( .A(n47073), .B(n47074), .Z(n47072) );
  XOR U47175 ( .A(n47073), .B(n47076), .Z(n47002) );
  NAND U47176 ( .A(b[1]), .B(a[11]), .Z(n47076) );
  IV U47177 ( .A(n47070), .Z(n47073) );
  NANDN U47178 ( .A(n5595), .B(n5596), .Z(n47070) );
  XOR U47179 ( .A(n47077), .B(n47078), .Z(n5596) );
  NAND U47180 ( .A(a[11]), .B(b[0]), .Z(n5595) );
  XNOR U47181 ( .A(n47058), .B(n47062), .Z(n47079) );
  XNOR U47182 ( .A(n47053), .B(n47057), .Z(n47080) );
  XNOR U47183 ( .A(n47048), .B(n47052), .Z(n47081) );
  XNOR U47184 ( .A(n47043), .B(n47047), .Z(n47082) );
  XNOR U47185 ( .A(n47038), .B(n47042), .Z(n47083) );
  XNOR U47186 ( .A(n47033), .B(n47037), .Z(n47084) );
  XNOR U47187 ( .A(n47028), .B(n47032), .Z(n47085) );
  XNOR U47188 ( .A(n47023), .B(n47027), .Z(n47086) );
  XNOR U47189 ( .A(n47018), .B(n47022), .Z(n47087) );
  XNOR U47190 ( .A(n47088), .B(n47017), .Z(n47018) );
  AND U47191 ( .A(a[0]), .B(b[13]), .Z(n47088) );
  XOR U47192 ( .A(n47089), .B(n47017), .Z(n47019) );
  XNOR U47193 ( .A(n47090), .B(n47091), .Z(n47017) );
  ANDN U47194 ( .B(n47092), .A(n47093), .Z(n47090) );
  AND U47195 ( .A(a[1]), .B(b[12]), .Z(n47089) );
  XOR U47196 ( .A(n47095), .B(n47096), .Z(n47022) );
  ANDN U47197 ( .B(n47097), .A(n47098), .Z(n47095) );
  AND U47198 ( .A(a[2]), .B(b[11]), .Z(n47094) );
  XOR U47199 ( .A(n47100), .B(n47101), .Z(n47027) );
  ANDN U47200 ( .B(n47102), .A(n47103), .Z(n47100) );
  AND U47201 ( .A(a[3]), .B(b[10]), .Z(n47099) );
  XOR U47202 ( .A(n47105), .B(n47106), .Z(n47032) );
  ANDN U47203 ( .B(n47107), .A(n47108), .Z(n47105) );
  AND U47204 ( .A(a[4]), .B(b[9]), .Z(n47104) );
  XOR U47205 ( .A(n47110), .B(n47111), .Z(n47037) );
  ANDN U47206 ( .B(n47112), .A(n47113), .Z(n47110) );
  AND U47207 ( .A(a[5]), .B(b[8]), .Z(n47109) );
  XOR U47208 ( .A(n47115), .B(n47116), .Z(n47042) );
  ANDN U47209 ( .B(n47117), .A(n47118), .Z(n47115) );
  AND U47210 ( .A(a[6]), .B(b[7]), .Z(n47114) );
  XOR U47211 ( .A(n47120), .B(n47121), .Z(n47047) );
  ANDN U47212 ( .B(n47122), .A(n47123), .Z(n47120) );
  AND U47213 ( .A(a[7]), .B(b[6]), .Z(n47119) );
  XOR U47214 ( .A(n47125), .B(n47126), .Z(n47052) );
  ANDN U47215 ( .B(n47127), .A(n47128), .Z(n47125) );
  AND U47216 ( .A(a[8]), .B(b[5]), .Z(n47124) );
  XOR U47217 ( .A(n47130), .B(n47131), .Z(n47057) );
  ANDN U47218 ( .B(n47132), .A(n47133), .Z(n47130) );
  AND U47219 ( .A(a[9]), .B(b[4]), .Z(n47129) );
  XOR U47220 ( .A(n47135), .B(n47136), .Z(n47062) );
  ANDN U47221 ( .B(n47074), .A(n47075), .Z(n47135) );
  AND U47222 ( .A(b[2]), .B(a[10]), .Z(n47137) );
  XNOR U47223 ( .A(n47132), .B(n47136), .Z(n47138) );
  XOR U47224 ( .A(n47139), .B(n47140), .Z(n47136) );
  OR U47225 ( .A(n47077), .B(n47078), .Z(n47140) );
  XNOR U47226 ( .A(n47142), .B(n47143), .Z(n47141) );
  XOR U47227 ( .A(n47142), .B(n47145), .Z(n47077) );
  NAND U47228 ( .A(b[1]), .B(a[10]), .Z(n47145) );
  IV U47229 ( .A(n47139), .Z(n47142) );
  NANDN U47230 ( .A(n12387), .B(n12388), .Z(n47139) );
  XOR U47231 ( .A(n47146), .B(n47147), .Z(n12388) );
  NAND U47232 ( .A(a[10]), .B(b[0]), .Z(n12387) );
  XNOR U47233 ( .A(n47127), .B(n47131), .Z(n47148) );
  XNOR U47234 ( .A(n47122), .B(n47126), .Z(n47149) );
  XNOR U47235 ( .A(n47117), .B(n47121), .Z(n47150) );
  XNOR U47236 ( .A(n47112), .B(n47116), .Z(n47151) );
  XNOR U47237 ( .A(n47107), .B(n47111), .Z(n47152) );
  XNOR U47238 ( .A(n47102), .B(n47106), .Z(n47153) );
  XNOR U47239 ( .A(n47097), .B(n47101), .Z(n47154) );
  XNOR U47240 ( .A(n47092), .B(n47096), .Z(n47155) );
  XOR U47241 ( .A(n47156), .B(n47091), .Z(n47092) );
  AND U47242 ( .A(a[0]), .B(b[12]), .Z(n47156) );
  XNOR U47243 ( .A(n47157), .B(n47091), .Z(n47093) );
  XNOR U47244 ( .A(n47158), .B(n47159), .Z(n47091) );
  ANDN U47245 ( .B(n47160), .A(n47161), .Z(n47158) );
  AND U47246 ( .A(a[1]), .B(b[11]), .Z(n47157) );
  XOR U47247 ( .A(n47163), .B(n47164), .Z(n47096) );
  ANDN U47248 ( .B(n47165), .A(n47166), .Z(n47163) );
  AND U47249 ( .A(a[2]), .B(b[10]), .Z(n47162) );
  XOR U47250 ( .A(n47168), .B(n47169), .Z(n47101) );
  ANDN U47251 ( .B(n47170), .A(n47171), .Z(n47168) );
  AND U47252 ( .A(a[3]), .B(b[9]), .Z(n47167) );
  XOR U47253 ( .A(n47173), .B(n47174), .Z(n47106) );
  ANDN U47254 ( .B(n47175), .A(n47176), .Z(n47173) );
  AND U47255 ( .A(a[4]), .B(b[8]), .Z(n47172) );
  XOR U47256 ( .A(n47178), .B(n47179), .Z(n47111) );
  ANDN U47257 ( .B(n47180), .A(n47181), .Z(n47178) );
  AND U47258 ( .A(a[5]), .B(b[7]), .Z(n47177) );
  XOR U47259 ( .A(n47183), .B(n47184), .Z(n47116) );
  ANDN U47260 ( .B(n47185), .A(n47186), .Z(n47183) );
  AND U47261 ( .A(a[6]), .B(b[6]), .Z(n47182) );
  XOR U47262 ( .A(n47188), .B(n47189), .Z(n47121) );
  ANDN U47263 ( .B(n47190), .A(n47191), .Z(n47188) );
  AND U47264 ( .A(a[7]), .B(b[5]), .Z(n47187) );
  XOR U47265 ( .A(n47193), .B(n47194), .Z(n47126) );
  ANDN U47266 ( .B(n47195), .A(n47196), .Z(n47193) );
  AND U47267 ( .A(a[8]), .B(b[4]), .Z(n47192) );
  XOR U47268 ( .A(n47198), .B(n47199), .Z(n47131) );
  ANDN U47269 ( .B(n47143), .A(n47144), .Z(n47198) );
  AND U47270 ( .A(a[9]), .B(b[2]), .Z(n47200) );
  XNOR U47271 ( .A(n47195), .B(n47199), .Z(n47201) );
  XOR U47272 ( .A(n47202), .B(n47203), .Z(n47199) );
  OR U47273 ( .A(n47146), .B(n47147), .Z(n47203) );
  XOR U47274 ( .A(n47202), .B(n47205), .Z(n47204) );
  XNOR U47275 ( .A(n47202), .B(n47207), .Z(n47146) );
  NAND U47276 ( .A(a[9]), .B(b[1]), .Z(n47207) );
  OR U47277 ( .A(n1), .B(n2), .Z(n47202) );
  XOR U47278 ( .A(n47208), .B(n47209), .Z(n2) );
  NAND U47279 ( .A(b[0]), .B(a[9]), .Z(n1) );
  XNOR U47280 ( .A(n47190), .B(n47194), .Z(n47210) );
  XNOR U47281 ( .A(n47185), .B(n47189), .Z(n47211) );
  XNOR U47282 ( .A(n47180), .B(n47184), .Z(n47212) );
  XNOR U47283 ( .A(n47175), .B(n47179), .Z(n47213) );
  XNOR U47284 ( .A(n47170), .B(n47174), .Z(n47214) );
  XNOR U47285 ( .A(n47165), .B(n47169), .Z(n47215) );
  XNOR U47286 ( .A(n47160), .B(n47164), .Z(n47216) );
  XNOR U47287 ( .A(n47217), .B(n47159), .Z(n47160) );
  AND U47288 ( .A(a[0]), .B(b[11]), .Z(n47217) );
  XOR U47289 ( .A(n47218), .B(n47159), .Z(n47161) );
  XNOR U47290 ( .A(n47219), .B(n47220), .Z(n47159) );
  ANDN U47291 ( .B(n47221), .A(n47222), .Z(n47219) );
  AND U47292 ( .A(a[1]), .B(b[10]), .Z(n47218) );
  XOR U47293 ( .A(n47224), .B(n47225), .Z(n47164) );
  ANDN U47294 ( .B(n47226), .A(n47227), .Z(n47224) );
  AND U47295 ( .A(a[2]), .B(b[9]), .Z(n47223) );
  XOR U47296 ( .A(n47229), .B(n47230), .Z(n47169) );
  ANDN U47297 ( .B(n47231), .A(n47232), .Z(n47229) );
  AND U47298 ( .A(a[3]), .B(b[8]), .Z(n47228) );
  XOR U47299 ( .A(n47234), .B(n47235), .Z(n47174) );
  ANDN U47300 ( .B(n47236), .A(n47237), .Z(n47234) );
  AND U47301 ( .A(a[4]), .B(b[7]), .Z(n47233) );
  XOR U47302 ( .A(n47239), .B(n47240), .Z(n47179) );
  ANDN U47303 ( .B(n47241), .A(n47242), .Z(n47239) );
  AND U47304 ( .A(a[5]), .B(b[6]), .Z(n47238) );
  XOR U47305 ( .A(n47244), .B(n47245), .Z(n47184) );
  ANDN U47306 ( .B(n47246), .A(n47247), .Z(n47244) );
  AND U47307 ( .A(a[6]), .B(b[5]), .Z(n47243) );
  XOR U47308 ( .A(n47249), .B(n47250), .Z(n47189) );
  ANDN U47309 ( .B(n47251), .A(n47252), .Z(n47249) );
  AND U47310 ( .A(a[7]), .B(b[4]), .Z(n47248) );
  XOR U47311 ( .A(n47254), .B(n47255), .Z(n47194) );
  ANDN U47312 ( .B(n47205), .A(n47206), .Z(n47254) );
  AND U47313 ( .A(a[8]), .B(b[2]), .Z(n47256) );
  XNOR U47314 ( .A(n47251), .B(n47255), .Z(n47257) );
  XOR U47315 ( .A(n47258), .B(n47259), .Z(n47255) );
  NANDN U47316 ( .A(n47209), .B(n47208), .Z(n47259) );
  XOR U47317 ( .A(n47258), .B(n47260), .Z(n47208) );
  NAND U47318 ( .A(a[8]), .B(b[1]), .Z(n47260) );
  XNOR U47319 ( .A(n47262), .B(n47263), .Z(n47261) );
  IV U47320 ( .A(n47258), .Z(n47262) );
  NANDN U47321 ( .A(n23), .B(n24), .Z(n47258) );
  XOR U47322 ( .A(n47265), .B(n47266), .Z(n24) );
  NAND U47323 ( .A(a[8]), .B(b[0]), .Z(n23) );
  XNOR U47324 ( .A(n47246), .B(n47250), .Z(n47267) );
  XNOR U47325 ( .A(n47241), .B(n47245), .Z(n47268) );
  XNOR U47326 ( .A(n47236), .B(n47240), .Z(n47269) );
  XNOR U47327 ( .A(n47231), .B(n47235), .Z(n47270) );
  XNOR U47328 ( .A(n47226), .B(n47230), .Z(n47271) );
  XNOR U47329 ( .A(n47221), .B(n47225), .Z(n47272) );
  XOR U47330 ( .A(n47273), .B(n47220), .Z(n47221) );
  AND U47331 ( .A(a[0]), .B(b[10]), .Z(n47273) );
  XNOR U47332 ( .A(n47274), .B(n47220), .Z(n47222) );
  XNOR U47333 ( .A(n47275), .B(n47276), .Z(n47220) );
  ANDN U47334 ( .B(n47277), .A(n47278), .Z(n47275) );
  AND U47335 ( .A(a[1]), .B(b[9]), .Z(n47274) );
  XOR U47336 ( .A(n47280), .B(n47281), .Z(n47225) );
  ANDN U47337 ( .B(n47282), .A(n47283), .Z(n47280) );
  AND U47338 ( .A(a[2]), .B(b[8]), .Z(n47279) );
  XOR U47339 ( .A(n47285), .B(n47286), .Z(n47230) );
  ANDN U47340 ( .B(n47287), .A(n47288), .Z(n47285) );
  AND U47341 ( .A(a[3]), .B(b[7]), .Z(n47284) );
  XOR U47342 ( .A(n47290), .B(n47291), .Z(n47235) );
  ANDN U47343 ( .B(n47292), .A(n47293), .Z(n47290) );
  AND U47344 ( .A(a[4]), .B(b[6]), .Z(n47289) );
  XOR U47345 ( .A(n47295), .B(n47296), .Z(n47240) );
  ANDN U47346 ( .B(n47297), .A(n47298), .Z(n47295) );
  AND U47347 ( .A(a[5]), .B(b[5]), .Z(n47294) );
  XOR U47348 ( .A(n47300), .B(n47301), .Z(n47245) );
  ANDN U47349 ( .B(n47302), .A(n47303), .Z(n47300) );
  AND U47350 ( .A(a[6]), .B(b[4]), .Z(n47299) );
  XOR U47351 ( .A(n47305), .B(n47306), .Z(n47250) );
  ANDN U47352 ( .B(n47263), .A(n47264), .Z(n47305) );
  AND U47353 ( .A(a[7]), .B(b[2]), .Z(n47307) );
  XNOR U47354 ( .A(n47302), .B(n47306), .Z(n47308) );
  XOR U47355 ( .A(n47309), .B(n47310), .Z(n47306) );
  OR U47356 ( .A(n47265), .B(n47266), .Z(n47310) );
  XNOR U47357 ( .A(n47312), .B(n47313), .Z(n47311) );
  XOR U47358 ( .A(n47312), .B(n47315), .Z(n47265) );
  NAND U47359 ( .A(a[7]), .B(b[1]), .Z(n47315) );
  IV U47360 ( .A(n47309), .Z(n47312) );
  NANDN U47361 ( .A(n45), .B(n46), .Z(n47309) );
  XOR U47362 ( .A(n47316), .B(n47317), .Z(n46) );
  NAND U47363 ( .A(a[7]), .B(b[0]), .Z(n45) );
  XNOR U47364 ( .A(n47297), .B(n47301), .Z(n47318) );
  XNOR U47365 ( .A(n47292), .B(n47296), .Z(n47319) );
  XNOR U47366 ( .A(n47287), .B(n47291), .Z(n47320) );
  XNOR U47367 ( .A(n47282), .B(n47286), .Z(n47321) );
  XNOR U47368 ( .A(n47277), .B(n47281), .Z(n47322) );
  XNOR U47369 ( .A(n47323), .B(n47276), .Z(n47277) );
  AND U47370 ( .A(a[0]), .B(b[9]), .Z(n47323) );
  XOR U47371 ( .A(n47324), .B(n47276), .Z(n47278) );
  XNOR U47372 ( .A(n47325), .B(n47326), .Z(n47276) );
  ANDN U47373 ( .B(n47327), .A(n47328), .Z(n47325) );
  AND U47374 ( .A(a[1]), .B(b[8]), .Z(n47324) );
  XOR U47375 ( .A(n47330), .B(n47331), .Z(n47281) );
  ANDN U47376 ( .B(n47332), .A(n47333), .Z(n47330) );
  AND U47377 ( .A(a[2]), .B(b[7]), .Z(n47329) );
  XOR U47378 ( .A(n47335), .B(n47336), .Z(n47286) );
  ANDN U47379 ( .B(n47337), .A(n47338), .Z(n47335) );
  AND U47380 ( .A(a[3]), .B(b[6]), .Z(n47334) );
  XOR U47381 ( .A(n47340), .B(n47341), .Z(n47291) );
  ANDN U47382 ( .B(n47342), .A(n47343), .Z(n47340) );
  AND U47383 ( .A(a[4]), .B(b[5]), .Z(n47339) );
  XOR U47384 ( .A(n47345), .B(n47346), .Z(n47296) );
  ANDN U47385 ( .B(n47347), .A(n47348), .Z(n47345) );
  AND U47386 ( .A(a[5]), .B(b[4]), .Z(n47344) );
  XOR U47387 ( .A(n47350), .B(n47351), .Z(n47301) );
  ANDN U47388 ( .B(n47313), .A(n47314), .Z(n47350) );
  AND U47389 ( .A(a[6]), .B(b[2]), .Z(n47352) );
  XNOR U47390 ( .A(n47347), .B(n47351), .Z(n47353) );
  XOR U47391 ( .A(n47354), .B(n47355), .Z(n47351) );
  OR U47392 ( .A(n47316), .B(n47317), .Z(n47355) );
  XNOR U47393 ( .A(n47357), .B(n47358), .Z(n47356) );
  XOR U47394 ( .A(n47357), .B(n47360), .Z(n47316) );
  NAND U47395 ( .A(a[6]), .B(b[1]), .Z(n47360) );
  IV U47396 ( .A(n47354), .Z(n47357) );
  NANDN U47397 ( .A(n67), .B(n68), .Z(n47354) );
  XOR U47398 ( .A(n47361), .B(n47362), .Z(n68) );
  NAND U47399 ( .A(a[6]), .B(b[0]), .Z(n67) );
  XNOR U47400 ( .A(n47342), .B(n47346), .Z(n47363) );
  XNOR U47401 ( .A(n47337), .B(n47341), .Z(n47364) );
  XNOR U47402 ( .A(n47332), .B(n47336), .Z(n47365) );
  XNOR U47403 ( .A(n47327), .B(n47331), .Z(n47366) );
  XOR U47404 ( .A(n47367), .B(n47326), .Z(n47327) );
  AND U47405 ( .A(a[0]), .B(b[8]), .Z(n47367) );
  XNOR U47406 ( .A(n47368), .B(n47326), .Z(n47328) );
  XNOR U47407 ( .A(n47369), .B(n47370), .Z(n47326) );
  ANDN U47408 ( .B(n47371), .A(n47372), .Z(n47369) );
  AND U47409 ( .A(a[1]), .B(b[7]), .Z(n47368) );
  XOR U47410 ( .A(n47374), .B(n47375), .Z(n47331) );
  ANDN U47411 ( .B(n47376), .A(n47377), .Z(n47374) );
  AND U47412 ( .A(a[2]), .B(b[6]), .Z(n47373) );
  XOR U47413 ( .A(n47379), .B(n47380), .Z(n47336) );
  ANDN U47414 ( .B(n47381), .A(n47382), .Z(n47379) );
  AND U47415 ( .A(a[3]), .B(b[5]), .Z(n47378) );
  XOR U47416 ( .A(n47384), .B(n47385), .Z(n47341) );
  ANDN U47417 ( .B(n47386), .A(n47387), .Z(n47384) );
  AND U47418 ( .A(a[4]), .B(b[4]), .Z(n47383) );
  XOR U47419 ( .A(n47389), .B(n47390), .Z(n47346) );
  ANDN U47420 ( .B(n47358), .A(n47359), .Z(n47389) );
  AND U47421 ( .A(a[5]), .B(b[2]), .Z(n47391) );
  XNOR U47422 ( .A(n47386), .B(n47390), .Z(n47392) );
  XOR U47423 ( .A(n47393), .B(n47394), .Z(n47390) );
  OR U47424 ( .A(n47361), .B(n47362), .Z(n47394) );
  XNOR U47425 ( .A(n47396), .B(n47397), .Z(n47395) );
  XOR U47426 ( .A(n47396), .B(n47399), .Z(n47361) );
  NAND U47427 ( .A(a[5]), .B(b[1]), .Z(n47399) );
  IV U47428 ( .A(n47393), .Z(n47396) );
  NANDN U47429 ( .A(n89), .B(n90), .Z(n47393) );
  XOR U47430 ( .A(n47400), .B(n47401), .Z(n90) );
  NAND U47431 ( .A(a[5]), .B(b[0]), .Z(n89) );
  XNOR U47432 ( .A(n47381), .B(n47385), .Z(n47402) );
  XNOR U47433 ( .A(n47376), .B(n47380), .Z(n47403) );
  XNOR U47434 ( .A(n47371), .B(n47375), .Z(n47404) );
  XNOR U47435 ( .A(n47405), .B(n47370), .Z(n47371) );
  AND U47436 ( .A(a[0]), .B(b[7]), .Z(n47405) );
  XOR U47437 ( .A(n47406), .B(n47370), .Z(n47372) );
  XNOR U47438 ( .A(n47407), .B(n47408), .Z(n47370) );
  ANDN U47439 ( .B(n47409), .A(n47410), .Z(n47407) );
  AND U47440 ( .A(a[1]), .B(b[6]), .Z(n47406) );
  XOR U47441 ( .A(n47412), .B(n47413), .Z(n47375) );
  ANDN U47442 ( .B(n47414), .A(n47415), .Z(n47412) );
  AND U47443 ( .A(a[2]), .B(b[5]), .Z(n47411) );
  XOR U47444 ( .A(n47417), .B(n47418), .Z(n47380) );
  ANDN U47445 ( .B(n47419), .A(n47420), .Z(n47417) );
  AND U47446 ( .A(a[3]), .B(b[4]), .Z(n47416) );
  XOR U47447 ( .A(n47422), .B(n47423), .Z(n47385) );
  ANDN U47448 ( .B(n47397), .A(n47398), .Z(n47422) );
  AND U47449 ( .A(a[4]), .B(b[2]), .Z(n47424) );
  XNOR U47450 ( .A(n47419), .B(n47423), .Z(n47425) );
  XOR U47451 ( .A(n47426), .B(n47427), .Z(n47423) );
  OR U47452 ( .A(n47400), .B(n47401), .Z(n47427) );
  XNOR U47453 ( .A(n47429), .B(n47430), .Z(n47428) );
  XOR U47454 ( .A(n47429), .B(n47432), .Z(n47400) );
  NAND U47455 ( .A(a[4]), .B(b[1]), .Z(n47432) );
  IV U47456 ( .A(n47426), .Z(n47429) );
  NANDN U47457 ( .A(n111), .B(n112), .Z(n47426) );
  XOR U47458 ( .A(n47433), .B(n47434), .Z(n112) );
  NAND U47459 ( .A(a[4]), .B(b[0]), .Z(n111) );
  XNOR U47460 ( .A(n47414), .B(n47418), .Z(n47435) );
  XNOR U47461 ( .A(n47409), .B(n47413), .Z(n47436) );
  XOR U47462 ( .A(n47437), .B(n47408), .Z(n47409) );
  AND U47463 ( .A(a[0]), .B(b[6]), .Z(n47437) );
  XNOR U47464 ( .A(n47438), .B(n47408), .Z(n47410) );
  XNOR U47465 ( .A(n47439), .B(n47440), .Z(n47408) );
  ANDN U47466 ( .B(n47441), .A(n47442), .Z(n47439) );
  AND U47467 ( .A(a[1]), .B(b[5]), .Z(n47438) );
  XOR U47468 ( .A(n47444), .B(n47445), .Z(n47413) );
  ANDN U47469 ( .B(n47446), .A(n47447), .Z(n47444) );
  AND U47470 ( .A(a[2]), .B(b[4]), .Z(n47443) );
  XOR U47471 ( .A(n47449), .B(n47450), .Z(n47418) );
  ANDN U47472 ( .B(n47430), .A(n47431), .Z(n47449) );
  AND U47473 ( .A(a[3]), .B(b[2]), .Z(n47451) );
  XNOR U47474 ( .A(n47446), .B(n47450), .Z(n47452) );
  XOR U47475 ( .A(n47453), .B(n47454), .Z(n47450) );
  OR U47476 ( .A(n47433), .B(n47434), .Z(n47454) );
  XNOR U47477 ( .A(n47456), .B(n47457), .Z(n47455) );
  XOR U47478 ( .A(n47456), .B(n47459), .Z(n47433) );
  NAND U47479 ( .A(a[3]), .B(b[1]), .Z(n47459) );
  IV U47480 ( .A(n47453), .Z(n47456) );
  NANDN U47481 ( .A(n133), .B(n134), .Z(n47453) );
  XOR U47482 ( .A(n47460), .B(n47461), .Z(n134) );
  NAND U47483 ( .A(a[3]), .B(b[0]), .Z(n133) );
  XNOR U47484 ( .A(n47441), .B(n47445), .Z(n47462) );
  XNOR U47485 ( .A(n47463), .B(n47440), .Z(n47441) );
  AND U47486 ( .A(a[0]), .B(b[5]), .Z(n47463) );
  XOR U47487 ( .A(n47464), .B(n47440), .Z(n47442) );
  XNOR U47488 ( .A(n47465), .B(n47466), .Z(n47440) );
  ANDN U47489 ( .B(n47467), .A(n47468), .Z(n47465) );
  AND U47490 ( .A(a[1]), .B(b[4]), .Z(n47464) );
  XOR U47491 ( .A(n47470), .B(n47471), .Z(n47445) );
  ANDN U47492 ( .B(n47457), .A(n47458), .Z(n47470) );
  AND U47493 ( .A(a[2]), .B(b[2]), .Z(n47472) );
  XNOR U47494 ( .A(n47467), .B(n47471), .Z(n47473) );
  XOR U47495 ( .A(n47474), .B(n47475), .Z(n47471) );
  OR U47496 ( .A(n47460), .B(n47461), .Z(n47475) );
  XNOR U47497 ( .A(n47477), .B(n47478), .Z(n47476) );
  XOR U47498 ( .A(n47477), .B(n47480), .Z(n47460) );
  NAND U47499 ( .A(a[2]), .B(b[1]), .Z(n47480) );
  IV U47500 ( .A(n47474), .Z(n47477) );
  NANDN U47501 ( .A(n155), .B(n156), .Z(n47474) );
  XOR U47502 ( .A(n47481), .B(n47482), .Z(n156) );
  NAND U47503 ( .A(a[2]), .B(b[0]), .Z(n155) );
  XOR U47504 ( .A(n47483), .B(n47466), .Z(n47467) );
  AND U47505 ( .A(a[0]), .B(b[4]), .Z(n47483) );
  XNOR U47506 ( .A(n47484), .B(n47466), .Z(n47468) );
  XNOR U47507 ( .A(n47485), .B(n47486), .Z(n47466) );
  ANDN U47508 ( .B(n47478), .A(n47479), .Z(n47485) );
  XOR U47509 ( .A(n47487), .B(n47486), .Z(n47479) );
  AND U47510 ( .A(a[1]), .B(b[2]), .Z(n47487) );
  XNOR U47511 ( .A(n47488), .B(n47486), .Z(n47478) );
  XNOR U47512 ( .A(n47489), .B(n47490), .Z(n47486) );
  OR U47513 ( .A(n47482), .B(n47481), .Z(n47490) );
  XNOR U47514 ( .A(n47489), .B(n47491), .Z(n47481) );
  NAND U47515 ( .A(a[1]), .B(b[1]), .Z(n47491) );
  XNOR U47516 ( .A(n47489), .B(n47492), .Z(n47482) );
  NAND U47517 ( .A(a[0]), .B(b[2]), .Z(n47492) );
  OR U47518 ( .A(n177), .B(n178), .Z(n47489) );
  NAND U47519 ( .A(b[1]), .B(a[0]), .Z(n178) );
  NAND U47520 ( .A(a[1]), .B(b[0]), .Z(n177) );
  AND U47521 ( .A(a[0]), .B(b[3]), .Z(n47488) );
  AND U47522 ( .A(a[1]), .B(b[3]), .Z(n47484) );
  AND U47523 ( .A(a[2]), .B(b[3]), .Z(n47469) );
  AND U47524 ( .A(a[3]), .B(b[3]), .Z(n47448) );
  AND U47525 ( .A(a[4]), .B(b[3]), .Z(n47421) );
  AND U47526 ( .A(a[5]), .B(b[3]), .Z(n47388) );
  AND U47527 ( .A(a[6]), .B(b[3]), .Z(n47349) );
  AND U47528 ( .A(a[7]), .B(b[3]), .Z(n47304) );
  AND U47529 ( .A(a[8]), .B(b[3]), .Z(n47253) );
  AND U47530 ( .A(a[9]), .B(b[3]), .Z(n47197) );
  AND U47531 ( .A(b[3]), .B(a[10]), .Z(n47134) );
  AND U47532 ( .A(b[3]), .B(a[11]), .Z(n47065) );
  AND U47533 ( .A(b[3]), .B(a[12]), .Z(n46990) );
  AND U47534 ( .A(b[3]), .B(a[13]), .Z(n46909) );
  AND U47535 ( .A(b[3]), .B(a[14]), .Z(n46822) );
  AND U47536 ( .A(b[3]), .B(a[15]), .Z(n46729) );
  AND U47537 ( .A(b[3]), .B(a[16]), .Z(n46630) );
  AND U47538 ( .A(b[3]), .B(a[17]), .Z(n46525) );
  AND U47539 ( .A(b[3]), .B(a[18]), .Z(n46414) );
  AND U47540 ( .A(b[3]), .B(a[19]), .Z(n46297) );
  AND U47541 ( .A(b[3]), .B(a[20]), .Z(n46174) );
  AND U47542 ( .A(b[3]), .B(a[21]), .Z(n46045) );
  AND U47543 ( .A(b[3]), .B(a[22]), .Z(n45910) );
  AND U47544 ( .A(b[3]), .B(a[23]), .Z(n45769) );
  AND U47545 ( .A(b[3]), .B(a[24]), .Z(n45622) );
  AND U47546 ( .A(b[3]), .B(a[25]), .Z(n45469) );
  AND U47547 ( .A(b[3]), .B(a[26]), .Z(n45310) );
  AND U47548 ( .A(b[3]), .B(a[27]), .Z(n45145) );
  AND U47549 ( .A(b[3]), .B(a[28]), .Z(n44974) );
  AND U47550 ( .A(b[3]), .B(a[29]), .Z(n44797) );
  AND U47551 ( .A(b[3]), .B(a[30]), .Z(n44614) );
  AND U47552 ( .A(b[3]), .B(a[31]), .Z(n44425) );
  AND U47553 ( .A(b[3]), .B(a[32]), .Z(n44230) );
  AND U47554 ( .A(b[3]), .B(a[33]), .Z(n44029) );
  AND U47555 ( .A(b[3]), .B(a[34]), .Z(n43822) );
  AND U47556 ( .A(b[3]), .B(a[35]), .Z(n43609) );
  AND U47557 ( .A(b[3]), .B(a[36]), .Z(n43390) );
  AND U47558 ( .A(b[3]), .B(a[37]), .Z(n43165) );
  AND U47559 ( .A(b[3]), .B(a[38]), .Z(n42934) );
  AND U47560 ( .A(b[3]), .B(a[39]), .Z(n42697) );
  AND U47561 ( .A(b[3]), .B(a[40]), .Z(n42454) );
  AND U47562 ( .A(b[3]), .B(a[41]), .Z(n42205) );
  AND U47563 ( .A(b[3]), .B(a[42]), .Z(n41950) );
  AND U47564 ( .A(b[3]), .B(a[43]), .Z(n41689) );
  AND U47565 ( .A(b[3]), .B(a[44]), .Z(n41422) );
  AND U47566 ( .A(b[3]), .B(a[45]), .Z(n41149) );
  AND U47567 ( .A(b[3]), .B(a[46]), .Z(n40870) );
  AND U47568 ( .A(b[3]), .B(a[47]), .Z(n40585) );
  AND U47569 ( .A(b[3]), .B(a[48]), .Z(n40294) );
  AND U47570 ( .A(b[3]), .B(a[49]), .Z(n39997) );
  AND U47571 ( .A(b[3]), .B(a[50]), .Z(n39694) );
  AND U47572 ( .A(b[3]), .B(a[51]), .Z(n39385) );
  AND U47573 ( .A(b[3]), .B(a[52]), .Z(n39070) );
  AND U47574 ( .A(b[3]), .B(a[53]), .Z(n38749) );
  AND U47575 ( .A(b[3]), .B(a[54]), .Z(n38422) );
  AND U47576 ( .A(b[3]), .B(a[55]), .Z(n38089) );
  AND U47577 ( .A(b[3]), .B(a[56]), .Z(n37750) );
  AND U47578 ( .A(b[3]), .B(a[57]), .Z(n37405) );
  AND U47579 ( .A(b[3]), .B(a[58]), .Z(n37054) );
  AND U47580 ( .A(b[3]), .B(a[59]), .Z(n36697) );
  AND U47581 ( .A(b[3]), .B(a[60]), .Z(n36334) );
  AND U47582 ( .A(b[3]), .B(a[61]), .Z(n35965) );
  AND U47583 ( .A(b[3]), .B(a[62]), .Z(n35590) );
  AND U47584 ( .A(b[3]), .B(a[63]), .Z(n35209) );
  AND U47585 ( .A(b[3]), .B(a[64]), .Z(n34822) );
  AND U47586 ( .A(b[3]), .B(a[65]), .Z(n34429) );
  AND U47587 ( .A(b[3]), .B(a[66]), .Z(n34030) );
  AND U47588 ( .A(b[3]), .B(a[67]), .Z(n33625) );
  AND U47589 ( .A(b[3]), .B(a[68]), .Z(n33214) );
  AND U47590 ( .A(b[3]), .B(a[69]), .Z(n32797) );
  AND U47591 ( .A(b[3]), .B(a[70]), .Z(n32374) );
  AND U47592 ( .A(b[3]), .B(a[71]), .Z(n31945) );
  AND U47593 ( .A(b[3]), .B(a[72]), .Z(n31510) );
  AND U47594 ( .A(b[3]), .B(a[73]), .Z(n31069) );
  AND U47595 ( .A(b[3]), .B(a[74]), .Z(n30622) );
  AND U47596 ( .A(b[3]), .B(a[75]), .Z(n30169) );
  AND U47597 ( .A(b[3]), .B(a[76]), .Z(n29710) );
  AND U47598 ( .A(b[3]), .B(a[77]), .Z(n29245) );
  AND U47599 ( .A(b[3]), .B(a[78]), .Z(n28774) );
  AND U47600 ( .A(b[3]), .B(a[79]), .Z(n28297) );
  AND U47601 ( .A(b[3]), .B(a[80]), .Z(n27814) );
  AND U47602 ( .A(b[3]), .B(a[81]), .Z(n27325) );
  AND U47603 ( .A(b[3]), .B(a[82]), .Z(n26828) );
  AND U47604 ( .A(b[3]), .B(a[83]), .Z(n26327) );
  AND U47605 ( .A(b[3]), .B(a[84]), .Z(n25819) );
  AND U47606 ( .A(b[3]), .B(a[85]), .Z(n25305) );
  AND U47607 ( .A(b[3]), .B(a[86]), .Z(n24782) );
  AND U47608 ( .A(b[3]), .B(a[87]), .Z(n24257) );
  AND U47609 ( .A(b[3]), .B(a[88]), .Z(n23726) );
  AND U47610 ( .A(b[3]), .B(a[89]), .Z(n23188) );
  AND U47611 ( .A(b[3]), .B(a[90]), .Z(n22644) );
  AND U47612 ( .A(b[3]), .B(a[91]), .Z(n22095) );
  AND U47613 ( .A(b[3]), .B(a[92]), .Z(n21540) );
  AND U47614 ( .A(b[3]), .B(a[93]), .Z(n20978) );
  AND U47615 ( .A(b[3]), .B(a[94]), .Z(n20411) );
  AND U47616 ( .A(b[3]), .B(a[95]), .Z(n19838) );
  AND U47617 ( .A(b[3]), .B(a[96]), .Z(n19259) );
  AND U47618 ( .A(b[3]), .B(a[97]), .Z(n18578) );
  NAND U47619 ( .A(a[100]), .B(b[0]), .Z(n17392) );
  AND U47620 ( .A(b[0]), .B(a[0]), .Z(c[0]) );
endmodule

