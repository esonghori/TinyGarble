
module FA_32 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_64 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_96 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_33 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_992 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_960 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_928 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_896 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_864 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_832 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_800 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_768 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_736 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_704 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_672 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_640 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_608 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_576 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_544 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_512 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_480 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_448 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_416 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_384 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_352 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_320 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_288 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_256 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_224 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_192 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_160 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_128 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_96 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_64 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_32 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_1025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_34 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_1055 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1054 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1053 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1052 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1051 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1050 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1049 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1048 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1047 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1046 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1045 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1044 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1043 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1042 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1041 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1040 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1039 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1038 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1037 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1036 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1035 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1034 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1033 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1032 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1031 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1030 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1029 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1028 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_1027 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_1026 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_1025 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_1057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_35 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1087 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1086 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1085 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1084 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1083 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1082 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1081 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1080 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1079 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1078 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1077 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1076 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1075 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1074 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1073 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1072 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1071 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1070 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1069 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1068 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1067 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1066 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1065 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1064 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1063 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1062 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1061 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1060 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_1059 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_1058 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1057 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_36 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1119 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1118 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1117 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1116 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1115 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1114 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1113 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1112 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1111 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1110 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1109 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1108 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1107 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1106 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1105 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1104 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1103 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1102 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1101 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1100 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1099 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1098 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1097 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1096 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1095 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1094 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1093 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_1092 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_1091 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1090 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1089 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_37 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1151 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1150 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1149 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1148 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1147 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1146 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1145 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1144 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1143 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1142 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1141 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1140 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1139 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1138 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1137 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1136 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1135 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1134 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1133 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1132 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1131 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1130 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1129 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1128 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1127 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1126 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_1125 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_1124 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1123 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1122 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1121 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_38 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1183 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1182 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1181 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1180 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1179 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1178 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1177 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1176 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1175 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1174 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1173 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1172 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1171 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1170 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1169 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1168 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1167 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1166 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1165 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1164 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1163 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1162 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1161 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1160 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1159 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_1158 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_1157 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1156 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1155 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1154 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1153 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_39 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1215 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1214 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1213 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1212 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1211 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1210 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1209 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1208 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1207 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1206 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1205 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1204 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1203 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1202 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1201 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1200 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1199 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1198 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1197 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1196 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1195 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1194 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1193 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1192 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_1191 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_1190 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1189 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1188 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1187 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1186 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1185 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_40 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1247 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1246 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1245 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1244 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1243 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1242 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1241 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1240 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1239 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1238 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1237 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1236 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1235 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1234 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1233 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1232 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1231 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1230 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1229 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1228 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1227 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1226 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1225 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_1224 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_1223 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1222 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1221 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1220 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1219 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1218 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1217 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_41 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1279 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1278 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1277 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1276 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1275 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1274 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1273 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1272 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1271 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1270 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1269 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1268 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1267 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1266 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1265 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1264 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1263 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1262 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1261 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1260 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1259 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1258 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_1257 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_1256 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1255 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1254 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1253 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1252 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1251 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1250 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1249 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_42 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1311 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1310 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1309 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1308 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1307 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1306 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1305 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1304 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1303 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1302 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1301 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1300 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1299 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1298 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1297 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1296 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1295 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1294 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1293 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1292 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1291 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_1290 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_1289 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1288 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1287 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1286 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1285 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1284 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1283 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1282 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1281 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_43 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1343 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1342 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1341 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1340 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1339 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1338 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1337 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1336 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1335 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1334 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1333 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1332 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1331 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1330 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1329 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1328 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1327 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1326 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1325 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1324 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_1323 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_1322 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1321 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1320 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1319 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1318 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1317 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1316 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1315 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1314 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1313 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_44 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1375 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1374 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1373 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1372 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1371 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1370 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1369 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1368 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1367 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1366 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1365 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1364 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1363 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1362 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1361 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1360 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1359 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1358 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1357 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_1356 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_1355 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1354 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1353 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1352 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1351 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1350 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1349 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1348 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1347 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1346 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1345 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_45 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1407 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1406 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1405 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1404 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1403 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1402 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1401 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1400 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1399 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1398 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1397 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1396 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1395 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1394 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1393 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1392 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1391 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1390 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_1389 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_1388 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1387 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1386 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1385 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1384 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1383 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1382 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1381 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1380 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1379 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1378 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1377 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_46 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1439 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1438 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1437 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1436 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1435 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1434 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1433 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1432 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1431 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1430 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1429 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1428 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1427 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1426 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1425 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1424 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1423 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_1422 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_1421 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1420 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1419 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1418 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1417 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1416 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1415 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1414 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1413 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1412 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1411 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1410 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1409 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_47 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1471 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1470 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1469 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1468 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1467 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1466 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1465 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1464 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1463 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1462 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1461 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1460 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1459 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1458 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1457 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1456 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_1455 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_1454 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1453 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1452 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1451 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1450 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1449 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1448 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1447 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1446 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1445 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1444 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1443 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1442 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1441 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_48 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1503 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1502 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1501 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1500 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1499 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1498 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1497 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1496 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1495 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1494 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1493 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1492 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1491 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1490 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1489 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_1488 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_1487 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1486 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1485 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1484 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1483 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1482 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1481 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1480 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1479 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1478 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1477 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1476 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1475 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1474 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1473 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_49 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1535 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1534 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1533 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1532 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1531 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1530 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1529 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1528 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1527 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1526 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1525 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1524 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1523 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1522 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_1521 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_1520 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1519 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1518 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1517 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1516 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1515 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1514 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1513 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1512 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1511 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1510 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1509 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1508 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1507 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1506 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1505 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_50 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1567 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1566 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1565 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1564 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1563 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1562 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1561 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1560 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1559 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1558 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1557 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1556 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1555 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_1554 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_1553 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1552 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1551 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1550 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1549 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1548 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1547 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1546 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1545 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1544 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1543 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1542 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1541 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1540 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1539 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1538 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1537 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_51 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1599 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1598 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1597 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1596 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1595 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1594 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1593 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1592 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1591 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1590 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1589 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1588 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_1587 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_1586 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1585 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1584 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1583 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1582 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1581 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1580 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1579 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1578 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1577 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1576 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1575 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1574 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1573 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1572 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1571 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1570 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1569 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_52 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1631 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1630 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1629 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1628 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1627 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1626 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1625 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1624 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1623 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1622 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1621 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_1620 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_1619 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1618 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1617 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1616 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1615 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1614 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1613 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1612 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1611 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1610 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1609 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1608 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1607 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1606 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1605 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1604 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1603 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1602 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1601 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_53 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1663 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1662 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1661 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1660 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1659 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1658 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1657 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1656 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1655 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1654 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_1653 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_1652 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1651 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1650 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1649 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1648 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1647 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1646 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1645 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1644 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1643 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1642 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1641 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1640 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1639 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1638 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1637 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1636 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1635 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1634 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1633 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_54 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1695 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1694 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1693 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1692 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1691 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1690 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1689 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1688 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1687 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_1686 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_1685 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1684 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1683 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1682 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1681 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1680 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1679 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1678 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1677 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1676 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1675 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1674 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1673 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1672 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1671 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1670 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1669 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1668 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1667 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1666 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1665 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_55 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1727 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1726 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1725 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1724 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1723 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1722 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1721 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1720 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_1719 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_1718 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1717 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1716 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1715 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1714 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1713 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1712 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1711 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1710 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1709 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1708 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1707 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1706 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1705 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1704 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1703 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1702 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1701 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1700 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1699 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1698 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1697 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_56 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1759 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1758 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1757 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1756 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1755 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1754 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1753 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_1752 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_1751 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1750 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1749 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1748 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1747 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1746 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1745 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1744 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1743 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1742 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1741 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1740 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1739 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1738 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1737 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1736 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1735 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1734 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1733 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1732 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1731 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1730 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1729 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_57 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1791 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1790 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1789 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1788 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1787 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1786 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_1785 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_1784 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1783 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1782 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1781 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1780 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1779 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1778 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1777 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1776 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1775 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1774 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1773 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1772 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1771 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1770 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1769 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1768 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1767 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1766 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1765 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1764 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1763 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1762 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1761 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_58 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1823 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1822 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1821 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1820 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1819 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_1818 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_1817 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1816 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1815 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1814 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1813 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1812 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1811 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1810 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1809 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1808 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1807 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1806 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1805 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1804 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1803 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1802 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1801 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1800 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1799 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1798 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1797 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1796 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1795 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1794 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1793 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_59 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1855 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1854 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1853 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1852 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_1851 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_1850 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1849 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1848 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1847 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1846 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1845 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1844 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1843 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1842 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1841 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1840 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1839 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1838 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1837 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1836 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1835 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1834 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1833 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1832 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1831 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1830 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1829 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1828 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1827 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1826 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1825 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_60 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1887 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1886 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1885 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_1884 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_1883 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1882 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1881 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1880 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1879 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1878 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1877 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1876 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1875 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1874 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1873 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1872 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1871 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1870 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1869 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1868 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1867 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1866 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1865 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1864 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1863 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1862 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1861 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1860 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1859 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1858 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1857 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_61 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1919 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1918 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_1917 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_1916 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_1915 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1914 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1913 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1912 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1911 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1910 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1909 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1908 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1907 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1906 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1905 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1904 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1903 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1902 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1901 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1900 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1899 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1898 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1897 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1896 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1895 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1894 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1893 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1892 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1891 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1890 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1889 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_1951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_62 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_1951 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_1950 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_1949 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_1948 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_1947 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1946 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1945 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1944 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1943 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1942 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1941 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1940 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1939 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1938 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1937 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1936 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1935 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1934 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1933 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1932 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1931 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1930 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1929 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1928 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1927 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1926 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1925 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1924 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1923 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1922 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1921 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_1953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_1983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_63 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_1983 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_1982 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_1981 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_1980 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_1979 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_1978 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_1977 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_1976 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_1975 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_1974 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_1973 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_1972 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_1971 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_1970 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_1969 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_1968 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_1967 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_1966 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_1965 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_1964 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_1963 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_1962 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_1961 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_1960 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_1959 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_1958 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_1957 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_1956 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_1955 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_1954 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_1953 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_1 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_63 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_62 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_61 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_60 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_59 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_58 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_57 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_56 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_55 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_54 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_53 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_52 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_51 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_50 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_49 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_48 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_47 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_46 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_45 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_44 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_43 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_42 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_41 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_40 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_39 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_38 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_37 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_36 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_35 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_34 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_33 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_1985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_1986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_32 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_2015 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_2014 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_2013 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_2012 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_2011 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2010 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2009 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2008 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2007 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2006 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2005 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2004 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2003 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2002 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2001 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2000 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1999 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1998 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1997 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1996 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1995 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1994 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1993 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1992 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1991 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1990 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1989 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1988 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1987 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1986 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1985 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module matrixMult_N_M_3_N5_M32 ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;

  wire   [31:0] xy;
  wire   [31:0] oi;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign o[0] = 1'b0;

  MULT_N32_1 MULT_ ( .A({x[31:1], 1'b0}), .B({1'b0, y[30:0]}), .O({xy[31:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_32 ADD_ ( .A({xy[31:1], 1'b0}), .B({o[31:1], 1'b0}), .CI(1'b0), .S({
        oi[31:1], SYNOPSYS_UNCONNECTED__1}) );
  DFF \o_reg[1]  ( .D(oi[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[1]) );
  DFF \o_reg[2]  ( .D(oi[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[2]) );
  DFF \o_reg[3]  ( .D(oi[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[3]) );
  DFF \o_reg[4]  ( .D(oi[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[4]) );
  DFF \o_reg[5]  ( .D(oi[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[5]) );
  DFF \o_reg[6]  ( .D(oi[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[6]) );
  DFF \o_reg[7]  ( .D(oi[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[7]) );
  DFF \o_reg[8]  ( .D(oi[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[8]) );
  DFF \o_reg[9]  ( .D(oi[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[9]) );
  DFF \o_reg[10]  ( .D(oi[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[10]) );
  DFF \o_reg[11]  ( .D(oi[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[11]) );
  DFF \o_reg[12]  ( .D(oi[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[12]) );
  DFF \o_reg[13]  ( .D(oi[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[13]) );
  DFF \o_reg[14]  ( .D(oi[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[14]) );
  DFF \o_reg[15]  ( .D(oi[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[15]) );
  DFF \o_reg[16]  ( .D(oi[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[16]) );
  DFF \o_reg[17]  ( .D(oi[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[17]) );
  DFF \o_reg[18]  ( .D(oi[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[18]) );
  DFF \o_reg[19]  ( .D(oi[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[19]) );
  DFF \o_reg[20]  ( .D(oi[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[20]) );
  DFF \o_reg[21]  ( .D(oi[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[21]) );
  DFF \o_reg[22]  ( .D(oi[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[22]) );
  DFF \o_reg[23]  ( .D(oi[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[23]) );
  DFF \o_reg[24]  ( .D(oi[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[24]) );
  DFF \o_reg[25]  ( .D(oi[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[25]) );
  DFF \o_reg[26]  ( .D(oi[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[26]) );
  DFF \o_reg[27]  ( .D(oi[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[27]) );
  DFF \o_reg[28]  ( .D(oi[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[28]) );
  DFF \o_reg[29]  ( .D(oi[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[29]) );
  DFF \o_reg[30]  ( .D(oi[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[30]) );
  DFF \o_reg[31]  ( .D(oi[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[31]) );
endmodule

