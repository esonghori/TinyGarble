
module sum_N1024_CC8 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n5) );
  NAND U6 ( .A(a[0]), .B(b[0]), .Z(n3) );
  NAND U7 ( .A(n1), .B(carry_on), .Z(n2) );
  NAND U8 ( .A(n3), .B(n2), .Z(n4) );
  XOR U9 ( .A(n5), .B(n4), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n9) );
  NAND U11 ( .A(a[1]), .B(b[1]), .Z(n7) );
  NAND U12 ( .A(n5), .B(n4), .Z(n6) );
  NAND U13 ( .A(n7), .B(n6), .Z(n8) );
  XOR U14 ( .A(n9), .B(n8), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n13) );
  NAND U16 ( .A(a[2]), .B(b[2]), .Z(n11) );
  NAND U17 ( .A(n9), .B(n8), .Z(n10) );
  NAND U18 ( .A(n11), .B(n10), .Z(n12) );
  XOR U19 ( .A(n13), .B(n12), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n17) );
  NAND U21 ( .A(a[3]), .B(b[3]), .Z(n15) );
  NAND U22 ( .A(n13), .B(n12), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n16) );
  XOR U24 ( .A(n17), .B(n16), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n21) );
  NAND U26 ( .A(a[4]), .B(b[4]), .Z(n19) );
  NAND U27 ( .A(n17), .B(n16), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n20) );
  XOR U29 ( .A(n21), .B(n20), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n25) );
  NAND U31 ( .A(a[5]), .B(b[5]), .Z(n23) );
  NAND U32 ( .A(n21), .B(n20), .Z(n22) );
  NAND U33 ( .A(n23), .B(n22), .Z(n24) );
  XOR U34 ( .A(n25), .B(n24), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n29) );
  NAND U36 ( .A(a[6]), .B(b[6]), .Z(n27) );
  NAND U37 ( .A(n25), .B(n24), .Z(n26) );
  NAND U38 ( .A(n27), .B(n26), .Z(n28) );
  XOR U39 ( .A(n29), .B(n28), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n33) );
  NAND U41 ( .A(a[7]), .B(b[7]), .Z(n31) );
  NAND U42 ( .A(n29), .B(n28), .Z(n30) );
  NAND U43 ( .A(n31), .B(n30), .Z(n32) );
  XOR U44 ( .A(n33), .B(n32), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n37) );
  NAND U46 ( .A(a[8]), .B(b[8]), .Z(n35) );
  NAND U47 ( .A(n33), .B(n32), .Z(n34) );
  NAND U48 ( .A(n35), .B(n34), .Z(n36) );
  XOR U49 ( .A(n37), .B(n36), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n41) );
  NAND U51 ( .A(a[9]), .B(b[9]), .Z(n39) );
  NAND U52 ( .A(n37), .B(n36), .Z(n38) );
  NAND U53 ( .A(n39), .B(n38), .Z(n40) );
  XOR U54 ( .A(n41), .B(n40), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n45) );
  NAND U56 ( .A(a[10]), .B(b[10]), .Z(n43) );
  NAND U57 ( .A(n41), .B(n40), .Z(n42) );
  NAND U58 ( .A(n43), .B(n42), .Z(n44) );
  XOR U59 ( .A(n45), .B(n44), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n49) );
  NAND U61 ( .A(a[11]), .B(b[11]), .Z(n47) );
  NAND U62 ( .A(n45), .B(n44), .Z(n46) );
  NAND U63 ( .A(n47), .B(n46), .Z(n48) );
  XOR U64 ( .A(n49), .B(n48), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n53) );
  NAND U66 ( .A(a[12]), .B(b[12]), .Z(n51) );
  NAND U67 ( .A(n49), .B(n48), .Z(n50) );
  NAND U68 ( .A(n51), .B(n50), .Z(n52) );
  XOR U69 ( .A(n53), .B(n52), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n57) );
  NAND U71 ( .A(a[13]), .B(b[13]), .Z(n55) );
  NAND U72 ( .A(n53), .B(n52), .Z(n54) );
  NAND U73 ( .A(n55), .B(n54), .Z(n56) );
  XOR U74 ( .A(n57), .B(n56), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n61) );
  NAND U76 ( .A(a[14]), .B(b[14]), .Z(n59) );
  NAND U77 ( .A(n57), .B(n56), .Z(n58) );
  NAND U78 ( .A(n59), .B(n58), .Z(n60) );
  XOR U79 ( .A(n61), .B(n60), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n65) );
  NAND U81 ( .A(a[15]), .B(b[15]), .Z(n63) );
  NAND U82 ( .A(n61), .B(n60), .Z(n62) );
  NAND U83 ( .A(n63), .B(n62), .Z(n64) );
  XOR U84 ( .A(n65), .B(n64), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n69) );
  NAND U86 ( .A(a[16]), .B(b[16]), .Z(n67) );
  NAND U87 ( .A(n65), .B(n64), .Z(n66) );
  NAND U88 ( .A(n67), .B(n66), .Z(n68) );
  XOR U89 ( .A(n69), .B(n68), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n73) );
  NAND U91 ( .A(a[17]), .B(b[17]), .Z(n71) );
  NAND U92 ( .A(n69), .B(n68), .Z(n70) );
  NAND U93 ( .A(n71), .B(n70), .Z(n72) );
  XOR U94 ( .A(n73), .B(n72), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n77) );
  NAND U96 ( .A(a[18]), .B(b[18]), .Z(n75) );
  NAND U97 ( .A(n73), .B(n72), .Z(n74) );
  NAND U98 ( .A(n75), .B(n74), .Z(n76) );
  XOR U99 ( .A(n77), .B(n76), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n81) );
  NAND U101 ( .A(a[19]), .B(b[19]), .Z(n79) );
  NAND U102 ( .A(n77), .B(n76), .Z(n78) );
  NAND U103 ( .A(n79), .B(n78), .Z(n80) );
  XOR U104 ( .A(n81), .B(n80), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n85) );
  NAND U106 ( .A(a[20]), .B(b[20]), .Z(n83) );
  NAND U107 ( .A(n81), .B(n80), .Z(n82) );
  NAND U108 ( .A(n83), .B(n82), .Z(n84) );
  XOR U109 ( .A(n85), .B(n84), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n89) );
  NAND U111 ( .A(a[21]), .B(b[21]), .Z(n87) );
  NAND U112 ( .A(n85), .B(n84), .Z(n86) );
  NAND U113 ( .A(n87), .B(n86), .Z(n88) );
  XOR U114 ( .A(n89), .B(n88), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n93) );
  NAND U116 ( .A(a[22]), .B(b[22]), .Z(n91) );
  NAND U117 ( .A(n89), .B(n88), .Z(n90) );
  NAND U118 ( .A(n91), .B(n90), .Z(n92) );
  XOR U119 ( .A(n93), .B(n92), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n97) );
  NAND U121 ( .A(a[23]), .B(b[23]), .Z(n95) );
  NAND U122 ( .A(n93), .B(n92), .Z(n94) );
  NAND U123 ( .A(n95), .B(n94), .Z(n96) );
  XOR U124 ( .A(n97), .B(n96), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n101) );
  NAND U126 ( .A(a[24]), .B(b[24]), .Z(n99) );
  NAND U127 ( .A(n97), .B(n96), .Z(n98) );
  NAND U128 ( .A(n99), .B(n98), .Z(n100) );
  XOR U129 ( .A(n101), .B(n100), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n105) );
  NAND U131 ( .A(a[25]), .B(b[25]), .Z(n103) );
  NAND U132 ( .A(n101), .B(n100), .Z(n102) );
  NAND U133 ( .A(n103), .B(n102), .Z(n104) );
  XOR U134 ( .A(n105), .B(n104), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n109) );
  NAND U136 ( .A(a[26]), .B(b[26]), .Z(n107) );
  NAND U137 ( .A(n105), .B(n104), .Z(n106) );
  NAND U138 ( .A(n107), .B(n106), .Z(n108) );
  XOR U139 ( .A(n109), .B(n108), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n113) );
  NAND U141 ( .A(a[27]), .B(b[27]), .Z(n111) );
  NAND U142 ( .A(n109), .B(n108), .Z(n110) );
  NAND U143 ( .A(n111), .B(n110), .Z(n112) );
  XOR U144 ( .A(n113), .B(n112), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n117) );
  NAND U146 ( .A(a[28]), .B(b[28]), .Z(n115) );
  NAND U147 ( .A(n113), .B(n112), .Z(n114) );
  NAND U148 ( .A(n115), .B(n114), .Z(n116) );
  XOR U149 ( .A(n117), .B(n116), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n121) );
  NAND U151 ( .A(a[29]), .B(b[29]), .Z(n119) );
  NAND U152 ( .A(n117), .B(n116), .Z(n118) );
  NAND U153 ( .A(n119), .B(n118), .Z(n120) );
  XOR U154 ( .A(n121), .B(n120), .Z(c[30]) );
  XOR U155 ( .A(a[31]), .B(b[31]), .Z(n125) );
  NAND U156 ( .A(a[30]), .B(b[30]), .Z(n123) );
  NAND U157 ( .A(n121), .B(n120), .Z(n122) );
  NAND U158 ( .A(n123), .B(n122), .Z(n124) );
  XOR U159 ( .A(n125), .B(n124), .Z(c[31]) );
  XOR U160 ( .A(a[32]), .B(b[32]), .Z(n129) );
  NAND U161 ( .A(a[31]), .B(b[31]), .Z(n127) );
  NAND U162 ( .A(n125), .B(n124), .Z(n126) );
  NAND U163 ( .A(n127), .B(n126), .Z(n128) );
  XOR U164 ( .A(n129), .B(n128), .Z(c[32]) );
  XOR U165 ( .A(a[33]), .B(b[33]), .Z(n133) );
  NAND U166 ( .A(a[32]), .B(b[32]), .Z(n131) );
  NAND U167 ( .A(n129), .B(n128), .Z(n130) );
  NAND U168 ( .A(n131), .B(n130), .Z(n132) );
  XOR U169 ( .A(n133), .B(n132), .Z(c[33]) );
  XOR U170 ( .A(a[34]), .B(b[34]), .Z(n137) );
  NAND U171 ( .A(a[33]), .B(b[33]), .Z(n135) );
  NAND U172 ( .A(n133), .B(n132), .Z(n134) );
  NAND U173 ( .A(n135), .B(n134), .Z(n136) );
  XOR U174 ( .A(n137), .B(n136), .Z(c[34]) );
  XOR U175 ( .A(a[35]), .B(b[35]), .Z(n141) );
  NAND U176 ( .A(a[34]), .B(b[34]), .Z(n139) );
  NAND U177 ( .A(n137), .B(n136), .Z(n138) );
  NAND U178 ( .A(n139), .B(n138), .Z(n140) );
  XOR U179 ( .A(n141), .B(n140), .Z(c[35]) );
  XOR U180 ( .A(a[36]), .B(b[36]), .Z(n145) );
  NAND U181 ( .A(a[35]), .B(b[35]), .Z(n143) );
  NAND U182 ( .A(n141), .B(n140), .Z(n142) );
  NAND U183 ( .A(n143), .B(n142), .Z(n144) );
  XOR U184 ( .A(n145), .B(n144), .Z(c[36]) );
  XOR U185 ( .A(a[37]), .B(b[37]), .Z(n149) );
  NAND U186 ( .A(a[36]), .B(b[36]), .Z(n147) );
  NAND U187 ( .A(n145), .B(n144), .Z(n146) );
  NAND U188 ( .A(n147), .B(n146), .Z(n148) );
  XOR U189 ( .A(n149), .B(n148), .Z(c[37]) );
  XOR U190 ( .A(a[38]), .B(b[38]), .Z(n153) );
  NAND U191 ( .A(a[37]), .B(b[37]), .Z(n151) );
  NAND U192 ( .A(n149), .B(n148), .Z(n150) );
  NAND U193 ( .A(n151), .B(n150), .Z(n152) );
  XOR U194 ( .A(n153), .B(n152), .Z(c[38]) );
  XOR U195 ( .A(a[39]), .B(b[39]), .Z(n157) );
  NAND U196 ( .A(a[38]), .B(b[38]), .Z(n155) );
  NAND U197 ( .A(n153), .B(n152), .Z(n154) );
  NAND U198 ( .A(n155), .B(n154), .Z(n156) );
  XOR U199 ( .A(n157), .B(n156), .Z(c[39]) );
  XOR U200 ( .A(a[40]), .B(b[40]), .Z(n161) );
  NAND U201 ( .A(a[39]), .B(b[39]), .Z(n159) );
  NAND U202 ( .A(n157), .B(n156), .Z(n158) );
  NAND U203 ( .A(n159), .B(n158), .Z(n160) );
  XOR U204 ( .A(n161), .B(n160), .Z(c[40]) );
  XOR U205 ( .A(a[41]), .B(b[41]), .Z(n165) );
  NAND U206 ( .A(a[40]), .B(b[40]), .Z(n163) );
  NAND U207 ( .A(n161), .B(n160), .Z(n162) );
  NAND U208 ( .A(n163), .B(n162), .Z(n164) );
  XOR U209 ( .A(n165), .B(n164), .Z(c[41]) );
  XOR U210 ( .A(a[42]), .B(b[42]), .Z(n169) );
  NAND U211 ( .A(a[41]), .B(b[41]), .Z(n167) );
  NAND U212 ( .A(n165), .B(n164), .Z(n166) );
  NAND U213 ( .A(n167), .B(n166), .Z(n168) );
  XOR U214 ( .A(n169), .B(n168), .Z(c[42]) );
  XOR U215 ( .A(a[43]), .B(b[43]), .Z(n173) );
  NAND U216 ( .A(a[42]), .B(b[42]), .Z(n171) );
  NAND U217 ( .A(n169), .B(n168), .Z(n170) );
  NAND U218 ( .A(n171), .B(n170), .Z(n172) );
  XOR U219 ( .A(n173), .B(n172), .Z(c[43]) );
  XOR U220 ( .A(a[44]), .B(b[44]), .Z(n177) );
  NAND U221 ( .A(a[43]), .B(b[43]), .Z(n175) );
  NAND U222 ( .A(n173), .B(n172), .Z(n174) );
  NAND U223 ( .A(n175), .B(n174), .Z(n176) );
  XOR U224 ( .A(n177), .B(n176), .Z(c[44]) );
  XOR U225 ( .A(a[45]), .B(b[45]), .Z(n181) );
  NAND U226 ( .A(a[44]), .B(b[44]), .Z(n179) );
  NAND U227 ( .A(n177), .B(n176), .Z(n178) );
  NAND U228 ( .A(n179), .B(n178), .Z(n180) );
  XOR U229 ( .A(n181), .B(n180), .Z(c[45]) );
  XOR U230 ( .A(a[46]), .B(b[46]), .Z(n185) );
  NAND U231 ( .A(a[45]), .B(b[45]), .Z(n183) );
  NAND U232 ( .A(n181), .B(n180), .Z(n182) );
  NAND U233 ( .A(n183), .B(n182), .Z(n184) );
  XOR U234 ( .A(n185), .B(n184), .Z(c[46]) );
  XOR U235 ( .A(a[47]), .B(b[47]), .Z(n189) );
  NAND U236 ( .A(a[46]), .B(b[46]), .Z(n187) );
  NAND U237 ( .A(n185), .B(n184), .Z(n186) );
  NAND U238 ( .A(n187), .B(n186), .Z(n188) );
  XOR U239 ( .A(n189), .B(n188), .Z(c[47]) );
  XOR U240 ( .A(a[48]), .B(b[48]), .Z(n193) );
  NAND U241 ( .A(a[47]), .B(b[47]), .Z(n191) );
  NAND U242 ( .A(n189), .B(n188), .Z(n190) );
  NAND U243 ( .A(n191), .B(n190), .Z(n192) );
  XOR U244 ( .A(n193), .B(n192), .Z(c[48]) );
  XOR U245 ( .A(a[49]), .B(b[49]), .Z(n197) );
  NAND U246 ( .A(a[48]), .B(b[48]), .Z(n195) );
  NAND U247 ( .A(n193), .B(n192), .Z(n194) );
  NAND U248 ( .A(n195), .B(n194), .Z(n196) );
  XOR U249 ( .A(n197), .B(n196), .Z(c[49]) );
  XOR U250 ( .A(a[50]), .B(b[50]), .Z(n201) );
  NAND U251 ( .A(a[49]), .B(b[49]), .Z(n199) );
  NAND U252 ( .A(n197), .B(n196), .Z(n198) );
  NAND U253 ( .A(n199), .B(n198), .Z(n200) );
  XOR U254 ( .A(n201), .B(n200), .Z(c[50]) );
  XOR U255 ( .A(a[51]), .B(b[51]), .Z(n205) );
  NAND U256 ( .A(a[50]), .B(b[50]), .Z(n203) );
  NAND U257 ( .A(n201), .B(n200), .Z(n202) );
  NAND U258 ( .A(n203), .B(n202), .Z(n204) );
  XOR U259 ( .A(n205), .B(n204), .Z(c[51]) );
  XOR U260 ( .A(a[52]), .B(b[52]), .Z(n209) );
  NAND U261 ( .A(a[51]), .B(b[51]), .Z(n207) );
  NAND U262 ( .A(n205), .B(n204), .Z(n206) );
  NAND U263 ( .A(n207), .B(n206), .Z(n208) );
  XOR U264 ( .A(n209), .B(n208), .Z(c[52]) );
  XOR U265 ( .A(a[53]), .B(b[53]), .Z(n213) );
  NAND U266 ( .A(a[52]), .B(b[52]), .Z(n211) );
  NAND U267 ( .A(n209), .B(n208), .Z(n210) );
  NAND U268 ( .A(n211), .B(n210), .Z(n212) );
  XOR U269 ( .A(n213), .B(n212), .Z(c[53]) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n217) );
  NAND U271 ( .A(a[53]), .B(b[53]), .Z(n215) );
  NAND U272 ( .A(n213), .B(n212), .Z(n214) );
  NAND U273 ( .A(n215), .B(n214), .Z(n216) );
  XOR U274 ( .A(n217), .B(n216), .Z(c[54]) );
  XOR U275 ( .A(a[55]), .B(b[55]), .Z(n221) );
  NAND U276 ( .A(a[54]), .B(b[54]), .Z(n219) );
  NAND U277 ( .A(n217), .B(n216), .Z(n218) );
  NAND U278 ( .A(n219), .B(n218), .Z(n220) );
  XOR U279 ( .A(n221), .B(n220), .Z(c[55]) );
  XOR U280 ( .A(a[56]), .B(b[56]), .Z(n225) );
  NAND U281 ( .A(a[55]), .B(b[55]), .Z(n223) );
  NAND U282 ( .A(n221), .B(n220), .Z(n222) );
  NAND U283 ( .A(n223), .B(n222), .Z(n224) );
  XOR U284 ( .A(n225), .B(n224), .Z(c[56]) );
  XOR U285 ( .A(a[57]), .B(b[57]), .Z(n229) );
  NAND U286 ( .A(a[56]), .B(b[56]), .Z(n227) );
  NAND U287 ( .A(n225), .B(n224), .Z(n226) );
  NAND U288 ( .A(n227), .B(n226), .Z(n228) );
  XOR U289 ( .A(n229), .B(n228), .Z(c[57]) );
  XOR U290 ( .A(a[58]), .B(b[58]), .Z(n233) );
  NAND U291 ( .A(a[57]), .B(b[57]), .Z(n231) );
  NAND U292 ( .A(n229), .B(n228), .Z(n230) );
  NAND U293 ( .A(n231), .B(n230), .Z(n232) );
  XOR U294 ( .A(n233), .B(n232), .Z(c[58]) );
  XOR U295 ( .A(a[59]), .B(b[59]), .Z(n237) );
  NAND U296 ( .A(a[58]), .B(b[58]), .Z(n235) );
  NAND U297 ( .A(n233), .B(n232), .Z(n234) );
  NAND U298 ( .A(n235), .B(n234), .Z(n236) );
  XOR U299 ( .A(n237), .B(n236), .Z(c[59]) );
  XOR U300 ( .A(a[60]), .B(b[60]), .Z(n241) );
  NAND U301 ( .A(a[59]), .B(b[59]), .Z(n239) );
  NAND U302 ( .A(n237), .B(n236), .Z(n238) );
  NAND U303 ( .A(n239), .B(n238), .Z(n240) );
  XOR U304 ( .A(n241), .B(n240), .Z(c[60]) );
  XOR U305 ( .A(a[61]), .B(b[61]), .Z(n245) );
  NAND U306 ( .A(a[60]), .B(b[60]), .Z(n243) );
  NAND U307 ( .A(n241), .B(n240), .Z(n242) );
  NAND U308 ( .A(n243), .B(n242), .Z(n244) );
  XOR U309 ( .A(n245), .B(n244), .Z(c[61]) );
  XOR U310 ( .A(a[62]), .B(b[62]), .Z(n249) );
  NAND U311 ( .A(a[61]), .B(b[61]), .Z(n247) );
  NAND U312 ( .A(n245), .B(n244), .Z(n246) );
  NAND U313 ( .A(n247), .B(n246), .Z(n248) );
  XOR U314 ( .A(n249), .B(n248), .Z(c[62]) );
  XOR U315 ( .A(a[63]), .B(b[63]), .Z(n253) );
  NAND U316 ( .A(a[62]), .B(b[62]), .Z(n251) );
  NAND U317 ( .A(n249), .B(n248), .Z(n250) );
  NAND U318 ( .A(n251), .B(n250), .Z(n252) );
  XOR U319 ( .A(n253), .B(n252), .Z(c[63]) );
  XOR U320 ( .A(a[64]), .B(b[64]), .Z(n257) );
  NAND U321 ( .A(a[63]), .B(b[63]), .Z(n255) );
  NAND U322 ( .A(n253), .B(n252), .Z(n254) );
  NAND U323 ( .A(n255), .B(n254), .Z(n256) );
  XOR U324 ( .A(n257), .B(n256), .Z(c[64]) );
  XOR U325 ( .A(a[65]), .B(b[65]), .Z(n261) );
  NAND U326 ( .A(a[64]), .B(b[64]), .Z(n259) );
  NAND U327 ( .A(n257), .B(n256), .Z(n258) );
  NAND U328 ( .A(n259), .B(n258), .Z(n260) );
  XOR U329 ( .A(n261), .B(n260), .Z(c[65]) );
  XOR U330 ( .A(a[66]), .B(b[66]), .Z(n265) );
  NAND U331 ( .A(a[65]), .B(b[65]), .Z(n263) );
  NAND U332 ( .A(n261), .B(n260), .Z(n262) );
  NAND U333 ( .A(n263), .B(n262), .Z(n264) );
  XOR U334 ( .A(n265), .B(n264), .Z(c[66]) );
  XOR U335 ( .A(a[67]), .B(b[67]), .Z(n269) );
  NAND U336 ( .A(a[66]), .B(b[66]), .Z(n267) );
  NAND U337 ( .A(n265), .B(n264), .Z(n266) );
  NAND U338 ( .A(n267), .B(n266), .Z(n268) );
  XOR U339 ( .A(n269), .B(n268), .Z(c[67]) );
  XOR U340 ( .A(a[68]), .B(b[68]), .Z(n273) );
  NAND U341 ( .A(a[67]), .B(b[67]), .Z(n271) );
  NAND U342 ( .A(n269), .B(n268), .Z(n270) );
  NAND U343 ( .A(n271), .B(n270), .Z(n272) );
  XOR U344 ( .A(n273), .B(n272), .Z(c[68]) );
  XOR U345 ( .A(a[69]), .B(b[69]), .Z(n277) );
  NAND U346 ( .A(a[68]), .B(b[68]), .Z(n275) );
  NAND U347 ( .A(n273), .B(n272), .Z(n274) );
  NAND U348 ( .A(n275), .B(n274), .Z(n276) );
  XOR U349 ( .A(n277), .B(n276), .Z(c[69]) );
  XOR U350 ( .A(a[70]), .B(b[70]), .Z(n281) );
  NAND U351 ( .A(a[69]), .B(b[69]), .Z(n279) );
  NAND U352 ( .A(n277), .B(n276), .Z(n278) );
  NAND U353 ( .A(n279), .B(n278), .Z(n280) );
  XOR U354 ( .A(n281), .B(n280), .Z(c[70]) );
  XOR U355 ( .A(a[71]), .B(b[71]), .Z(n285) );
  NAND U356 ( .A(a[70]), .B(b[70]), .Z(n283) );
  NAND U357 ( .A(n281), .B(n280), .Z(n282) );
  NAND U358 ( .A(n283), .B(n282), .Z(n284) );
  XOR U359 ( .A(n285), .B(n284), .Z(c[71]) );
  XOR U360 ( .A(a[72]), .B(b[72]), .Z(n289) );
  NAND U361 ( .A(a[71]), .B(b[71]), .Z(n287) );
  NAND U362 ( .A(n285), .B(n284), .Z(n286) );
  NAND U363 ( .A(n287), .B(n286), .Z(n288) );
  XOR U364 ( .A(n289), .B(n288), .Z(c[72]) );
  XOR U365 ( .A(a[73]), .B(b[73]), .Z(n293) );
  NAND U366 ( .A(a[72]), .B(b[72]), .Z(n291) );
  NAND U367 ( .A(n289), .B(n288), .Z(n290) );
  NAND U368 ( .A(n291), .B(n290), .Z(n292) );
  XOR U369 ( .A(n293), .B(n292), .Z(c[73]) );
  XOR U370 ( .A(a[74]), .B(b[74]), .Z(n297) );
  NAND U371 ( .A(a[73]), .B(b[73]), .Z(n295) );
  NAND U372 ( .A(n293), .B(n292), .Z(n294) );
  NAND U373 ( .A(n295), .B(n294), .Z(n296) );
  XOR U374 ( .A(n297), .B(n296), .Z(c[74]) );
  XOR U375 ( .A(a[75]), .B(b[75]), .Z(n301) );
  NAND U376 ( .A(a[74]), .B(b[74]), .Z(n299) );
  NAND U377 ( .A(n297), .B(n296), .Z(n298) );
  NAND U378 ( .A(n299), .B(n298), .Z(n300) );
  XOR U379 ( .A(n301), .B(n300), .Z(c[75]) );
  XOR U380 ( .A(a[76]), .B(b[76]), .Z(n305) );
  NAND U381 ( .A(a[75]), .B(b[75]), .Z(n303) );
  NAND U382 ( .A(n301), .B(n300), .Z(n302) );
  NAND U383 ( .A(n303), .B(n302), .Z(n304) );
  XOR U384 ( .A(n305), .B(n304), .Z(c[76]) );
  XOR U385 ( .A(a[77]), .B(b[77]), .Z(n309) );
  NAND U386 ( .A(a[76]), .B(b[76]), .Z(n307) );
  NAND U387 ( .A(n305), .B(n304), .Z(n306) );
  NAND U388 ( .A(n307), .B(n306), .Z(n308) );
  XOR U389 ( .A(n309), .B(n308), .Z(c[77]) );
  XOR U390 ( .A(a[78]), .B(b[78]), .Z(n313) );
  NAND U391 ( .A(a[77]), .B(b[77]), .Z(n311) );
  NAND U392 ( .A(n309), .B(n308), .Z(n310) );
  NAND U393 ( .A(n311), .B(n310), .Z(n312) );
  XOR U394 ( .A(n313), .B(n312), .Z(c[78]) );
  XOR U395 ( .A(a[79]), .B(b[79]), .Z(n317) );
  NAND U396 ( .A(a[78]), .B(b[78]), .Z(n315) );
  NAND U397 ( .A(n313), .B(n312), .Z(n314) );
  NAND U398 ( .A(n315), .B(n314), .Z(n316) );
  XOR U399 ( .A(n317), .B(n316), .Z(c[79]) );
  XOR U400 ( .A(a[80]), .B(b[80]), .Z(n321) );
  NAND U401 ( .A(a[79]), .B(b[79]), .Z(n319) );
  NAND U402 ( .A(n317), .B(n316), .Z(n318) );
  NAND U403 ( .A(n319), .B(n318), .Z(n320) );
  XOR U404 ( .A(n321), .B(n320), .Z(c[80]) );
  XOR U405 ( .A(a[81]), .B(b[81]), .Z(n325) );
  NAND U406 ( .A(a[80]), .B(b[80]), .Z(n323) );
  NAND U407 ( .A(n321), .B(n320), .Z(n322) );
  NAND U408 ( .A(n323), .B(n322), .Z(n324) );
  XOR U409 ( .A(n325), .B(n324), .Z(c[81]) );
  XOR U410 ( .A(a[82]), .B(b[82]), .Z(n329) );
  NAND U411 ( .A(a[81]), .B(b[81]), .Z(n327) );
  NAND U412 ( .A(n325), .B(n324), .Z(n326) );
  NAND U413 ( .A(n327), .B(n326), .Z(n328) );
  XOR U414 ( .A(n329), .B(n328), .Z(c[82]) );
  XOR U415 ( .A(a[83]), .B(b[83]), .Z(n333) );
  NAND U416 ( .A(a[82]), .B(b[82]), .Z(n331) );
  NAND U417 ( .A(n329), .B(n328), .Z(n330) );
  NAND U418 ( .A(n331), .B(n330), .Z(n332) );
  XOR U419 ( .A(n333), .B(n332), .Z(c[83]) );
  XOR U420 ( .A(a[84]), .B(b[84]), .Z(n337) );
  NAND U421 ( .A(a[83]), .B(b[83]), .Z(n335) );
  NAND U422 ( .A(n333), .B(n332), .Z(n334) );
  NAND U423 ( .A(n335), .B(n334), .Z(n336) );
  XOR U424 ( .A(n337), .B(n336), .Z(c[84]) );
  XOR U425 ( .A(a[85]), .B(b[85]), .Z(n341) );
  NAND U426 ( .A(a[84]), .B(b[84]), .Z(n339) );
  NAND U427 ( .A(n337), .B(n336), .Z(n338) );
  NAND U428 ( .A(n339), .B(n338), .Z(n340) );
  XOR U429 ( .A(n341), .B(n340), .Z(c[85]) );
  XOR U430 ( .A(a[86]), .B(b[86]), .Z(n345) );
  NAND U431 ( .A(a[85]), .B(b[85]), .Z(n343) );
  NAND U432 ( .A(n341), .B(n340), .Z(n342) );
  NAND U433 ( .A(n343), .B(n342), .Z(n344) );
  XOR U434 ( .A(n345), .B(n344), .Z(c[86]) );
  XOR U435 ( .A(a[87]), .B(b[87]), .Z(n349) );
  NAND U436 ( .A(a[86]), .B(b[86]), .Z(n347) );
  NAND U437 ( .A(n345), .B(n344), .Z(n346) );
  NAND U438 ( .A(n347), .B(n346), .Z(n348) );
  XOR U439 ( .A(n349), .B(n348), .Z(c[87]) );
  XOR U440 ( .A(a[88]), .B(b[88]), .Z(n353) );
  NAND U441 ( .A(a[87]), .B(b[87]), .Z(n351) );
  NAND U442 ( .A(n349), .B(n348), .Z(n350) );
  NAND U443 ( .A(n351), .B(n350), .Z(n352) );
  XOR U444 ( .A(n353), .B(n352), .Z(c[88]) );
  XOR U445 ( .A(a[89]), .B(b[89]), .Z(n357) );
  NAND U446 ( .A(a[88]), .B(b[88]), .Z(n355) );
  NAND U447 ( .A(n353), .B(n352), .Z(n354) );
  NAND U448 ( .A(n355), .B(n354), .Z(n356) );
  XOR U449 ( .A(n357), .B(n356), .Z(c[89]) );
  XOR U450 ( .A(a[90]), .B(b[90]), .Z(n361) );
  NAND U451 ( .A(a[89]), .B(b[89]), .Z(n359) );
  NAND U452 ( .A(n357), .B(n356), .Z(n358) );
  NAND U453 ( .A(n359), .B(n358), .Z(n360) );
  XOR U454 ( .A(n361), .B(n360), .Z(c[90]) );
  XOR U455 ( .A(a[91]), .B(b[91]), .Z(n365) );
  NAND U456 ( .A(a[90]), .B(b[90]), .Z(n363) );
  NAND U457 ( .A(n361), .B(n360), .Z(n362) );
  NAND U458 ( .A(n363), .B(n362), .Z(n364) );
  XOR U459 ( .A(n365), .B(n364), .Z(c[91]) );
  XOR U460 ( .A(a[92]), .B(b[92]), .Z(n369) );
  NAND U461 ( .A(a[91]), .B(b[91]), .Z(n367) );
  NAND U462 ( .A(n365), .B(n364), .Z(n366) );
  NAND U463 ( .A(n367), .B(n366), .Z(n368) );
  XOR U464 ( .A(n369), .B(n368), .Z(c[92]) );
  XOR U465 ( .A(a[93]), .B(b[93]), .Z(n373) );
  NAND U466 ( .A(a[92]), .B(b[92]), .Z(n371) );
  NAND U467 ( .A(n369), .B(n368), .Z(n370) );
  NAND U468 ( .A(n371), .B(n370), .Z(n372) );
  XOR U469 ( .A(n373), .B(n372), .Z(c[93]) );
  XOR U470 ( .A(a[94]), .B(b[94]), .Z(n377) );
  NAND U471 ( .A(a[93]), .B(b[93]), .Z(n375) );
  NAND U472 ( .A(n373), .B(n372), .Z(n374) );
  NAND U473 ( .A(n375), .B(n374), .Z(n376) );
  XOR U474 ( .A(n377), .B(n376), .Z(c[94]) );
  XOR U475 ( .A(a[95]), .B(b[95]), .Z(n381) );
  NAND U476 ( .A(a[94]), .B(b[94]), .Z(n379) );
  NAND U477 ( .A(n377), .B(n376), .Z(n378) );
  NAND U478 ( .A(n379), .B(n378), .Z(n380) );
  XOR U479 ( .A(n381), .B(n380), .Z(c[95]) );
  XOR U480 ( .A(a[96]), .B(b[96]), .Z(n385) );
  NAND U481 ( .A(a[95]), .B(b[95]), .Z(n383) );
  NAND U482 ( .A(n381), .B(n380), .Z(n382) );
  NAND U483 ( .A(n383), .B(n382), .Z(n384) );
  XOR U484 ( .A(n385), .B(n384), .Z(c[96]) );
  XOR U485 ( .A(a[97]), .B(b[97]), .Z(n389) );
  NAND U486 ( .A(a[96]), .B(b[96]), .Z(n387) );
  NAND U487 ( .A(n385), .B(n384), .Z(n386) );
  NAND U488 ( .A(n387), .B(n386), .Z(n388) );
  XOR U489 ( .A(n389), .B(n388), .Z(c[97]) );
  XOR U490 ( .A(a[98]), .B(b[98]), .Z(n393) );
  NAND U491 ( .A(a[97]), .B(b[97]), .Z(n391) );
  NAND U492 ( .A(n389), .B(n388), .Z(n390) );
  NAND U493 ( .A(n391), .B(n390), .Z(n392) );
  XOR U494 ( .A(n393), .B(n392), .Z(c[98]) );
  XOR U495 ( .A(a[99]), .B(b[99]), .Z(n397) );
  NAND U496 ( .A(a[98]), .B(b[98]), .Z(n395) );
  NAND U497 ( .A(n393), .B(n392), .Z(n394) );
  NAND U498 ( .A(n395), .B(n394), .Z(n396) );
  XOR U499 ( .A(n397), .B(n396), .Z(c[99]) );
  XOR U500 ( .A(a[100]), .B(b[100]), .Z(n401) );
  NAND U501 ( .A(a[99]), .B(b[99]), .Z(n399) );
  NAND U502 ( .A(n397), .B(n396), .Z(n398) );
  NAND U503 ( .A(n399), .B(n398), .Z(n400) );
  XOR U504 ( .A(n401), .B(n400), .Z(c[100]) );
  XOR U505 ( .A(a[101]), .B(b[101]), .Z(n405) );
  NAND U506 ( .A(a[100]), .B(b[100]), .Z(n403) );
  NAND U507 ( .A(n401), .B(n400), .Z(n402) );
  NAND U508 ( .A(n403), .B(n402), .Z(n404) );
  XOR U509 ( .A(n405), .B(n404), .Z(c[101]) );
  XOR U510 ( .A(a[102]), .B(b[102]), .Z(n409) );
  NAND U511 ( .A(a[101]), .B(b[101]), .Z(n407) );
  NAND U512 ( .A(n405), .B(n404), .Z(n406) );
  NAND U513 ( .A(n407), .B(n406), .Z(n408) );
  XOR U514 ( .A(n409), .B(n408), .Z(c[102]) );
  XOR U515 ( .A(a[103]), .B(b[103]), .Z(n413) );
  NAND U516 ( .A(a[102]), .B(b[102]), .Z(n411) );
  NAND U517 ( .A(n409), .B(n408), .Z(n410) );
  NAND U518 ( .A(n411), .B(n410), .Z(n412) );
  XOR U519 ( .A(n413), .B(n412), .Z(c[103]) );
  XOR U520 ( .A(a[104]), .B(b[104]), .Z(n417) );
  NAND U521 ( .A(a[103]), .B(b[103]), .Z(n415) );
  NAND U522 ( .A(n413), .B(n412), .Z(n414) );
  NAND U523 ( .A(n415), .B(n414), .Z(n416) );
  XOR U524 ( .A(n417), .B(n416), .Z(c[104]) );
  XOR U525 ( .A(a[105]), .B(b[105]), .Z(n421) );
  NAND U526 ( .A(a[104]), .B(b[104]), .Z(n419) );
  NAND U527 ( .A(n417), .B(n416), .Z(n418) );
  NAND U528 ( .A(n419), .B(n418), .Z(n420) );
  XOR U529 ( .A(n421), .B(n420), .Z(c[105]) );
  XOR U530 ( .A(a[106]), .B(b[106]), .Z(n425) );
  NAND U531 ( .A(a[105]), .B(b[105]), .Z(n423) );
  NAND U532 ( .A(n421), .B(n420), .Z(n422) );
  NAND U533 ( .A(n423), .B(n422), .Z(n424) );
  XOR U534 ( .A(n425), .B(n424), .Z(c[106]) );
  XOR U535 ( .A(a[107]), .B(b[107]), .Z(n429) );
  NAND U536 ( .A(a[106]), .B(b[106]), .Z(n427) );
  NAND U537 ( .A(n425), .B(n424), .Z(n426) );
  NAND U538 ( .A(n427), .B(n426), .Z(n428) );
  XOR U539 ( .A(n429), .B(n428), .Z(c[107]) );
  XOR U540 ( .A(a[108]), .B(b[108]), .Z(n433) );
  NAND U541 ( .A(a[107]), .B(b[107]), .Z(n431) );
  NAND U542 ( .A(n429), .B(n428), .Z(n430) );
  NAND U543 ( .A(n431), .B(n430), .Z(n432) );
  XOR U544 ( .A(n433), .B(n432), .Z(c[108]) );
  XOR U545 ( .A(a[109]), .B(b[109]), .Z(n437) );
  NAND U546 ( .A(a[108]), .B(b[108]), .Z(n435) );
  NAND U547 ( .A(n433), .B(n432), .Z(n434) );
  NAND U548 ( .A(n435), .B(n434), .Z(n436) );
  XOR U549 ( .A(n437), .B(n436), .Z(c[109]) );
  XOR U550 ( .A(a[110]), .B(b[110]), .Z(n441) );
  NAND U551 ( .A(a[109]), .B(b[109]), .Z(n439) );
  NAND U552 ( .A(n437), .B(n436), .Z(n438) );
  NAND U553 ( .A(n439), .B(n438), .Z(n440) );
  XOR U554 ( .A(n441), .B(n440), .Z(c[110]) );
  XOR U555 ( .A(a[111]), .B(b[111]), .Z(n445) );
  NAND U556 ( .A(a[110]), .B(b[110]), .Z(n443) );
  NAND U557 ( .A(n441), .B(n440), .Z(n442) );
  NAND U558 ( .A(n443), .B(n442), .Z(n444) );
  XOR U559 ( .A(n445), .B(n444), .Z(c[111]) );
  XOR U560 ( .A(a[112]), .B(b[112]), .Z(n449) );
  NAND U561 ( .A(a[111]), .B(b[111]), .Z(n447) );
  NAND U562 ( .A(n445), .B(n444), .Z(n446) );
  NAND U563 ( .A(n447), .B(n446), .Z(n448) );
  XOR U564 ( .A(n449), .B(n448), .Z(c[112]) );
  XOR U565 ( .A(a[113]), .B(b[113]), .Z(n453) );
  NAND U566 ( .A(a[112]), .B(b[112]), .Z(n451) );
  NAND U567 ( .A(n449), .B(n448), .Z(n450) );
  NAND U568 ( .A(n451), .B(n450), .Z(n452) );
  XOR U569 ( .A(n453), .B(n452), .Z(c[113]) );
  XOR U570 ( .A(a[114]), .B(b[114]), .Z(n457) );
  NAND U571 ( .A(a[113]), .B(b[113]), .Z(n455) );
  NAND U572 ( .A(n453), .B(n452), .Z(n454) );
  NAND U573 ( .A(n455), .B(n454), .Z(n456) );
  XOR U574 ( .A(n457), .B(n456), .Z(c[114]) );
  XOR U575 ( .A(a[115]), .B(b[115]), .Z(n461) );
  NAND U576 ( .A(a[114]), .B(b[114]), .Z(n459) );
  NAND U577 ( .A(n457), .B(n456), .Z(n458) );
  NAND U578 ( .A(n459), .B(n458), .Z(n460) );
  XOR U579 ( .A(n461), .B(n460), .Z(c[115]) );
  XOR U580 ( .A(a[116]), .B(b[116]), .Z(n465) );
  NAND U581 ( .A(a[115]), .B(b[115]), .Z(n463) );
  NAND U582 ( .A(n461), .B(n460), .Z(n462) );
  NAND U583 ( .A(n463), .B(n462), .Z(n464) );
  XOR U584 ( .A(n465), .B(n464), .Z(c[116]) );
  XOR U585 ( .A(a[117]), .B(b[117]), .Z(n469) );
  NAND U586 ( .A(a[116]), .B(b[116]), .Z(n467) );
  NAND U587 ( .A(n465), .B(n464), .Z(n466) );
  NAND U588 ( .A(n467), .B(n466), .Z(n468) );
  XOR U589 ( .A(n469), .B(n468), .Z(c[117]) );
  XOR U590 ( .A(a[118]), .B(b[118]), .Z(n473) );
  NAND U591 ( .A(a[117]), .B(b[117]), .Z(n471) );
  NAND U592 ( .A(n469), .B(n468), .Z(n470) );
  NAND U593 ( .A(n471), .B(n470), .Z(n472) );
  XOR U594 ( .A(n473), .B(n472), .Z(c[118]) );
  XOR U595 ( .A(a[119]), .B(b[119]), .Z(n477) );
  NAND U596 ( .A(a[118]), .B(b[118]), .Z(n475) );
  NAND U597 ( .A(n473), .B(n472), .Z(n474) );
  NAND U598 ( .A(n475), .B(n474), .Z(n476) );
  XOR U599 ( .A(n477), .B(n476), .Z(c[119]) );
  XOR U600 ( .A(a[120]), .B(b[120]), .Z(n481) );
  NAND U601 ( .A(a[119]), .B(b[119]), .Z(n479) );
  NAND U602 ( .A(n477), .B(n476), .Z(n478) );
  NAND U603 ( .A(n479), .B(n478), .Z(n480) );
  XOR U604 ( .A(n481), .B(n480), .Z(c[120]) );
  XOR U605 ( .A(a[121]), .B(b[121]), .Z(n485) );
  NAND U606 ( .A(a[120]), .B(b[120]), .Z(n483) );
  NAND U607 ( .A(n481), .B(n480), .Z(n482) );
  NAND U608 ( .A(n483), .B(n482), .Z(n484) );
  XOR U609 ( .A(n485), .B(n484), .Z(c[121]) );
  XOR U610 ( .A(a[122]), .B(b[122]), .Z(n489) );
  NAND U611 ( .A(a[121]), .B(b[121]), .Z(n487) );
  NAND U612 ( .A(n485), .B(n484), .Z(n486) );
  NAND U613 ( .A(n487), .B(n486), .Z(n488) );
  XOR U614 ( .A(n489), .B(n488), .Z(c[122]) );
  XOR U615 ( .A(a[123]), .B(b[123]), .Z(n493) );
  NAND U616 ( .A(a[122]), .B(b[122]), .Z(n491) );
  NAND U617 ( .A(n489), .B(n488), .Z(n490) );
  NAND U618 ( .A(n491), .B(n490), .Z(n492) );
  XOR U619 ( .A(n493), .B(n492), .Z(c[123]) );
  XOR U620 ( .A(a[124]), .B(b[124]), .Z(n497) );
  NAND U621 ( .A(a[123]), .B(b[123]), .Z(n495) );
  NAND U622 ( .A(n493), .B(n492), .Z(n494) );
  NAND U623 ( .A(n495), .B(n494), .Z(n496) );
  XOR U624 ( .A(n497), .B(n496), .Z(c[124]) );
  XOR U625 ( .A(a[125]), .B(b[125]), .Z(n501) );
  NAND U626 ( .A(a[124]), .B(b[124]), .Z(n499) );
  NAND U627 ( .A(n497), .B(n496), .Z(n498) );
  NAND U628 ( .A(n499), .B(n498), .Z(n500) );
  XOR U629 ( .A(n501), .B(n500), .Z(c[125]) );
  XOR U630 ( .A(a[126]), .B(b[126]), .Z(n505) );
  NAND U631 ( .A(a[125]), .B(b[125]), .Z(n503) );
  NAND U632 ( .A(n501), .B(n500), .Z(n502) );
  NAND U633 ( .A(n503), .B(n502), .Z(n504) );
  XOR U634 ( .A(n505), .B(n504), .Z(c[126]) );
  NAND U635 ( .A(a[126]), .B(b[126]), .Z(n507) );
  NAND U636 ( .A(n505), .B(n504), .Z(n506) );
  AND U637 ( .A(n507), .B(n506), .Z(n509) );
  XOR U638 ( .A(a[127]), .B(b[127]), .Z(n508) );
  XNOR U639 ( .A(n509), .B(n508), .Z(c[127]) );
  NAND U640 ( .A(a[127]), .B(b[127]), .Z(n511) );
  NANDN U641 ( .A(n509), .B(n508), .Z(n510) );
  NAND U642 ( .A(n511), .B(n510), .Z(carry_on_d) );
endmodule

