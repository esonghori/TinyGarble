
module aes_seq_CC5 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [255:0] key;
  output [127:0] out;
  input clk, rst;
  wire   \w0[1][127] , \w0[1][126] , \w0[1][125] , \w0[1][124] , \w0[1][123] ,
         \w0[1][122] , \w0[1][121] , \w0[1][120] , \w0[1][119] , \w0[1][118] ,
         \w0[1][117] , \w0[1][116] , \w0[1][115] , \w0[1][114] , \w0[1][113] ,
         \w0[1][112] , \w0[1][111] , \w0[1][110] , \w0[1][109] , \w0[1][108] ,
         \w0[1][107] , \w0[1][106] , \w0[1][105] , \w0[1][104] , \w0[1][103] ,
         \w0[1][102] , \w0[1][101] , \w0[1][100] , \w0[1][99] , \w0[1][98] ,
         \w0[1][97] , \w0[1][96] , \w0[1][95] , \w0[1][94] , \w0[1][93] ,
         \w0[1][92] , \w0[1][91] , \w0[1][90] , \w0[1][89] , \w0[1][88] ,
         \w0[1][87] , \w0[1][86] , \w0[1][85] , \w0[1][84] , \w0[1][83] ,
         \w0[1][82] , \w0[1][81] , \w0[1][80] , \w0[1][79] , \w0[1][78] ,
         \w0[1][77] , \w0[1][76] , \w0[1][75] , \w0[1][74] , \w0[1][73] ,
         \w0[1][72] , \w0[1][71] , \w0[1][70] , \w0[1][69] , \w0[1][68] ,
         \w0[1][67] , \w0[1][66] , \w0[1][65] , \w0[1][64] , \w0[1][63] ,
         \w0[1][62] , \w0[1][61] , \w0[1][60] , \w0[1][59] , \w0[1][58] ,
         \w0[1][57] , \w0[1][56] , \w0[1][55] , \w0[1][54] , \w0[1][53] ,
         \w0[1][52] , \w0[1][51] , \w0[1][50] , \w0[1][49] , \w0[1][48] ,
         \w0[1][47] , \w0[1][46] , \w0[1][45] , \w0[1][44] , \w0[1][43] ,
         \w0[1][42] , \w0[1][41] , \w0[1][40] , \w0[1][39] , \w0[1][38] ,
         \w0[1][37] , \w0[1][36] , \w0[1][35] , \w0[1][34] , \w0[1][33] ,
         \w0[1][32] , \w0[1][31] , \w0[1][30] , \w0[1][29] , \w0[1][28] ,
         \w0[1][27] , \w0[1][26] , \w0[1][25] , \w0[1][24] , \w0[1][23] ,
         \w0[1][22] , \w0[1][21] , \w0[1][20] , \w0[1][19] , \w0[1][18] ,
         \w0[1][17] , \w0[1][16] , \w0[1][15] , \w0[1][14] , \w0[1][13] ,
         \w0[1][12] , \w0[1][11] , \w0[1][10] , \w0[1][9] , \w0[1][8] ,
         \w0[1][7] , \w0[1][6] , \w0[1][5] , \w0[1][4] , \w0[1][3] ,
         \w0[1][2] , \w0[1][1] , \w0[1][0] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394;
  wire   [127:0] state;

  DFF \state_reg[0]  ( .D(\w0[1][0] ), .CLK(clk), .RST(rst), .I(msg[0]), .Q(
        state[0]) );
  DFF \state_reg[1]  ( .D(\w0[1][1] ), .CLK(clk), .RST(rst), .I(msg[1]), .Q(
        state[1]) );
  DFF \state_reg[2]  ( .D(\w0[1][2] ), .CLK(clk), .RST(rst), .I(msg[2]), .Q(
        state[2]) );
  DFF \state_reg[3]  ( .D(\w0[1][3] ), .CLK(clk), .RST(rst), .I(msg[3]), .Q(
        state[3]) );
  DFF \state_reg[4]  ( .D(\w0[1][4] ), .CLK(clk), .RST(rst), .I(msg[4]), .Q(
        state[4]) );
  DFF \state_reg[5]  ( .D(\w0[1][5] ), .CLK(clk), .RST(rst), .I(msg[5]), .Q(
        state[5]) );
  DFF \state_reg[6]  ( .D(\w0[1][6] ), .CLK(clk), .RST(rst), .I(msg[6]), .Q(
        state[6]) );
  DFF \state_reg[7]  ( .D(\w0[1][7] ), .CLK(clk), .RST(rst), .I(msg[7]), .Q(
        state[7]) );
  DFF \state_reg[8]  ( .D(\w0[1][8] ), .CLK(clk), .RST(rst), .I(msg[8]), .Q(
        state[8]) );
  DFF \state_reg[9]  ( .D(\w0[1][9] ), .CLK(clk), .RST(rst), .I(msg[9]), .Q(
        state[9]) );
  DFF \state_reg[10]  ( .D(\w0[1][10] ), .CLK(clk), .RST(rst), .I(msg[10]), 
        .Q(state[10]) );
  DFF \state_reg[11]  ( .D(\w0[1][11] ), .CLK(clk), .RST(rst), .I(msg[11]), 
        .Q(state[11]) );
  DFF \state_reg[12]  ( .D(\w0[1][12] ), .CLK(clk), .RST(rst), .I(msg[12]), 
        .Q(state[12]) );
  DFF \state_reg[13]  ( .D(\w0[1][13] ), .CLK(clk), .RST(rst), .I(msg[13]), 
        .Q(state[13]) );
  DFF \state_reg[14]  ( .D(\w0[1][14] ), .CLK(clk), .RST(rst), .I(msg[14]), 
        .Q(state[14]) );
  DFF \state_reg[15]  ( .D(\w0[1][15] ), .CLK(clk), .RST(rst), .I(msg[15]), 
        .Q(state[15]) );
  DFF \state_reg[16]  ( .D(\w0[1][16] ), .CLK(clk), .RST(rst), .I(msg[16]), 
        .Q(state[16]) );
  DFF \state_reg[17]  ( .D(\w0[1][17] ), .CLK(clk), .RST(rst), .I(msg[17]), 
        .Q(state[17]) );
  DFF \state_reg[18]  ( .D(\w0[1][18] ), .CLK(clk), .RST(rst), .I(msg[18]), 
        .Q(state[18]) );
  DFF \state_reg[19]  ( .D(\w0[1][19] ), .CLK(clk), .RST(rst), .I(msg[19]), 
        .Q(state[19]) );
  DFF \state_reg[20]  ( .D(\w0[1][20] ), .CLK(clk), .RST(rst), .I(msg[20]), 
        .Q(state[20]) );
  DFF \state_reg[21]  ( .D(\w0[1][21] ), .CLK(clk), .RST(rst), .I(msg[21]), 
        .Q(state[21]) );
  DFF \state_reg[22]  ( .D(\w0[1][22] ), .CLK(clk), .RST(rst), .I(msg[22]), 
        .Q(state[22]) );
  DFF \state_reg[23]  ( .D(\w0[1][23] ), .CLK(clk), .RST(rst), .I(msg[23]), 
        .Q(state[23]) );
  DFF \state_reg[24]  ( .D(\w0[1][24] ), .CLK(clk), .RST(rst), .I(msg[24]), 
        .Q(state[24]) );
  DFF \state_reg[25]  ( .D(\w0[1][25] ), .CLK(clk), .RST(rst), .I(msg[25]), 
        .Q(state[25]) );
  DFF \state_reg[26]  ( .D(\w0[1][26] ), .CLK(clk), .RST(rst), .I(msg[26]), 
        .Q(state[26]) );
  DFF \state_reg[27]  ( .D(\w0[1][27] ), .CLK(clk), .RST(rst), .I(msg[27]), 
        .Q(state[27]) );
  DFF \state_reg[28]  ( .D(\w0[1][28] ), .CLK(clk), .RST(rst), .I(msg[28]), 
        .Q(state[28]) );
  DFF \state_reg[29]  ( .D(\w0[1][29] ), .CLK(clk), .RST(rst), .I(msg[29]), 
        .Q(state[29]) );
  DFF \state_reg[30]  ( .D(\w0[1][30] ), .CLK(clk), .RST(rst), .I(msg[30]), 
        .Q(state[30]) );
  DFF \state_reg[31]  ( .D(\w0[1][31] ), .CLK(clk), .RST(rst), .I(msg[31]), 
        .Q(state[31]) );
  DFF \state_reg[32]  ( .D(\w0[1][32] ), .CLK(clk), .RST(rst), .I(msg[32]), 
        .Q(state[32]) );
  DFF \state_reg[33]  ( .D(\w0[1][33] ), .CLK(clk), .RST(rst), .I(msg[33]), 
        .Q(state[33]) );
  DFF \state_reg[34]  ( .D(\w0[1][34] ), .CLK(clk), .RST(rst), .I(msg[34]), 
        .Q(state[34]) );
  DFF \state_reg[35]  ( .D(\w0[1][35] ), .CLK(clk), .RST(rst), .I(msg[35]), 
        .Q(state[35]) );
  DFF \state_reg[36]  ( .D(\w0[1][36] ), .CLK(clk), .RST(rst), .I(msg[36]), 
        .Q(state[36]) );
  DFF \state_reg[37]  ( .D(\w0[1][37] ), .CLK(clk), .RST(rst), .I(msg[37]), 
        .Q(state[37]) );
  DFF \state_reg[38]  ( .D(\w0[1][38] ), .CLK(clk), .RST(rst), .I(msg[38]), 
        .Q(state[38]) );
  DFF \state_reg[39]  ( .D(\w0[1][39] ), .CLK(clk), .RST(rst), .I(msg[39]), 
        .Q(state[39]) );
  DFF \state_reg[40]  ( .D(\w0[1][40] ), .CLK(clk), .RST(rst), .I(msg[40]), 
        .Q(state[40]) );
  DFF \state_reg[41]  ( .D(\w0[1][41] ), .CLK(clk), .RST(rst), .I(msg[41]), 
        .Q(state[41]) );
  DFF \state_reg[42]  ( .D(\w0[1][42] ), .CLK(clk), .RST(rst), .I(msg[42]), 
        .Q(state[42]) );
  DFF \state_reg[43]  ( .D(\w0[1][43] ), .CLK(clk), .RST(rst), .I(msg[43]), 
        .Q(state[43]) );
  DFF \state_reg[44]  ( .D(\w0[1][44] ), .CLK(clk), .RST(rst), .I(msg[44]), 
        .Q(state[44]) );
  DFF \state_reg[45]  ( .D(\w0[1][45] ), .CLK(clk), .RST(rst), .I(msg[45]), 
        .Q(state[45]) );
  DFF \state_reg[46]  ( .D(\w0[1][46] ), .CLK(clk), .RST(rst), .I(msg[46]), 
        .Q(state[46]) );
  DFF \state_reg[47]  ( .D(\w0[1][47] ), .CLK(clk), .RST(rst), .I(msg[47]), 
        .Q(state[47]) );
  DFF \state_reg[48]  ( .D(\w0[1][48] ), .CLK(clk), .RST(rst), .I(msg[48]), 
        .Q(state[48]) );
  DFF \state_reg[49]  ( .D(\w0[1][49] ), .CLK(clk), .RST(rst), .I(msg[49]), 
        .Q(state[49]) );
  DFF \state_reg[50]  ( .D(\w0[1][50] ), .CLK(clk), .RST(rst), .I(msg[50]), 
        .Q(state[50]) );
  DFF \state_reg[51]  ( .D(\w0[1][51] ), .CLK(clk), .RST(rst), .I(msg[51]), 
        .Q(state[51]) );
  DFF \state_reg[52]  ( .D(\w0[1][52] ), .CLK(clk), .RST(rst), .I(msg[52]), 
        .Q(state[52]) );
  DFF \state_reg[53]  ( .D(\w0[1][53] ), .CLK(clk), .RST(rst), .I(msg[53]), 
        .Q(state[53]) );
  DFF \state_reg[54]  ( .D(\w0[1][54] ), .CLK(clk), .RST(rst), .I(msg[54]), 
        .Q(state[54]) );
  DFF \state_reg[55]  ( .D(\w0[1][55] ), .CLK(clk), .RST(rst), .I(msg[55]), 
        .Q(state[55]) );
  DFF \state_reg[56]  ( .D(\w0[1][56] ), .CLK(clk), .RST(rst), .I(msg[56]), 
        .Q(state[56]) );
  DFF \state_reg[57]  ( .D(\w0[1][57] ), .CLK(clk), .RST(rst), .I(msg[57]), 
        .Q(state[57]) );
  DFF \state_reg[58]  ( .D(\w0[1][58] ), .CLK(clk), .RST(rst), .I(msg[58]), 
        .Q(state[58]) );
  DFF \state_reg[59]  ( .D(\w0[1][59] ), .CLK(clk), .RST(rst), .I(msg[59]), 
        .Q(state[59]) );
  DFF \state_reg[60]  ( .D(\w0[1][60] ), .CLK(clk), .RST(rst), .I(msg[60]), 
        .Q(state[60]) );
  DFF \state_reg[61]  ( .D(\w0[1][61] ), .CLK(clk), .RST(rst), .I(msg[61]), 
        .Q(state[61]) );
  DFF \state_reg[62]  ( .D(\w0[1][62] ), .CLK(clk), .RST(rst), .I(msg[62]), 
        .Q(state[62]) );
  DFF \state_reg[63]  ( .D(\w0[1][63] ), .CLK(clk), .RST(rst), .I(msg[63]), 
        .Q(state[63]) );
  DFF \state_reg[64]  ( .D(\w0[1][64] ), .CLK(clk), .RST(rst), .I(msg[64]), 
        .Q(state[64]) );
  DFF \state_reg[65]  ( .D(\w0[1][65] ), .CLK(clk), .RST(rst), .I(msg[65]), 
        .Q(state[65]) );
  DFF \state_reg[66]  ( .D(\w0[1][66] ), .CLK(clk), .RST(rst), .I(msg[66]), 
        .Q(state[66]) );
  DFF \state_reg[67]  ( .D(\w0[1][67] ), .CLK(clk), .RST(rst), .I(msg[67]), 
        .Q(state[67]) );
  DFF \state_reg[68]  ( .D(\w0[1][68] ), .CLK(clk), .RST(rst), .I(msg[68]), 
        .Q(state[68]) );
  DFF \state_reg[69]  ( .D(\w0[1][69] ), .CLK(clk), .RST(rst), .I(msg[69]), 
        .Q(state[69]) );
  DFF \state_reg[70]  ( .D(\w0[1][70] ), .CLK(clk), .RST(rst), .I(msg[70]), 
        .Q(state[70]) );
  DFF \state_reg[71]  ( .D(\w0[1][71] ), .CLK(clk), .RST(rst), .I(msg[71]), 
        .Q(state[71]) );
  DFF \state_reg[72]  ( .D(\w0[1][72] ), .CLK(clk), .RST(rst), .I(msg[72]), 
        .Q(state[72]) );
  DFF \state_reg[73]  ( .D(\w0[1][73] ), .CLK(clk), .RST(rst), .I(msg[73]), 
        .Q(state[73]) );
  DFF \state_reg[74]  ( .D(\w0[1][74] ), .CLK(clk), .RST(rst), .I(msg[74]), 
        .Q(state[74]) );
  DFF \state_reg[75]  ( .D(\w0[1][75] ), .CLK(clk), .RST(rst), .I(msg[75]), 
        .Q(state[75]) );
  DFF \state_reg[76]  ( .D(\w0[1][76] ), .CLK(clk), .RST(rst), .I(msg[76]), 
        .Q(state[76]) );
  DFF \state_reg[77]  ( .D(\w0[1][77] ), .CLK(clk), .RST(rst), .I(msg[77]), 
        .Q(state[77]) );
  DFF \state_reg[78]  ( .D(\w0[1][78] ), .CLK(clk), .RST(rst), .I(msg[78]), 
        .Q(state[78]) );
  DFF \state_reg[79]  ( .D(\w0[1][79] ), .CLK(clk), .RST(rst), .I(msg[79]), 
        .Q(state[79]) );
  DFF \state_reg[80]  ( .D(\w0[1][80] ), .CLK(clk), .RST(rst), .I(msg[80]), 
        .Q(state[80]) );
  DFF \state_reg[81]  ( .D(\w0[1][81] ), .CLK(clk), .RST(rst), .I(msg[81]), 
        .Q(state[81]) );
  DFF \state_reg[82]  ( .D(\w0[1][82] ), .CLK(clk), .RST(rst), .I(msg[82]), 
        .Q(state[82]) );
  DFF \state_reg[83]  ( .D(\w0[1][83] ), .CLK(clk), .RST(rst), .I(msg[83]), 
        .Q(state[83]) );
  DFF \state_reg[84]  ( .D(\w0[1][84] ), .CLK(clk), .RST(rst), .I(msg[84]), 
        .Q(state[84]) );
  DFF \state_reg[85]  ( .D(\w0[1][85] ), .CLK(clk), .RST(rst), .I(msg[85]), 
        .Q(state[85]) );
  DFF \state_reg[86]  ( .D(\w0[1][86] ), .CLK(clk), .RST(rst), .I(msg[86]), 
        .Q(state[86]) );
  DFF \state_reg[87]  ( .D(\w0[1][87] ), .CLK(clk), .RST(rst), .I(msg[87]), 
        .Q(state[87]) );
  DFF \state_reg[88]  ( .D(\w0[1][88] ), .CLK(clk), .RST(rst), .I(msg[88]), 
        .Q(state[88]) );
  DFF \state_reg[89]  ( .D(\w0[1][89] ), .CLK(clk), .RST(rst), .I(msg[89]), 
        .Q(state[89]) );
  DFF \state_reg[90]  ( .D(\w0[1][90] ), .CLK(clk), .RST(rst), .I(msg[90]), 
        .Q(state[90]) );
  DFF \state_reg[91]  ( .D(\w0[1][91] ), .CLK(clk), .RST(rst), .I(msg[91]), 
        .Q(state[91]) );
  DFF \state_reg[92]  ( .D(\w0[1][92] ), .CLK(clk), .RST(rst), .I(msg[92]), 
        .Q(state[92]) );
  DFF \state_reg[93]  ( .D(\w0[1][93] ), .CLK(clk), .RST(rst), .I(msg[93]), 
        .Q(state[93]) );
  DFF \state_reg[94]  ( .D(\w0[1][94] ), .CLK(clk), .RST(rst), .I(msg[94]), 
        .Q(state[94]) );
  DFF \state_reg[95]  ( .D(\w0[1][95] ), .CLK(clk), .RST(rst), .I(msg[95]), 
        .Q(state[95]) );
  DFF \state_reg[96]  ( .D(\w0[1][96] ), .CLK(clk), .RST(rst), .I(msg[96]), 
        .Q(state[96]) );
  DFF \state_reg[97]  ( .D(\w0[1][97] ), .CLK(clk), .RST(rst), .I(msg[97]), 
        .Q(state[97]) );
  DFF \state_reg[98]  ( .D(\w0[1][98] ), .CLK(clk), .RST(rst), .I(msg[98]), 
        .Q(state[98]) );
  DFF \state_reg[99]  ( .D(\w0[1][99] ), .CLK(clk), .RST(rst), .I(msg[99]), 
        .Q(state[99]) );
  DFF \state_reg[100]  ( .D(\w0[1][100] ), .CLK(clk), .RST(rst), .I(msg[100]), 
        .Q(state[100]) );
  DFF \state_reg[101]  ( .D(\w0[1][101] ), .CLK(clk), .RST(rst), .I(msg[101]), 
        .Q(state[101]) );
  DFF \state_reg[102]  ( .D(\w0[1][102] ), .CLK(clk), .RST(rst), .I(msg[102]), 
        .Q(state[102]) );
  DFF \state_reg[103]  ( .D(\w0[1][103] ), .CLK(clk), .RST(rst), .I(msg[103]), 
        .Q(state[103]) );
  DFF \state_reg[104]  ( .D(\w0[1][104] ), .CLK(clk), .RST(rst), .I(msg[104]), 
        .Q(state[104]) );
  DFF \state_reg[105]  ( .D(\w0[1][105] ), .CLK(clk), .RST(rst), .I(msg[105]), 
        .Q(state[105]) );
  DFF \state_reg[106]  ( .D(\w0[1][106] ), .CLK(clk), .RST(rst), .I(msg[106]), 
        .Q(state[106]) );
  DFF \state_reg[107]  ( .D(\w0[1][107] ), .CLK(clk), .RST(rst), .I(msg[107]), 
        .Q(state[107]) );
  DFF \state_reg[108]  ( .D(\w0[1][108] ), .CLK(clk), .RST(rst), .I(msg[108]), 
        .Q(state[108]) );
  DFF \state_reg[109]  ( .D(\w0[1][109] ), .CLK(clk), .RST(rst), .I(msg[109]), 
        .Q(state[109]) );
  DFF \state_reg[110]  ( .D(\w0[1][110] ), .CLK(clk), .RST(rst), .I(msg[110]), 
        .Q(state[110]) );
  DFF \state_reg[111]  ( .D(\w0[1][111] ), .CLK(clk), .RST(rst), .I(msg[111]), 
        .Q(state[111]) );
  DFF \state_reg[112]  ( .D(\w0[1][112] ), .CLK(clk), .RST(rst), .I(msg[112]), 
        .Q(state[112]) );
  DFF \state_reg[113]  ( .D(\w0[1][113] ), .CLK(clk), .RST(rst), .I(msg[113]), 
        .Q(state[113]) );
  DFF \state_reg[114]  ( .D(\w0[1][114] ), .CLK(clk), .RST(rst), .I(msg[114]), 
        .Q(state[114]) );
  DFF \state_reg[115]  ( .D(\w0[1][115] ), .CLK(clk), .RST(rst), .I(msg[115]), 
        .Q(state[115]) );
  DFF \state_reg[116]  ( .D(\w0[1][116] ), .CLK(clk), .RST(rst), .I(msg[116]), 
        .Q(state[116]) );
  DFF \state_reg[117]  ( .D(\w0[1][117] ), .CLK(clk), .RST(rst), .I(msg[117]), 
        .Q(state[117]) );
  DFF \state_reg[118]  ( .D(\w0[1][118] ), .CLK(clk), .RST(rst), .I(msg[118]), 
        .Q(state[118]) );
  DFF \state_reg[119]  ( .D(\w0[1][119] ), .CLK(clk), .RST(rst), .I(msg[119]), 
        .Q(state[119]) );
  DFF \state_reg[120]  ( .D(\w0[1][120] ), .CLK(clk), .RST(rst), .I(msg[120]), 
        .Q(state[120]) );
  DFF \state_reg[121]  ( .D(\w0[1][121] ), .CLK(clk), .RST(rst), .I(msg[121]), 
        .Q(state[121]) );
  DFF \state_reg[122]  ( .D(\w0[1][122] ), .CLK(clk), .RST(rst), .I(msg[122]), 
        .Q(state[122]) );
  DFF \state_reg[123]  ( .D(\w0[1][123] ), .CLK(clk), .RST(rst), .I(msg[123]), 
        .Q(state[123]) );
  DFF \state_reg[124]  ( .D(\w0[1][124] ), .CLK(clk), .RST(rst), .I(msg[124]), 
        .Q(state[124]) );
  DFF \state_reg[125]  ( .D(\w0[1][125] ), .CLK(clk), .RST(rst), .I(msg[125]), 
        .Q(state[125]) );
  DFF \state_reg[126]  ( .D(\w0[1][126] ), .CLK(clk), .RST(rst), .I(msg[126]), 
        .Q(state[126]) );
  DFF \state_reg[127]  ( .D(\w0[1][127] ), .CLK(clk), .RST(rst), .I(msg[127]), 
        .Q(state[127]) );
  XNOR U3 ( .A(n3700), .B(n3690), .Z(n3697) );
  XNOR U4 ( .A(n5019), .B(n5010), .Z(n5017) );
  XNOR U5 ( .A(n2785), .B(n2776), .Z(n2783) );
  XNOR U6 ( .A(n2678), .B(n2669), .Z(n2676) );
  XNOR U7 ( .A(n2476), .B(n2466), .Z(n2474) );
  XNOR U8 ( .A(n3462), .B(n3453), .Z(n3460) );
  XNOR U9 ( .A(n3580), .B(n3571), .Z(n3578) );
  XOR U10 ( .A(n5323), .B(n5337), .Z(n5334) );
  XNOR U11 ( .A(n4337), .B(n4327), .Z(n4334) );
  XNOR U12 ( .A(n4545), .B(n4535), .Z(n4542) );
  XNOR U13 ( .A(n2139), .B(n2096), .Z(n2193) );
  XOR U14 ( .A(n4465), .B(n4472), .Z(n4471) );
  XOR U15 ( .A(n2564), .B(n2551), .Z(n2354) );
  XOR U16 ( .A(n3341), .B(n3332), .Z(n3216) );
  XOR U17 ( .A(n5111), .B(n5098), .Z(n4936) );
  NOR U18 ( .A(n5020), .B(n5019), .Z(n5016) );
  NOR U19 ( .A(n5332), .B(n5331), .Z(n5328) );
  XOR U20 ( .A(n5227), .B(n5214), .Z(n4915) );
  XOR U21 ( .A(n524), .B(n515), .Z(n444) );
  OR U22 ( .A(n3649), .B(n3266), .Z(n3648) );
  XNOR U23 ( .A(n4783), .B(n4896), .Z(n4798) );
  XNOR U24 ( .A(n4821), .B(n4834), .Z(n4833) );
  XOR U25 ( .A(n425), .B(n1651), .Z(n1082) );
  XNOR U26 ( .A(n785), .B(n2036), .Z(n807) );
  XNOR U27 ( .A(n2562), .B(n2553), .Z(n2560) );
  XNOR U28 ( .A(n5109), .B(n5100), .Z(n5107) );
  XNOR U29 ( .A(n5331), .B(n5322), .Z(n5329) );
  XNOR U30 ( .A(n5225), .B(n5216), .Z(n5223) );
  XOR U31 ( .A(n5011), .B(n5025), .Z(n5022) );
  XOR U32 ( .A(n4627), .B(n4638), .Z(n4635) );
  XNOR U33 ( .A(n4628), .B(n4613), .Z(n4620) );
  XNOR U34 ( .A(n1880), .B(n867), .Z(n4746) );
  XNOR U35 ( .A(n1920), .B(n1851), .Z(n1974) );
  XNOR U36 ( .A(n1710), .B(n1667), .Z(n1764) );
  XNOR U37 ( .A(n1303), .B(n1260), .Z(n1357) );
  XNOR U38 ( .A(n1110), .B(n1064), .Z(n1164) );
  XNOR U39 ( .A(n907), .B(n848), .Z(n961) );
  XNOR U40 ( .A(n292), .B(n249), .Z(n346) );
  XNOR U41 ( .A(n89), .B(n43), .Z(n143) );
  NOR U42 ( .A(n2377), .B(n2452), .Z(n2493) );
  NOR U43 ( .A(n2366), .B(n2629), .Z(n2802) );
  XOR U44 ( .A(n3726), .B(n3733), .Z(n3732) );
  XOR U45 ( .A(n4361), .B(n4368), .Z(n4367) );
  XOR U46 ( .A(n4296), .B(n4279), .Z(n4294) );
  NOR U47 ( .A(n4633), .B(n4632), .Z(n4629) );
  XOR U48 ( .A(n4569), .B(n4576), .Z(n4575) );
  XOR U49 ( .A(n4525), .B(n4309), .Z(n4523) );
  XNOR U50 ( .A(n4026), .B(n4016), .Z(n4023) );
  XNOR U51 ( .A(n2787), .B(n2774), .Z(n2365) );
  XOR U52 ( .A(n2680), .B(n2667), .Z(n2254) );
  XNOR U53 ( .A(n2478), .B(n2464), .Z(n2376) );
  XOR U54 ( .A(n3464), .B(n3451), .Z(n3224) );
  XNOR U55 ( .A(n3394), .B(n3392), .Z(n3233) );
  XOR U56 ( .A(n3582), .B(n3569), .Z(n3209) );
  XOR U57 ( .A(n4442), .B(n4433), .Z(n4187) );
  XOR U58 ( .A(n3218), .B(n3213), .Z(n3148) );
  XOR U59 ( .A(n4847), .B(n4842), .Z(n4805) );
  XNOR U60 ( .A(n4887), .B(n4991), .Z(n4837) );
  XOR U61 ( .A(n862), .B(n857), .Z(n423) );
  XOR U62 ( .A(n1846), .B(n1841), .Z(n1830) );
  XOR U63 ( .A(n1662), .B(n1657), .Z(n1645) );
  XOR U64 ( .A(n1466), .B(n1461), .Z(n1450) );
  XOR U65 ( .A(n1255), .B(n1250), .Z(n1239) );
  XOR U66 ( .A(n1059), .B(n1054), .Z(n1043) );
  XOR U67 ( .A(n843), .B(n838), .Z(n827) );
  XOR U68 ( .A(n446), .B(n441), .Z(n428) );
  XOR U69 ( .A(n244), .B(n239), .Z(n228) );
  XOR U70 ( .A(n38), .B(n33), .Z(n22) );
  XOR U71 ( .A(n3771), .B(n3766), .Z(n3061) );
  XOR U72 ( .A(n2891), .B(n2886), .Z(n2875) );
  XOR U73 ( .A(n2091), .B(n2086), .Z(n2075) );
  XNOR U74 ( .A(n2277), .B(n2742), .Z(n2445) );
  XNOR U75 ( .A(n2230), .B(n2379), .Z(n814) );
  XNOR U76 ( .A(n3275), .B(n3169), .Z(n3408) );
  XOR U77 ( .A(n3184), .B(n3183), .Z(n3182) );
  XOR U78 ( .A(n4799), .B(n4782), .Z(n4796) );
  XNOR U79 ( .A(n4815), .B(n4851), .Z(n4848) );
  XNOR U80 ( .A(n1031), .B(n405), .Z(n1022) );
  XOR U81 ( .A(n819), .B(n1408), .Z(n2237) );
  XNOR U82 ( .A(n3649), .B(n3265), .Z(n3719) );
  XOR U83 ( .A(n2777), .B(n2791), .Z(n2788) );
  XOR U84 ( .A(n2554), .B(n2568), .Z(n2565) );
  XOR U85 ( .A(n2670), .B(n2684), .Z(n2681) );
  XOR U86 ( .A(n2467), .B(n2482), .Z(n2479) );
  XOR U87 ( .A(n3454), .B(n3468), .Z(n3465) );
  XOR U88 ( .A(n3572), .B(n3586), .Z(n3583) );
  XNOR U89 ( .A(n3347), .B(n3334), .Z(n3342) );
  XOR U90 ( .A(n5101), .B(n5115), .Z(n5112) );
  XOR U91 ( .A(n5217), .B(n5231), .Z(n5228) );
  XNOR U92 ( .A(n4285), .B(n4101), .Z(n4355) );
  XNOR U93 ( .A(n4270), .B(n4264), .Z(n4268) );
  XNOR U94 ( .A(n4409), .B(n4192), .Z(n4459) );
  XNOR U95 ( .A(n4441), .B(n4431), .Z(n4438) );
  XNOR U96 ( .A(n4513), .B(n4178), .Z(n4563) );
  XNOR U97 ( .A(n2417), .B(n2401), .Z(n2415) );
  XOR U98 ( .A(n2517), .B(n2524), .Z(n2520) );
  XOR U99 ( .A(n2826), .B(n2833), .Z(n2829) );
  XNOR U100 ( .A(n2659), .B(n2644), .Z(n2657) );
  XNOR U101 ( .A(n3435), .B(n3430), .Z(n3433) );
  XNOR U102 ( .A(n3553), .B(n3548), .Z(n3551) );
  XNOR U103 ( .A(n5327), .B(n5317), .Z(n5319) );
  XNOR U104 ( .A(n4963), .B(n4947), .Z(n4961) );
  XNOR U105 ( .A(n4990), .B(n4973), .Z(n4988) );
  XNOR U106 ( .A(n5221), .B(n5211), .Z(n5213) );
  XNOR U107 ( .A(n4721), .B(n4711), .Z(n4718) );
  XNOR U108 ( .A(n1950), .B(n1940), .Z(n1947) );
  XNOR U109 ( .A(n1740), .B(n1730), .Z(n1737) );
  XNOR U110 ( .A(n1544), .B(n1534), .Z(n1541) );
  XNOR U111 ( .A(n1333), .B(n1323), .Z(n1330) );
  XNOR U112 ( .A(n1140), .B(n1130), .Z(n1137) );
  XNOR U113 ( .A(n937), .B(n927), .Z(n934) );
  XNOR U114 ( .A(n780), .B(n800), .Z(n777) );
  XNOR U115 ( .A(n656), .B(n692), .Z(n686) );
  XNOR U116 ( .A(n322), .B(n312), .Z(n319) );
  XNOR U117 ( .A(n119), .B(n109), .Z(n116) );
  XNOR U118 ( .A(n3849), .B(n3839), .Z(n3846) );
  XNOR U119 ( .A(n2969), .B(n2959), .Z(n2966) );
  XNOR U120 ( .A(n2169), .B(n2159), .Z(n2166) );
  NOR U121 ( .A(n2477), .B(n2476), .Z(n2473) );
  NOR U122 ( .A(n2786), .B(n2785), .Z(n2782) );
  NOR U123 ( .A(n2563), .B(n2562), .Z(n2559) );
  NOR U124 ( .A(n2679), .B(n2678), .Z(n2675) );
  NOR U125 ( .A(n3463), .B(n3462), .Z(n3459) );
  XOR U126 ( .A(n3701), .B(n3692), .Z(n3654) );
  NOR U127 ( .A(n3581), .B(n3580), .Z(n3577) );
  NOR U128 ( .A(n5110), .B(n5109), .Z(n5106) );
  XOR U129 ( .A(n5333), .B(n5320), .Z(n4828) );
  NOR U130 ( .A(n5226), .B(n5225), .Z(n5222) );
  XOR U131 ( .A(n5021), .B(n5008), .Z(n4926) );
  XOR U132 ( .A(n4338), .B(n4329), .Z(n4152) );
  XNOR U133 ( .A(n4675), .B(n4673), .Z(n4255) );
  XOR U134 ( .A(n4546), .B(n4537), .Z(n4172) );
  XOR U135 ( .A(n4634), .B(n4625), .Z(n4208) );
  NANDN U136 ( .A(n4700), .B(n1442), .Z(n1878) );
  NANDN U137 ( .A(n3070), .B(n2850), .Z(n2064) );
  XOR U138 ( .A(n3090), .B(n3081), .Z(n2053) );
  NANDN U139 ( .A(n1929), .B(n1887), .Z(n1918) );
  NANDN U140 ( .A(n1719), .B(n1677), .Z(n1708) );
  NANDN U141 ( .A(n1523), .B(n1481), .Z(n1512) );
  NANDN U142 ( .A(n1312), .B(n1270), .Z(n1301) );
  NANDN U143 ( .A(n1119), .B(n1074), .Z(n1108) );
  NANDN U144 ( .A(n916), .B(n874), .Z(n905) );
  XOR U145 ( .A(n727), .B(n718), .Z(n650) );
  NANDN U146 ( .A(n301), .B(n259), .Z(n290) );
  NANDN U147 ( .A(n98), .B(n53), .Z(n87) );
  NANDN U148 ( .A(n3828), .B(n3786), .Z(n3817) );
  NANDN U149 ( .A(n2948), .B(n2906), .Z(n2937) );
  NANDN U150 ( .A(n2148), .B(n2106), .Z(n2137) );
  XOR U151 ( .A(n2367), .B(n2361), .Z(n2276) );
  XOR U152 ( .A(n2378), .B(n2372), .Z(n2245) );
  XOR U153 ( .A(n2355), .B(n2349), .Z(n2238) );
  XOR U154 ( .A(n2255), .B(n2250), .Z(n2231) );
  XOR U155 ( .A(n3148), .B(n3167), .Z(n3210) );
  XNOR U156 ( .A(n3142), .B(n3161), .Z(n1633) );
  XOR U157 ( .A(n4875), .B(n4870), .Z(n4799) );
  XOR U158 ( .A(n4805), .B(n4841), .Z(n4838) );
  AND U159 ( .A(n4436), .B(n4421), .Z(n4427) );
  XOR U160 ( .A(n640), .B(n1438), .Z(n422) );
  XOR U161 ( .A(n1835), .B(n1883), .Z(n1829) );
  XOR U162 ( .A(n1650), .B(n1673), .Z(n1644) );
  XOR U163 ( .A(n1455), .B(n1477), .Z(n1449) );
  XOR U164 ( .A(n1244), .B(n1266), .Z(n1238) );
  XOR U165 ( .A(n1048), .B(n1070), .Z(n1042) );
  XOR U166 ( .A(n832), .B(n870), .Z(n826) );
  XNOR U167 ( .A(n469), .B(n457), .Z(n427) );
  XOR U168 ( .A(n233), .B(n255), .Z(n227) );
  XOR U169 ( .A(n27), .B(n49), .Z(n21) );
  XNOR U170 ( .A(n12), .B(n19), .Z(n13) );
  XOR U171 ( .A(n3950), .B(n3957), .Z(n10) );
  XOR U172 ( .A(n3066), .B(n3782), .Z(n3060) );
  XOR U173 ( .A(n2880), .B(n2902), .Z(n2874) );
  XOR U174 ( .A(n2080), .B(n2102), .Z(n2074) );
  XOR U175 ( .A(n3199), .B(n3184), .Z(n178) );
  XOR U176 ( .A(n814), .B(n1392), .Z(n2390) );
  XOR U177 ( .A(n187), .B(n188), .Z(n186) );
  XOR U178 ( .A(n1036), .B(n1035), .Z(n1032) );
  XNOR U179 ( .A(n1224), .B(n1221), .Z(n1815) );
  XOR U180 ( .A(n1), .B(n2), .Z(out[9]) );
  XNOR U181 ( .A(n3), .B(n4), .Z(n2) );
  XOR U182 ( .A(key[137]), .B(n5), .Z(n1) );
  XOR U183 ( .A(n6), .B(n7), .Z(out[99]) );
  XNOR U184 ( .A(n8), .B(n9), .Z(n7) );
  XOR U185 ( .A(n10), .B(n11), .Z(n6) );
  XNOR U186 ( .A(key[227]), .B(n12), .Z(n11) );
  XNOR U187 ( .A(key[226]), .B(n13), .Z(out[98]) );
  XOR U188 ( .A(n14), .B(n15), .Z(out[97]) );
  XNOR U189 ( .A(n8), .B(n16), .Z(n15) );
  XNOR U190 ( .A(key[225]), .B(n12), .Z(n14) );
  XOR U191 ( .A(n17), .B(n18), .Z(out[96]) );
  XNOR U192 ( .A(key[224]), .B(n19), .Z(n18) );
  XOR U193 ( .A(n20), .B(n21), .Z(out[95]) );
  XOR U194 ( .A(n22), .B(n23), .Z(n20) );
  XOR U195 ( .A(key[223]), .B(n24), .Z(n23) );
  XNOR U196 ( .A(n25), .B(n26), .Z(out[94]) );
  XNOR U197 ( .A(key[222]), .B(n27), .Z(n26) );
  XOR U198 ( .A(n28), .B(n29), .Z(out[93]) );
  XNOR U199 ( .A(n30), .B(n31), .Z(n29) );
  XOR U200 ( .A(n22), .B(n32), .Z(n31) );
  XNOR U201 ( .A(n34), .B(n35), .Z(n33) );
  NANDN U202 ( .A(n36), .B(n37), .Z(n35) );
  XOR U203 ( .A(n39), .B(n40), .Z(n28) );
  XOR U204 ( .A(key[221]), .B(n41), .Z(n40) );
  ANDN U205 ( .B(n42), .A(n43), .Z(n39) );
  XNOR U206 ( .A(n44), .B(n45), .Z(out[92]) );
  XNOR U207 ( .A(key[220]), .B(n46), .Z(n45) );
  XOR U208 ( .A(n47), .B(n48), .Z(out[91]) );
  XNOR U209 ( .A(n49), .B(n25), .Z(n48) );
  XNOR U210 ( .A(n50), .B(n51), .Z(n25) );
  XNOR U211 ( .A(n52), .B(n41), .Z(n51) );
  ANDN U212 ( .B(n53), .A(n54), .Z(n41) );
  NOR U213 ( .A(n55), .B(n56), .Z(n52) );
  XNOR U214 ( .A(n57), .B(n58), .Z(n47) );
  XOR U215 ( .A(key[219]), .B(n24), .Z(n58) );
  XOR U216 ( .A(key[218]), .B(n44), .Z(out[90]) );
  XNOR U217 ( .A(n59), .B(n60), .Z(n44) );
  XNOR U218 ( .A(n61), .B(n62), .Z(out[8]) );
  XNOR U219 ( .A(key[136]), .B(n63), .Z(n62) );
  XOR U220 ( .A(n64), .B(n21), .Z(out[89]) );
  XNOR U221 ( .A(n50), .B(n65), .Z(n49) );
  XNOR U222 ( .A(n66), .B(n67), .Z(n65) );
  NANDN U223 ( .A(n68), .B(n37), .Z(n67) );
  XNOR U224 ( .A(n32), .B(n69), .Z(n50) );
  XNOR U225 ( .A(n70), .B(n71), .Z(n69) );
  NANDN U226 ( .A(n72), .B(n73), .Z(n71) );
  XOR U227 ( .A(n60), .B(n57), .Z(n27) );
  XNOR U228 ( .A(n32), .B(n74), .Z(n57) );
  XNOR U229 ( .A(n66), .B(n75), .Z(n74) );
  NANDN U230 ( .A(n76), .B(n77), .Z(n75) );
  OR U231 ( .A(n78), .B(n79), .Z(n66) );
  XOR U232 ( .A(n80), .B(n70), .Z(n32) );
  NANDN U233 ( .A(n81), .B(n82), .Z(n70) );
  ANDN U234 ( .B(n83), .A(n84), .Z(n80) );
  XNOR U235 ( .A(key[217]), .B(n59), .Z(n64) );
  IV U236 ( .A(n24), .Z(n59) );
  XOR U237 ( .A(n85), .B(n86), .Z(n24) );
  XNOR U238 ( .A(n87), .B(n88), .Z(n86) );
  NAND U239 ( .A(n42), .B(n89), .Z(n88) );
  XNOR U240 ( .A(n30), .B(n90), .Z(out[88]) );
  XOR U241 ( .A(key[216]), .B(n60), .Z(n90) );
  XNOR U242 ( .A(n85), .B(n91), .Z(n60) );
  XOR U243 ( .A(n92), .B(n34), .Z(n91) );
  OR U244 ( .A(n93), .B(n78), .Z(n34) );
  XNOR U245 ( .A(n37), .B(n77), .Z(n78) );
  ANDN U246 ( .B(n94), .A(n95), .Z(n92) );
  IV U247 ( .A(n46), .Z(n30) );
  XOR U248 ( .A(n38), .B(n96), .Z(n46) );
  XOR U249 ( .A(n97), .B(n87), .Z(n96) );
  XNOR U250 ( .A(n56), .B(n42), .Z(n53) );
  NOR U251 ( .A(n99), .B(n56), .Z(n97) );
  XNOR U252 ( .A(n85), .B(n100), .Z(n38) );
  XNOR U253 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U254 ( .A(n72), .B(n103), .Z(n102) );
  XOR U255 ( .A(n104), .B(n101), .Z(n85) );
  OR U256 ( .A(n81), .B(n105), .Z(n101) );
  XOR U257 ( .A(n106), .B(n72), .Z(n81) );
  XNOR U258 ( .A(n77), .B(n42), .Z(n72) );
  XOR U259 ( .A(n107), .B(n108), .Z(n42) );
  NANDN U260 ( .A(n109), .B(n110), .Z(n108) );
  IV U261 ( .A(n95), .Z(n77) );
  XNOR U262 ( .A(n111), .B(n112), .Z(n95) );
  NANDN U263 ( .A(n109), .B(n113), .Z(n112) );
  ANDN U264 ( .B(n106), .A(n114), .Z(n104) );
  IV U265 ( .A(n84), .Z(n106) );
  XOR U266 ( .A(n56), .B(n37), .Z(n84) );
  XNOR U267 ( .A(n115), .B(n111), .Z(n37) );
  NANDN U268 ( .A(n116), .B(n117), .Z(n111) );
  XOR U269 ( .A(n113), .B(n118), .Z(n117) );
  ANDN U270 ( .B(n118), .A(n119), .Z(n115) );
  XOR U271 ( .A(n120), .B(n107), .Z(n56) );
  NANDN U272 ( .A(n116), .B(n121), .Z(n107) );
  XOR U273 ( .A(n122), .B(n110), .Z(n121) );
  XNOR U274 ( .A(n123), .B(n124), .Z(n109) );
  XOR U275 ( .A(n125), .B(n126), .Z(n124) );
  XNOR U276 ( .A(n127), .B(n128), .Z(n123) );
  XNOR U277 ( .A(n129), .B(n130), .Z(n128) );
  ANDN U278 ( .B(n122), .A(n126), .Z(n129) );
  ANDN U279 ( .B(n122), .A(n119), .Z(n120) );
  XNOR U280 ( .A(n125), .B(n131), .Z(n119) );
  XOR U281 ( .A(n132), .B(n130), .Z(n131) );
  NAND U282 ( .A(n133), .B(n134), .Z(n130) );
  XNOR U283 ( .A(n127), .B(n110), .Z(n134) );
  IV U284 ( .A(n122), .Z(n127) );
  XNOR U285 ( .A(n113), .B(n126), .Z(n133) );
  IV U286 ( .A(n118), .Z(n126) );
  XOR U287 ( .A(n135), .B(n136), .Z(n118) );
  XNOR U288 ( .A(n137), .B(n138), .Z(n136) );
  XNOR U289 ( .A(n139), .B(n140), .Z(n135) );
  NOR U290 ( .A(n55), .B(n99), .Z(n139) );
  AND U291 ( .A(n110), .B(n113), .Z(n132) );
  XNOR U292 ( .A(n110), .B(n113), .Z(n125) );
  XNOR U293 ( .A(n141), .B(n142), .Z(n113) );
  XNOR U294 ( .A(n143), .B(n138), .Z(n142) );
  XOR U295 ( .A(n144), .B(n145), .Z(n141) );
  XNOR U296 ( .A(n146), .B(n140), .Z(n145) );
  OR U297 ( .A(n54), .B(n98), .Z(n140) );
  XOR U298 ( .A(n99), .B(n89), .Z(n98) );
  XNOR U299 ( .A(n55), .B(n43), .Z(n54) );
  ANDN U300 ( .B(n89), .A(n43), .Z(n146) );
  XNOR U301 ( .A(n147), .B(n148), .Z(n110) );
  XNOR U302 ( .A(n138), .B(n149), .Z(n148) );
  XOR U303 ( .A(n68), .B(n144), .Z(n149) );
  XNOR U304 ( .A(n99), .B(n150), .Z(n138) );
  XNOR U305 ( .A(n151), .B(n152), .Z(n147) );
  XNOR U306 ( .A(n153), .B(n154), .Z(n152) );
  ANDN U307 ( .B(n94), .A(n76), .Z(n153) );
  XNOR U308 ( .A(n155), .B(n156), .Z(n122) );
  XNOR U309 ( .A(n143), .B(n157), .Z(n156) );
  XNOR U310 ( .A(n76), .B(n137), .Z(n157) );
  XOR U311 ( .A(n144), .B(n158), .Z(n137) );
  XNOR U312 ( .A(n159), .B(n160), .Z(n158) );
  NAND U313 ( .A(n103), .B(n73), .Z(n160) );
  XNOR U314 ( .A(n161), .B(n159), .Z(n144) );
  NANDN U315 ( .A(n105), .B(n82), .Z(n159) );
  XOR U316 ( .A(n83), .B(n73), .Z(n82) );
  XNOR U317 ( .A(n162), .B(n43), .Z(n73) );
  XOR U318 ( .A(n114), .B(n103), .Z(n105) );
  XOR U319 ( .A(n94), .B(n89), .Z(n103) );
  ANDN U320 ( .B(n83), .A(n114), .Z(n161) );
  XOR U321 ( .A(n151), .B(n99), .Z(n114) );
  XOR U322 ( .A(n163), .B(n164), .Z(n99) );
  XOR U323 ( .A(n165), .B(n166), .Z(n164) );
  XOR U324 ( .A(n167), .B(n150), .Z(n83) );
  XNOR U325 ( .A(n168), .B(n169), .Z(n43) );
  XNOR U326 ( .A(n170), .B(n166), .Z(n169) );
  XNOR U327 ( .A(n166), .B(n168), .Z(n89) );
  XNOR U328 ( .A(n94), .B(n171), .Z(n155) );
  XNOR U329 ( .A(n172), .B(n154), .Z(n171) );
  OR U330 ( .A(n79), .B(n93), .Z(n154) );
  XNOR U331 ( .A(n151), .B(n94), .Z(n93) );
  XOR U332 ( .A(n68), .B(n162), .Z(n79) );
  IV U333 ( .A(n76), .Z(n162) );
  XOR U334 ( .A(n150), .B(n173), .Z(n76) );
  XNOR U335 ( .A(n170), .B(n163), .Z(n173) );
  XOR U336 ( .A(key[218]), .B(\w0[1][90] ), .Z(n163) );
  XOR U337 ( .A(n174), .B(n175), .Z(\w0[1][90] ) );
  XOR U338 ( .A(n176), .B(n177), .Z(n175) );
  XOR U339 ( .A(n178), .B(n179), .Z(n174) );
  IV U340 ( .A(n55), .Z(n150) );
  XNOR U341 ( .A(n168), .B(n180), .Z(n55) );
  XNOR U342 ( .A(n166), .B(n181), .Z(n180) );
  ANDN U343 ( .B(n167), .A(n36), .Z(n172) );
  IV U344 ( .A(n68), .Z(n167) );
  XNOR U345 ( .A(n168), .B(n182), .Z(n68) );
  XNOR U346 ( .A(n166), .B(n183), .Z(n182) );
  XOR U347 ( .A(n36), .B(n184), .Z(n166) );
  XOR U348 ( .A(key[222]), .B(\w0[1][94] ), .Z(n184) );
  XNOR U349 ( .A(n185), .B(n186), .Z(\w0[1][94] ) );
  IV U350 ( .A(n151), .Z(n36) );
  XOR U351 ( .A(key[221]), .B(\w0[1][93] ), .Z(n168) );
  XOR U352 ( .A(n189), .B(n190), .Z(\w0[1][93] ) );
  XOR U353 ( .A(n191), .B(n192), .Z(n190) );
  XOR U354 ( .A(n193), .B(n194), .Z(n189) );
  XOR U355 ( .A(n195), .B(n196), .Z(n94) );
  XNOR U356 ( .A(n183), .B(n181), .Z(n196) );
  XOR U357 ( .A(key[223]), .B(\w0[1][95] ), .Z(n181) );
  XNOR U358 ( .A(n197), .B(n198), .Z(\w0[1][95] ) );
  XOR U359 ( .A(n199), .B(n200), .Z(n198) );
  XOR U360 ( .A(key[220]), .B(\w0[1][92] ), .Z(n183) );
  XOR U361 ( .A(n201), .B(n202), .Z(\w0[1][92] ) );
  XOR U362 ( .A(n203), .B(n204), .Z(n202) );
  XOR U363 ( .A(n205), .B(n206), .Z(n201) );
  XNOR U364 ( .A(n151), .B(n165), .Z(n195) );
  XOR U365 ( .A(n170), .B(n207), .Z(n165) );
  XOR U366 ( .A(key[219]), .B(\w0[1][91] ), .Z(n207) );
  XOR U367 ( .A(n208), .B(n209), .Z(\w0[1][91] ) );
  XOR U368 ( .A(n210), .B(n211), .Z(n209) );
  XOR U369 ( .A(n212), .B(n213), .Z(n208) );
  XOR U370 ( .A(key[217]), .B(\w0[1][89] ), .Z(n170) );
  XOR U371 ( .A(n214), .B(n215), .Z(\w0[1][89] ) );
  XOR U372 ( .A(n216), .B(n217), .Z(n215) );
  XOR U373 ( .A(n218), .B(n219), .Z(n214) );
  XOR U374 ( .A(key[216]), .B(\w0[1][88] ), .Z(n151) );
  XOR U375 ( .A(n220), .B(n221), .Z(\w0[1][88] ) );
  XOR U376 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U377 ( .A(n224), .B(n225), .Z(n220) );
  XOR U378 ( .A(n226), .B(n227), .Z(out[87]) );
  XOR U379 ( .A(n228), .B(n229), .Z(n226) );
  XNOR U380 ( .A(key[215]), .B(n230), .Z(n229) );
  XNOR U381 ( .A(n231), .B(n232), .Z(out[86]) );
  XNOR U382 ( .A(key[214]), .B(n233), .Z(n232) );
  XOR U383 ( .A(n234), .B(n235), .Z(out[85]) );
  XNOR U384 ( .A(n236), .B(n237), .Z(n235) );
  XOR U385 ( .A(n228), .B(n238), .Z(n237) );
  XNOR U386 ( .A(n240), .B(n241), .Z(n239) );
  NANDN U387 ( .A(n242), .B(n243), .Z(n241) );
  XOR U388 ( .A(n245), .B(n246), .Z(n234) );
  XOR U389 ( .A(key[213]), .B(n247), .Z(n246) );
  ANDN U390 ( .B(n248), .A(n249), .Z(n245) );
  XNOR U391 ( .A(n250), .B(n251), .Z(out[84]) );
  XNOR U392 ( .A(key[212]), .B(n252), .Z(n251) );
  XOR U393 ( .A(n253), .B(n254), .Z(out[83]) );
  XNOR U394 ( .A(n255), .B(n231), .Z(n254) );
  XNOR U395 ( .A(n256), .B(n257), .Z(n231) );
  XNOR U396 ( .A(n258), .B(n247), .Z(n257) );
  ANDN U397 ( .B(n259), .A(n260), .Z(n247) );
  NOR U398 ( .A(n261), .B(n262), .Z(n258) );
  XNOR U399 ( .A(n263), .B(n264), .Z(n253) );
  XOR U400 ( .A(key[211]), .B(n265), .Z(n264) );
  XOR U401 ( .A(key[210]), .B(n250), .Z(out[82]) );
  XNOR U402 ( .A(n230), .B(n266), .Z(n250) );
  IV U403 ( .A(n265), .Z(n230) );
  XOR U404 ( .A(n267), .B(n227), .Z(out[81]) );
  XNOR U405 ( .A(n256), .B(n268), .Z(n255) );
  XNOR U406 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U407 ( .A(n271), .B(n243), .Z(n270) );
  XNOR U408 ( .A(n238), .B(n272), .Z(n256) );
  XNOR U409 ( .A(n273), .B(n274), .Z(n272) );
  NANDN U410 ( .A(n275), .B(n276), .Z(n274) );
  XOR U411 ( .A(n266), .B(n263), .Z(n233) );
  XNOR U412 ( .A(n238), .B(n277), .Z(n263) );
  XNOR U413 ( .A(n269), .B(n278), .Z(n277) );
  NANDN U414 ( .A(n279), .B(n280), .Z(n278) );
  OR U415 ( .A(n281), .B(n282), .Z(n269) );
  XOR U416 ( .A(n283), .B(n273), .Z(n238) );
  NANDN U417 ( .A(n284), .B(n285), .Z(n273) );
  ANDN U418 ( .B(n286), .A(n287), .Z(n283) );
  XOR U419 ( .A(key[209]), .B(n265), .Z(n267) );
  XOR U420 ( .A(n288), .B(n289), .Z(n265) );
  XNOR U421 ( .A(n290), .B(n291), .Z(n289) );
  NAND U422 ( .A(n248), .B(n292), .Z(n291) );
  XNOR U423 ( .A(n236), .B(n293), .Z(out[80]) );
  XOR U424 ( .A(key[208]), .B(n266), .Z(n293) );
  XNOR U425 ( .A(n288), .B(n294), .Z(n266) );
  XOR U426 ( .A(n295), .B(n240), .Z(n294) );
  OR U427 ( .A(n296), .B(n281), .Z(n240) );
  XNOR U428 ( .A(n243), .B(n280), .Z(n281) );
  ANDN U429 ( .B(n297), .A(n298), .Z(n295) );
  IV U430 ( .A(n252), .Z(n236) );
  XOR U431 ( .A(n244), .B(n299), .Z(n252) );
  XOR U432 ( .A(n300), .B(n290), .Z(n299) );
  XNOR U433 ( .A(n262), .B(n248), .Z(n259) );
  NOR U434 ( .A(n302), .B(n262), .Z(n300) );
  XNOR U435 ( .A(n288), .B(n303), .Z(n244) );
  XNOR U436 ( .A(n304), .B(n305), .Z(n303) );
  NANDN U437 ( .A(n275), .B(n306), .Z(n305) );
  XOR U438 ( .A(n307), .B(n304), .Z(n288) );
  OR U439 ( .A(n284), .B(n308), .Z(n304) );
  XOR U440 ( .A(n309), .B(n275), .Z(n284) );
  XNOR U441 ( .A(n280), .B(n248), .Z(n275) );
  XOR U442 ( .A(n310), .B(n311), .Z(n248) );
  NANDN U443 ( .A(n312), .B(n313), .Z(n311) );
  IV U444 ( .A(n298), .Z(n280) );
  XNOR U445 ( .A(n314), .B(n315), .Z(n298) );
  NANDN U446 ( .A(n312), .B(n316), .Z(n315) );
  ANDN U447 ( .B(n309), .A(n317), .Z(n307) );
  IV U448 ( .A(n287), .Z(n309) );
  XOR U449 ( .A(n262), .B(n243), .Z(n287) );
  XNOR U450 ( .A(n318), .B(n314), .Z(n243) );
  NANDN U451 ( .A(n319), .B(n320), .Z(n314) );
  XOR U452 ( .A(n316), .B(n321), .Z(n320) );
  ANDN U453 ( .B(n321), .A(n322), .Z(n318) );
  XOR U454 ( .A(n323), .B(n310), .Z(n262) );
  NANDN U455 ( .A(n319), .B(n324), .Z(n310) );
  XOR U456 ( .A(n325), .B(n313), .Z(n324) );
  XNOR U457 ( .A(n326), .B(n327), .Z(n312) );
  XOR U458 ( .A(n328), .B(n329), .Z(n327) );
  XNOR U459 ( .A(n330), .B(n331), .Z(n326) );
  XNOR U460 ( .A(n332), .B(n333), .Z(n331) );
  ANDN U461 ( .B(n325), .A(n329), .Z(n332) );
  ANDN U462 ( .B(n325), .A(n322), .Z(n323) );
  XNOR U463 ( .A(n328), .B(n334), .Z(n322) );
  XOR U464 ( .A(n335), .B(n333), .Z(n334) );
  NAND U465 ( .A(n336), .B(n337), .Z(n333) );
  XNOR U466 ( .A(n330), .B(n313), .Z(n337) );
  IV U467 ( .A(n325), .Z(n330) );
  XNOR U468 ( .A(n316), .B(n329), .Z(n336) );
  IV U469 ( .A(n321), .Z(n329) );
  XOR U470 ( .A(n338), .B(n339), .Z(n321) );
  XNOR U471 ( .A(n340), .B(n341), .Z(n339) );
  XNOR U472 ( .A(n342), .B(n343), .Z(n338) );
  NOR U473 ( .A(n261), .B(n302), .Z(n342) );
  AND U474 ( .A(n313), .B(n316), .Z(n335) );
  XNOR U475 ( .A(n313), .B(n316), .Z(n328) );
  XNOR U476 ( .A(n344), .B(n345), .Z(n316) );
  XNOR U477 ( .A(n346), .B(n341), .Z(n345) );
  XOR U478 ( .A(n347), .B(n348), .Z(n344) );
  XNOR U479 ( .A(n349), .B(n343), .Z(n348) );
  OR U480 ( .A(n260), .B(n301), .Z(n343) );
  XOR U481 ( .A(n302), .B(n292), .Z(n301) );
  XNOR U482 ( .A(n261), .B(n249), .Z(n260) );
  ANDN U483 ( .B(n292), .A(n249), .Z(n349) );
  XNOR U484 ( .A(n350), .B(n351), .Z(n313) );
  XNOR U485 ( .A(n341), .B(n352), .Z(n351) );
  XOR U486 ( .A(n271), .B(n347), .Z(n352) );
  XNOR U487 ( .A(n302), .B(n353), .Z(n341) );
  XNOR U488 ( .A(n354), .B(n355), .Z(n350) );
  XNOR U489 ( .A(n356), .B(n357), .Z(n355) );
  ANDN U490 ( .B(n297), .A(n279), .Z(n356) );
  XNOR U491 ( .A(n358), .B(n359), .Z(n325) );
  XNOR U492 ( .A(n346), .B(n360), .Z(n359) );
  XNOR U493 ( .A(n279), .B(n340), .Z(n360) );
  XOR U494 ( .A(n347), .B(n361), .Z(n340) );
  XNOR U495 ( .A(n362), .B(n363), .Z(n361) );
  NAND U496 ( .A(n306), .B(n276), .Z(n363) );
  XNOR U497 ( .A(n364), .B(n362), .Z(n347) );
  NANDN U498 ( .A(n308), .B(n285), .Z(n362) );
  XOR U499 ( .A(n286), .B(n276), .Z(n285) );
  XNOR U500 ( .A(n365), .B(n249), .Z(n276) );
  XOR U501 ( .A(n317), .B(n306), .Z(n308) );
  XOR U502 ( .A(n297), .B(n292), .Z(n306) );
  ANDN U503 ( .B(n286), .A(n317), .Z(n364) );
  XOR U504 ( .A(n354), .B(n302), .Z(n317) );
  XOR U505 ( .A(n366), .B(n367), .Z(n302) );
  XOR U506 ( .A(n368), .B(n369), .Z(n367) );
  XOR U507 ( .A(n370), .B(n353), .Z(n286) );
  XNOR U508 ( .A(n371), .B(n372), .Z(n249) );
  XNOR U509 ( .A(n373), .B(n369), .Z(n372) );
  XNOR U510 ( .A(n369), .B(n371), .Z(n292) );
  XNOR U511 ( .A(n297), .B(n374), .Z(n358) );
  XNOR U512 ( .A(n375), .B(n357), .Z(n374) );
  OR U513 ( .A(n282), .B(n296), .Z(n357) );
  XNOR U514 ( .A(n354), .B(n297), .Z(n296) );
  XOR U515 ( .A(n271), .B(n365), .Z(n282) );
  IV U516 ( .A(n279), .Z(n365) );
  XOR U517 ( .A(n353), .B(n376), .Z(n279) );
  XNOR U518 ( .A(n373), .B(n366), .Z(n376) );
  XOR U519 ( .A(key[178]), .B(\w0[1][50] ), .Z(n366) );
  XNOR U520 ( .A(n377), .B(n378), .Z(\w0[1][50] ) );
  XNOR U521 ( .A(n379), .B(n380), .Z(n378) );
  IV U522 ( .A(n261), .Z(n353) );
  XNOR U523 ( .A(n371), .B(n381), .Z(n261) );
  XNOR U524 ( .A(n369), .B(n382), .Z(n381) );
  ANDN U525 ( .B(n370), .A(n242), .Z(n375) );
  IV U526 ( .A(n271), .Z(n370) );
  XNOR U527 ( .A(n371), .B(n383), .Z(n271) );
  XNOR U528 ( .A(n369), .B(n384), .Z(n383) );
  XOR U529 ( .A(n242), .B(n385), .Z(n369) );
  XOR U530 ( .A(key[182]), .B(\w0[1][54] ), .Z(n385) );
  XNOR U531 ( .A(n386), .B(n387), .Z(\w0[1][54] ) );
  XNOR U532 ( .A(n388), .B(n389), .Z(n387) );
  IV U533 ( .A(n354), .Z(n242) );
  XOR U534 ( .A(key[181]), .B(\w0[1][53] ), .Z(n371) );
  XNOR U535 ( .A(n390), .B(n391), .Z(\w0[1][53] ) );
  XOR U536 ( .A(n392), .B(n393), .Z(n391) );
  XOR U537 ( .A(n394), .B(n395), .Z(n297) );
  XNOR U538 ( .A(n384), .B(n382), .Z(n395) );
  XOR U539 ( .A(key[183]), .B(\w0[1][55] ), .Z(n382) );
  XNOR U540 ( .A(n396), .B(n397), .Z(\w0[1][55] ) );
  XOR U541 ( .A(n398), .B(n399), .Z(n397) );
  XOR U542 ( .A(key[180]), .B(\w0[1][52] ), .Z(n384) );
  XOR U543 ( .A(n400), .B(n401), .Z(\w0[1][52] ) );
  XNOR U544 ( .A(n402), .B(n403), .Z(n401) );
  XOR U545 ( .A(n404), .B(n405), .Z(n400) );
  XNOR U546 ( .A(n354), .B(n368), .Z(n394) );
  XOR U547 ( .A(n373), .B(n406), .Z(n368) );
  XOR U548 ( .A(key[179]), .B(\w0[1][51] ), .Z(n406) );
  XOR U549 ( .A(n407), .B(n408), .Z(\w0[1][51] ) );
  XNOR U550 ( .A(n409), .B(n410), .Z(n408) );
  XOR U551 ( .A(n411), .B(n412), .Z(n407) );
  XOR U552 ( .A(key[177]), .B(\w0[1][49] ), .Z(n373) );
  XNOR U553 ( .A(n413), .B(n414), .Z(\w0[1][49] ) );
  XOR U554 ( .A(n415), .B(n416), .Z(n414) );
  XOR U555 ( .A(key[176]), .B(\w0[1][48] ), .Z(n354) );
  XOR U556 ( .A(n417), .B(n418), .Z(\w0[1][48] ) );
  XNOR U557 ( .A(n419), .B(n420), .Z(n418) );
  XOR U558 ( .A(n421), .B(n422), .Z(out[7]) );
  XOR U559 ( .A(n423), .B(n424), .Z(n421) );
  XOR U560 ( .A(key[135]), .B(n425), .Z(n424) );
  XOR U561 ( .A(n426), .B(n427), .Z(out[79]) );
  XOR U562 ( .A(n428), .B(n429), .Z(n426) );
  XNOR U563 ( .A(key[207]), .B(n430), .Z(n429) );
  XOR U564 ( .A(n431), .B(n432), .Z(out[78]) );
  XNOR U565 ( .A(n433), .B(n434), .Z(n432) );
  XNOR U566 ( .A(key[206]), .B(n435), .Z(n431) );
  XOR U567 ( .A(n436), .B(n437), .Z(out[77]) );
  XNOR U568 ( .A(n438), .B(n439), .Z(n437) );
  XOR U569 ( .A(n428), .B(n440), .Z(n439) );
  XNOR U570 ( .A(n442), .B(n443), .Z(n441) );
  OR U571 ( .A(n444), .B(n445), .Z(n443) );
  XOR U572 ( .A(n447), .B(n448), .Z(n436) );
  XOR U573 ( .A(key[205]), .B(n449), .Z(n448) );
  ANDN U574 ( .B(n450), .A(n451), .Z(n447) );
  XNOR U575 ( .A(n452), .B(n453), .Z(out[76]) );
  XNOR U576 ( .A(key[204]), .B(n454), .Z(n453) );
  XOR U577 ( .A(n455), .B(n456), .Z(out[75]) );
  XNOR U578 ( .A(n457), .B(n434), .Z(n456) );
  XNOR U579 ( .A(n458), .B(n459), .Z(n434) );
  XNOR U580 ( .A(n460), .B(n449), .Z(n459) );
  NOR U581 ( .A(n461), .B(n462), .Z(n449) );
  NOR U582 ( .A(n463), .B(n464), .Z(n460) );
  XOR U583 ( .A(n465), .B(n466), .Z(n455) );
  XOR U584 ( .A(key[203]), .B(n467), .Z(n466) );
  XOR U585 ( .A(key[202]), .B(n452), .Z(out[74]) );
  XNOR U586 ( .A(n430), .B(n435), .Z(n452) );
  XOR U587 ( .A(n468), .B(n427), .Z(out[73]) );
  XNOR U588 ( .A(n458), .B(n470), .Z(n457) );
  XOR U589 ( .A(n471), .B(n472), .Z(n470) );
  ANDN U590 ( .B(n473), .A(n444), .Z(n471) );
  XNOR U591 ( .A(n440), .B(n474), .Z(n458) );
  XNOR U592 ( .A(n475), .B(n476), .Z(n474) );
  NAND U593 ( .A(n477), .B(n478), .Z(n476) );
  XOR U594 ( .A(n435), .B(n465), .Z(n469) );
  IV U595 ( .A(n433), .Z(n465) );
  XNOR U596 ( .A(n440), .B(n479), .Z(n433) );
  XNOR U597 ( .A(n472), .B(n480), .Z(n479) );
  NANDN U598 ( .A(n481), .B(n482), .Z(n480) );
  OR U599 ( .A(n483), .B(n484), .Z(n472) );
  XOR U600 ( .A(n485), .B(n475), .Z(n440) );
  NANDN U601 ( .A(n486), .B(n487), .Z(n475) );
  AND U602 ( .A(n488), .B(n489), .Z(n485) );
  XNOR U603 ( .A(key[201]), .B(n430), .Z(n468) );
  IV U604 ( .A(n467), .Z(n430) );
  XOR U605 ( .A(n490), .B(n491), .Z(n467) );
  XNOR U606 ( .A(n492), .B(n493), .Z(n491) );
  NANDN U607 ( .A(n451), .B(n494), .Z(n493) );
  XNOR U608 ( .A(n438), .B(n495), .Z(out[72]) );
  XOR U609 ( .A(key[200]), .B(n435), .Z(n495) );
  XNOR U610 ( .A(n490), .B(n496), .Z(n435) );
  XOR U611 ( .A(n497), .B(n442), .Z(n496) );
  OR U612 ( .A(n498), .B(n483), .Z(n442) );
  XNOR U613 ( .A(n444), .B(n481), .Z(n483) );
  NOR U614 ( .A(n499), .B(n481), .Z(n497) );
  IV U615 ( .A(n454), .Z(n438) );
  XOR U616 ( .A(n446), .B(n500), .Z(n454) );
  XNOR U617 ( .A(n492), .B(n501), .Z(n500) );
  OR U618 ( .A(n464), .B(n502), .Z(n501) );
  OR U619 ( .A(n503), .B(n461), .Z(n492) );
  XOR U620 ( .A(n464), .B(n504), .Z(n461) );
  XNOR U621 ( .A(n490), .B(n505), .Z(n446) );
  XNOR U622 ( .A(n506), .B(n507), .Z(n505) );
  NAND U623 ( .A(n478), .B(n508), .Z(n507) );
  XOR U624 ( .A(n509), .B(n506), .Z(n490) );
  OR U625 ( .A(n486), .B(n510), .Z(n506) );
  XNOR U626 ( .A(n488), .B(n478), .Z(n486) );
  XOR U627 ( .A(n481), .B(n451), .Z(n478) );
  IV U628 ( .A(n504), .Z(n451) );
  XOR U629 ( .A(n511), .B(n512), .Z(n504) );
  NANDN U630 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U631 ( .A(n515), .B(n516), .Z(n481) );
  OR U632 ( .A(n513), .B(n517), .Z(n516) );
  ANDN U633 ( .B(n488), .A(n518), .Z(n509) );
  XOR U634 ( .A(n444), .B(n464), .Z(n488) );
  XNOR U635 ( .A(n511), .B(n519), .Z(n464) );
  NANDN U636 ( .A(n520), .B(n521), .Z(n519) );
  NANDN U637 ( .A(n522), .B(n523), .Z(n511) );
  OR U638 ( .A(n525), .B(n522), .Z(n515) );
  XOR U639 ( .A(n526), .B(n513), .Z(n522) );
  XNOR U640 ( .A(n527), .B(n528), .Z(n513) );
  XOR U641 ( .A(n529), .B(n521), .Z(n528) );
  XNOR U642 ( .A(n530), .B(n531), .Z(n527) );
  XNOR U643 ( .A(n532), .B(n533), .Z(n531) );
  ANDN U644 ( .B(n521), .A(n534), .Z(n532) );
  IV U645 ( .A(n535), .Z(n521) );
  ANDN U646 ( .B(n526), .A(n534), .Z(n524) );
  IV U647 ( .A(n520), .Z(n526) );
  XNOR U648 ( .A(n529), .B(n536), .Z(n520) );
  XNOR U649 ( .A(n533), .B(n537), .Z(n536) );
  NANDN U650 ( .A(n517), .B(n514), .Z(n537) );
  NANDN U651 ( .A(n525), .B(n523), .Z(n533) );
  XNOR U652 ( .A(n514), .B(n535), .Z(n523) );
  XOR U653 ( .A(n538), .B(n539), .Z(n535) );
  XOR U654 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U655 ( .A(n482), .B(n542), .Z(n541) );
  XNOR U656 ( .A(n543), .B(n544), .Z(n538) );
  XNOR U657 ( .A(n545), .B(n546), .Z(n544) );
  ANDN U658 ( .B(n473), .A(n445), .Z(n545) );
  XNOR U659 ( .A(n534), .B(n517), .Z(n525) );
  IV U660 ( .A(n530), .Z(n534) );
  XOR U661 ( .A(n547), .B(n548), .Z(n530) );
  XNOR U662 ( .A(n549), .B(n542), .Z(n548) );
  XOR U663 ( .A(n550), .B(n551), .Z(n542) );
  XNOR U664 ( .A(n552), .B(n553), .Z(n551) );
  NAND U665 ( .A(n508), .B(n477), .Z(n553) );
  XNOR U666 ( .A(n554), .B(n555), .Z(n547) );
  ANDN U667 ( .B(n556), .A(n502), .Z(n554) );
  XOR U668 ( .A(n517), .B(n514), .Z(n529) );
  XNOR U669 ( .A(n557), .B(n558), .Z(n514) );
  XNOR U670 ( .A(n550), .B(n559), .Z(n558) );
  XNOR U671 ( .A(n549), .B(n473), .Z(n559) );
  XNOR U672 ( .A(n560), .B(n561), .Z(n557) );
  XNOR U673 ( .A(n562), .B(n546), .Z(n561) );
  OR U674 ( .A(n484), .B(n498), .Z(n546) );
  XNOR U675 ( .A(n560), .B(n543), .Z(n498) );
  XNOR U676 ( .A(n473), .B(n482), .Z(n484) );
  ANDN U677 ( .B(n482), .A(n499), .Z(n562) );
  XOR U678 ( .A(n563), .B(n564), .Z(n517) );
  XOR U679 ( .A(n550), .B(n540), .Z(n564) );
  XNOR U680 ( .A(n494), .B(n450), .Z(n540) );
  XOR U681 ( .A(n565), .B(n552), .Z(n550) );
  NANDN U682 ( .A(n510), .B(n487), .Z(n552) );
  XOR U683 ( .A(n489), .B(n477), .Z(n487) );
  XOR U684 ( .A(n450), .B(n482), .Z(n477) );
  XNOR U685 ( .A(n556), .B(n566), .Z(n482) );
  XNOR U686 ( .A(n567), .B(n568), .Z(n566) );
  XOR U687 ( .A(n518), .B(n508), .Z(n510) );
  XNOR U688 ( .A(n499), .B(n494), .Z(n508) );
  IV U689 ( .A(n543), .Z(n499) );
  XOR U690 ( .A(n569), .B(n570), .Z(n543) );
  XNOR U691 ( .A(n571), .B(n572), .Z(n570) );
  XNOR U692 ( .A(n560), .B(n573), .Z(n569) );
  ANDN U693 ( .B(n489), .A(n518), .Z(n565) );
  XNOR U694 ( .A(n560), .B(n574), .Z(n518) );
  XOR U695 ( .A(n556), .B(n473), .Z(n489) );
  XNOR U696 ( .A(n575), .B(n576), .Z(n473) );
  XOR U697 ( .A(n577), .B(n572), .Z(n576) );
  XNOR U698 ( .A(key[140]), .B(\w0[1][12] ), .Z(n572) );
  XNOR U699 ( .A(n578), .B(n579), .Z(\w0[1][12] ) );
  XOR U700 ( .A(n580), .B(n581), .Z(n579) );
  XOR U701 ( .A(n549), .B(n582), .Z(n563) );
  XNOR U702 ( .A(n583), .B(n555), .Z(n582) );
  OR U703 ( .A(n462), .B(n503), .Z(n555) );
  XNOR U704 ( .A(n574), .B(n494), .Z(n503) );
  XNOR U705 ( .A(n556), .B(n450), .Z(n462) );
  IV U706 ( .A(n463), .Z(n556) );
  AND U707 ( .A(n450), .B(n494), .Z(n583) );
  XOR U708 ( .A(n577), .B(n575), .Z(n494) );
  XNOR U709 ( .A(n575), .B(n584), .Z(n450) );
  XOR U710 ( .A(n567), .B(n585), .Z(n584) );
  XNOR U711 ( .A(n502), .B(n463), .Z(n549) );
  XOR U712 ( .A(n575), .B(n586), .Z(n463) );
  XOR U713 ( .A(n577), .B(n571), .Z(n586) );
  XNOR U714 ( .A(key[143]), .B(\w0[1][15] ), .Z(n571) );
  XNOR U715 ( .A(n587), .B(n588), .Z(\w0[1][15] ) );
  XOR U716 ( .A(n589), .B(n590), .Z(n588) );
  XNOR U717 ( .A(key[141]), .B(\w0[1][13] ), .Z(n575) );
  XOR U718 ( .A(n591), .B(n592), .Z(\w0[1][13] ) );
  XOR U719 ( .A(n593), .B(n594), .Z(n592) );
  XNOR U720 ( .A(n595), .B(n596), .Z(n591) );
  IV U721 ( .A(n574), .Z(n502) );
  XNOR U722 ( .A(n568), .B(n597), .Z(n574) );
  XNOR U723 ( .A(n573), .B(n585), .Z(n597) );
  IV U724 ( .A(n577), .Z(n585) );
  XOR U725 ( .A(n445), .B(n598), .Z(n577) );
  XOR U726 ( .A(key[142]), .B(\w0[1][14] ), .Z(n598) );
  XNOR U727 ( .A(n599), .B(n600), .Z(\w0[1][14] ) );
  XNOR U728 ( .A(n601), .B(n602), .Z(n600) );
  IV U729 ( .A(n560), .Z(n445) );
  XOR U730 ( .A(key[136]), .B(\w0[1][8] ), .Z(n560) );
  XOR U731 ( .A(n603), .B(n604), .Z(\w0[1][8] ) );
  XNOR U732 ( .A(n605), .B(n606), .Z(n604) );
  XNOR U733 ( .A(n607), .B(n608), .Z(n603) );
  XOR U734 ( .A(n567), .B(n609), .Z(n573) );
  XOR U735 ( .A(key[139]), .B(\w0[1][11] ), .Z(n609) );
  XOR U736 ( .A(n610), .B(n611), .Z(\w0[1][11] ) );
  XNOR U737 ( .A(n612), .B(n613), .Z(n611) );
  XNOR U738 ( .A(n614), .B(n615), .Z(n610) );
  XOR U739 ( .A(key[137]), .B(\w0[1][9] ), .Z(n567) );
  XOR U740 ( .A(n616), .B(n617), .Z(\w0[1][9] ) );
  XOR U741 ( .A(n618), .B(n619), .Z(n617) );
  XNOR U742 ( .A(n620), .B(n621), .Z(n616) );
  XOR U743 ( .A(key[138]), .B(\w0[1][10] ), .Z(n568) );
  XOR U744 ( .A(n622), .B(n623), .Z(\w0[1][10] ) );
  XNOR U745 ( .A(n624), .B(n625), .Z(n623) );
  XNOR U746 ( .A(n626), .B(n627), .Z(n622) );
  XOR U747 ( .A(n628), .B(n629), .Z(out[71]) );
  XNOR U748 ( .A(n630), .B(n631), .Z(n628) );
  XNOR U749 ( .A(key[199]), .B(n632), .Z(n631) );
  XOR U750 ( .A(n633), .B(n634), .Z(out[70]) );
  XNOR U751 ( .A(n635), .B(n636), .Z(n634) );
  XNOR U752 ( .A(key[198]), .B(n637), .Z(n633) );
  XNOR U753 ( .A(n638), .B(n639), .Z(out[6]) );
  XNOR U754 ( .A(key[134]), .B(n640), .Z(n639) );
  XOR U755 ( .A(n641), .B(n642), .Z(out[69]) );
  XNOR U756 ( .A(n643), .B(n644), .Z(n642) );
  XNOR U757 ( .A(n632), .B(n645), .Z(n644) );
  XNOR U758 ( .A(n646), .B(n647), .Z(n632) );
  XNOR U759 ( .A(n648), .B(n649), .Z(n647) );
  OR U760 ( .A(n650), .B(n651), .Z(n649) );
  XNOR U761 ( .A(n652), .B(n653), .Z(n641) );
  XOR U762 ( .A(key[197]), .B(n654), .Z(n653) );
  ANDN U763 ( .B(n655), .A(n656), .Z(n654) );
  XNOR U764 ( .A(n657), .B(n658), .Z(out[68]) );
  XNOR U765 ( .A(key[196]), .B(n659), .Z(n658) );
  XOR U766 ( .A(n660), .B(n661), .Z(out[67]) );
  XNOR U767 ( .A(n662), .B(n636), .Z(n661) );
  XNOR U768 ( .A(n663), .B(n664), .Z(n636) );
  XNOR U769 ( .A(n652), .B(n665), .Z(n664) );
  OR U770 ( .A(n666), .B(n667), .Z(n665) );
  NANDN U771 ( .A(n668), .B(n669), .Z(n652) );
  XNOR U772 ( .A(n670), .B(n671), .Z(n660) );
  XNOR U773 ( .A(key[195]), .B(n635), .Z(n671) );
  XOR U774 ( .A(key[194]), .B(n657), .Z(out[66]) );
  XNOR U775 ( .A(n637), .B(n662), .Z(n657) );
  XOR U776 ( .A(n672), .B(n629), .Z(out[65]) );
  XNOR U777 ( .A(n670), .B(n662), .Z(n629) );
  XNOR U778 ( .A(n673), .B(n674), .Z(n662) );
  XNOR U779 ( .A(n675), .B(n676), .Z(n674) );
  NAND U780 ( .A(n677), .B(n655), .Z(n676) );
  XNOR U781 ( .A(n663), .B(n678), .Z(n670) );
  XNOR U782 ( .A(n679), .B(n680), .Z(n678) );
  NANDN U783 ( .A(n650), .B(n681), .Z(n680) );
  XNOR U784 ( .A(n645), .B(n682), .Z(n663) );
  XNOR U785 ( .A(n683), .B(n684), .Z(n682) );
  NANDN U786 ( .A(n685), .B(n686), .Z(n684) );
  XNOR U787 ( .A(key[193]), .B(n630), .Z(n672) );
  XOR U788 ( .A(n687), .B(n635), .Z(n630) );
  XNOR U789 ( .A(n645), .B(n688), .Z(n635) );
  XOR U790 ( .A(n689), .B(n679), .Z(n688) );
  OR U791 ( .A(n690), .B(n691), .Z(n679) );
  AND U792 ( .A(n692), .B(n693), .Z(n689) );
  XOR U793 ( .A(n694), .B(n683), .Z(n645) );
  NANDN U794 ( .A(n695), .B(n696), .Z(n683) );
  AND U795 ( .A(n697), .B(n698), .Z(n694) );
  XNOR U796 ( .A(n643), .B(n699), .Z(out[64]) );
  XNOR U797 ( .A(key[192]), .B(n687), .Z(n699) );
  IV U798 ( .A(n637), .Z(n687) );
  XNOR U799 ( .A(n673), .B(n700), .Z(n637) );
  XOR U800 ( .A(n701), .B(n648), .Z(n700) );
  OR U801 ( .A(n702), .B(n690), .Z(n648) );
  XOR U802 ( .A(n650), .B(n693), .Z(n690) );
  ANDN U803 ( .B(n693), .A(n703), .Z(n701) );
  IV U804 ( .A(n659), .Z(n643) );
  XOR U805 ( .A(n646), .B(n704), .Z(n659) );
  XOR U806 ( .A(n705), .B(n675), .Z(n704) );
  NANDN U807 ( .A(n706), .B(n669), .Z(n675) );
  XNOR U808 ( .A(n666), .B(n655), .Z(n669) );
  NOR U809 ( .A(n707), .B(n666), .Z(n705) );
  XNOR U810 ( .A(n673), .B(n708), .Z(n646) );
  XNOR U811 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U812 ( .A(n685), .B(n711), .Z(n710) );
  XOR U813 ( .A(n712), .B(n709), .Z(n673) );
  OR U814 ( .A(n695), .B(n713), .Z(n709) );
  XOR U815 ( .A(n697), .B(n685), .Z(n695) );
  XNOR U816 ( .A(n693), .B(n655), .Z(n685) );
  XOR U817 ( .A(n714), .B(n715), .Z(n655) );
  NANDN U818 ( .A(n716), .B(n717), .Z(n715) );
  XOR U819 ( .A(n718), .B(n719), .Z(n693) );
  OR U820 ( .A(n716), .B(n720), .Z(n719) );
  ANDN U821 ( .B(n697), .A(n721), .Z(n712) );
  XOR U822 ( .A(n650), .B(n666), .Z(n697) );
  XOR U823 ( .A(n722), .B(n714), .Z(n666) );
  NANDN U824 ( .A(n723), .B(n724), .Z(n714) );
  ANDN U825 ( .B(n725), .A(n726), .Z(n722) );
  NANDN U826 ( .A(n723), .B(n728), .Z(n718) );
  XOR U827 ( .A(n729), .B(n716), .Z(n723) );
  XNOR U828 ( .A(n730), .B(n731), .Z(n716) );
  XOR U829 ( .A(n732), .B(n725), .Z(n731) );
  XNOR U830 ( .A(n733), .B(n734), .Z(n730) );
  XNOR U831 ( .A(n735), .B(n736), .Z(n734) );
  ANDN U832 ( .B(n725), .A(n737), .Z(n735) );
  IV U833 ( .A(n738), .Z(n725) );
  ANDN U834 ( .B(n729), .A(n737), .Z(n727) );
  IV U835 ( .A(n733), .Z(n737) );
  IV U836 ( .A(n726), .Z(n729) );
  XNOR U837 ( .A(n732), .B(n739), .Z(n726) );
  XOR U838 ( .A(n740), .B(n736), .Z(n739) );
  NAND U839 ( .A(n728), .B(n724), .Z(n736) );
  XNOR U840 ( .A(n717), .B(n738), .Z(n724) );
  XOR U841 ( .A(n741), .B(n742), .Z(n738) );
  XOR U842 ( .A(n743), .B(n744), .Z(n742) );
  XNOR U843 ( .A(n692), .B(n745), .Z(n744) );
  XNOR U844 ( .A(n746), .B(n747), .Z(n741) );
  XNOR U845 ( .A(n748), .B(n749), .Z(n747) );
  ANDN U846 ( .B(n681), .A(n651), .Z(n748) );
  XNOR U847 ( .A(n733), .B(n720), .Z(n728) );
  XOR U848 ( .A(n750), .B(n751), .Z(n733) );
  XNOR U849 ( .A(n752), .B(n745), .Z(n751) );
  XOR U850 ( .A(n753), .B(n754), .Z(n745) );
  XNOR U851 ( .A(n755), .B(n756), .Z(n754) );
  NAND U852 ( .A(n711), .B(n686), .Z(n756) );
  XNOR U853 ( .A(n757), .B(n758), .Z(n750) );
  ANDN U854 ( .B(n759), .A(n707), .Z(n757) );
  ANDN U855 ( .B(n717), .A(n720), .Z(n740) );
  XOR U856 ( .A(n720), .B(n717), .Z(n732) );
  XNOR U857 ( .A(n760), .B(n761), .Z(n717) );
  XNOR U858 ( .A(n753), .B(n762), .Z(n761) );
  XNOR U859 ( .A(n752), .B(n681), .Z(n762) );
  XNOR U860 ( .A(n763), .B(n764), .Z(n760) );
  XNOR U861 ( .A(n765), .B(n749), .Z(n764) );
  OR U862 ( .A(n691), .B(n702), .Z(n749) );
  XNOR U863 ( .A(n763), .B(n746), .Z(n702) );
  XNOR U864 ( .A(n681), .B(n692), .Z(n691) );
  ANDN U865 ( .B(n692), .A(n703), .Z(n765) );
  XOR U866 ( .A(n766), .B(n767), .Z(n720) );
  XOR U867 ( .A(n753), .B(n743), .Z(n767) );
  XOR U868 ( .A(n677), .B(n656), .Z(n743) );
  XOR U869 ( .A(n768), .B(n755), .Z(n753) );
  NANDN U870 ( .A(n713), .B(n696), .Z(n755) );
  XOR U871 ( .A(n698), .B(n686), .Z(n696) );
  XNOR U872 ( .A(n759), .B(n769), .Z(n692) );
  XOR U873 ( .A(n770), .B(n771), .Z(n769) );
  XOR U874 ( .A(n721), .B(n711), .Z(n713) );
  XNOR U875 ( .A(n703), .B(n677), .Z(n711) );
  IV U876 ( .A(n746), .Z(n703) );
  XOR U877 ( .A(n772), .B(n773), .Z(n746) );
  XNOR U878 ( .A(n774), .B(n775), .Z(n773) );
  XNOR U879 ( .A(n763), .B(n776), .Z(n772) );
  ANDN U880 ( .B(n698), .A(n721), .Z(n768) );
  XNOR U881 ( .A(n763), .B(n777), .Z(n721) );
  XOR U882 ( .A(n759), .B(n681), .Z(n698) );
  XNOR U883 ( .A(n778), .B(n779), .Z(n681) );
  XNOR U884 ( .A(n780), .B(n775), .Z(n779) );
  XOR U885 ( .A(key[228]), .B(\w0[1][100] ), .Z(n775) );
  XOR U886 ( .A(n781), .B(n782), .Z(\w0[1][100] ) );
  XNOR U887 ( .A(n783), .B(n784), .Z(n782) );
  XOR U888 ( .A(n785), .B(n786), .Z(n781) );
  IV U889 ( .A(n667), .Z(n759) );
  XOR U890 ( .A(n752), .B(n787), .Z(n766) );
  XNOR U891 ( .A(n788), .B(n758), .Z(n787) );
  OR U892 ( .A(n668), .B(n706), .Z(n758) );
  XNOR U893 ( .A(n777), .B(n677), .Z(n706) );
  XNOR U894 ( .A(n667), .B(n656), .Z(n668) );
  ANDN U895 ( .B(n677), .A(n656), .Z(n788) );
  XOR U896 ( .A(n778), .B(n789), .Z(n656) );
  XNOR U897 ( .A(n790), .B(n780), .Z(n789) );
  XOR U898 ( .A(n780), .B(n778), .Z(n677) );
  XNOR U899 ( .A(n707), .B(n667), .Z(n752) );
  XOR U900 ( .A(n778), .B(n791), .Z(n667) );
  XNOR U901 ( .A(n780), .B(n774), .Z(n791) );
  XOR U902 ( .A(key[231]), .B(\w0[1][103] ), .Z(n774) );
  XNOR U903 ( .A(n792), .B(n793), .Z(\w0[1][103] ) );
  XOR U904 ( .A(n794), .B(n795), .Z(n793) );
  XNOR U905 ( .A(key[229]), .B(\w0[1][101] ), .Z(n778) );
  XNOR U906 ( .A(n796), .B(n797), .Z(\w0[1][101] ) );
  XOR U907 ( .A(n798), .B(n799), .Z(n797) );
  IV U908 ( .A(n777), .Z(n707) );
  XOR U909 ( .A(n770), .B(n776), .Z(n800) );
  XNOR U910 ( .A(n771), .B(n801), .Z(n776) );
  XOR U911 ( .A(key[227]), .B(\w0[1][99] ), .Z(n801) );
  XOR U912 ( .A(n802), .B(n803), .Z(\w0[1][99] ) );
  XOR U913 ( .A(n804), .B(n805), .Z(n803) );
  XOR U914 ( .A(n806), .B(n807), .Z(n802) );
  IV U915 ( .A(n790), .Z(n771) );
  XOR U916 ( .A(key[225]), .B(\w0[1][97] ), .Z(n790) );
  XNOR U917 ( .A(n808), .B(n809), .Z(\w0[1][97] ) );
  XNOR U918 ( .A(n810), .B(n811), .Z(n809) );
  XOR U919 ( .A(key[226]), .B(\w0[1][98] ), .Z(n770) );
  XNOR U920 ( .A(n812), .B(n813), .Z(\w0[1][98] ) );
  XNOR U921 ( .A(n814), .B(n815), .Z(n813) );
  XOR U922 ( .A(n651), .B(n816), .Z(n780) );
  XOR U923 ( .A(key[230]), .B(\w0[1][102] ), .Z(n816) );
  XNOR U924 ( .A(n817), .B(n818), .Z(\w0[1][102] ) );
  XNOR U925 ( .A(n819), .B(n820), .Z(n818) );
  IV U926 ( .A(n763), .Z(n651) );
  XOR U927 ( .A(key[224]), .B(\w0[1][96] ), .Z(n763) );
  XNOR U928 ( .A(n821), .B(n822), .Z(\w0[1][96] ) );
  XOR U929 ( .A(n823), .B(n824), .Z(n822) );
  XOR U930 ( .A(n825), .B(n826), .Z(out[63]) );
  XOR U931 ( .A(n827), .B(n828), .Z(n825) );
  XOR U932 ( .A(key[191]), .B(n829), .Z(n828) );
  XNOR U933 ( .A(n830), .B(n831), .Z(out[62]) );
  XNOR U934 ( .A(key[190]), .B(n832), .Z(n831) );
  XOR U935 ( .A(n833), .B(n834), .Z(out[61]) );
  XNOR U936 ( .A(n835), .B(n836), .Z(n834) );
  XOR U937 ( .A(n827), .B(n837), .Z(n836) );
  XNOR U938 ( .A(n839), .B(n840), .Z(n838) );
  NANDN U939 ( .A(n841), .B(n842), .Z(n840) );
  XOR U940 ( .A(n844), .B(n845), .Z(n833) );
  XOR U941 ( .A(key[189]), .B(n846), .Z(n845) );
  ANDN U942 ( .B(n847), .A(n848), .Z(n844) );
  XNOR U943 ( .A(n849), .B(n850), .Z(out[60]) );
  XNOR U944 ( .A(key[188]), .B(n851), .Z(n850) );
  XOR U945 ( .A(n852), .B(n853), .Z(out[5]) );
  XNOR U946 ( .A(n854), .B(n855), .Z(n853) );
  XOR U947 ( .A(n423), .B(n856), .Z(n855) );
  XNOR U948 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U949 ( .A(n860), .B(n861), .Z(n859) );
  XOR U950 ( .A(n863), .B(n864), .Z(n852) );
  XOR U951 ( .A(key[133]), .B(n865), .Z(n864) );
  ANDN U952 ( .B(n866), .A(n867), .Z(n863) );
  XOR U953 ( .A(n868), .B(n869), .Z(out[59]) );
  XNOR U954 ( .A(n870), .B(n830), .Z(n869) );
  XNOR U955 ( .A(n871), .B(n872), .Z(n830) );
  XNOR U956 ( .A(n873), .B(n846), .Z(n872) );
  ANDN U957 ( .B(n874), .A(n875), .Z(n846) );
  NOR U958 ( .A(n876), .B(n877), .Z(n873) );
  XNOR U959 ( .A(n878), .B(n879), .Z(n868) );
  XOR U960 ( .A(key[187]), .B(n829), .Z(n879) );
  XOR U961 ( .A(key[186]), .B(n849), .Z(out[58]) );
  XNOR U962 ( .A(n880), .B(n881), .Z(n849) );
  XOR U963 ( .A(n882), .B(n826), .Z(out[57]) );
  XNOR U964 ( .A(n871), .B(n883), .Z(n870) );
  XNOR U965 ( .A(n884), .B(n885), .Z(n883) );
  NANDN U966 ( .A(n886), .B(n842), .Z(n885) );
  XNOR U967 ( .A(n837), .B(n887), .Z(n871) );
  XNOR U968 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U969 ( .A(n890), .B(n891), .Z(n889) );
  XOR U970 ( .A(n881), .B(n878), .Z(n832) );
  XNOR U971 ( .A(n837), .B(n892), .Z(n878) );
  XNOR U972 ( .A(n884), .B(n893), .Z(n892) );
  NANDN U973 ( .A(n894), .B(n895), .Z(n893) );
  OR U974 ( .A(n896), .B(n897), .Z(n884) );
  XOR U975 ( .A(n898), .B(n888), .Z(n837) );
  NANDN U976 ( .A(n899), .B(n900), .Z(n888) );
  ANDN U977 ( .B(n901), .A(n902), .Z(n898) );
  XNOR U978 ( .A(key[185]), .B(n880), .Z(n882) );
  IV U979 ( .A(n829), .Z(n880) );
  XOR U980 ( .A(n903), .B(n904), .Z(n829) );
  XNOR U981 ( .A(n905), .B(n906), .Z(n904) );
  NAND U982 ( .A(n847), .B(n907), .Z(n906) );
  XNOR U983 ( .A(n835), .B(n908), .Z(out[56]) );
  XOR U984 ( .A(key[184]), .B(n881), .Z(n908) );
  XNOR U985 ( .A(n903), .B(n909), .Z(n881) );
  XOR U986 ( .A(n910), .B(n839), .Z(n909) );
  OR U987 ( .A(n911), .B(n896), .Z(n839) );
  XNOR U988 ( .A(n842), .B(n895), .Z(n896) );
  ANDN U989 ( .B(n912), .A(n913), .Z(n910) );
  IV U990 ( .A(n851), .Z(n835) );
  XOR U991 ( .A(n843), .B(n914), .Z(n851) );
  XOR U992 ( .A(n915), .B(n905), .Z(n914) );
  XNOR U993 ( .A(n877), .B(n847), .Z(n874) );
  NOR U994 ( .A(n917), .B(n877), .Z(n915) );
  XNOR U995 ( .A(n903), .B(n918), .Z(n843) );
  XNOR U996 ( .A(n919), .B(n920), .Z(n918) );
  NANDN U997 ( .A(n890), .B(n921), .Z(n920) );
  XOR U998 ( .A(n922), .B(n919), .Z(n903) );
  OR U999 ( .A(n899), .B(n923), .Z(n919) );
  XOR U1000 ( .A(n924), .B(n890), .Z(n899) );
  XNOR U1001 ( .A(n895), .B(n847), .Z(n890) );
  XOR U1002 ( .A(n925), .B(n926), .Z(n847) );
  NANDN U1003 ( .A(n927), .B(n928), .Z(n926) );
  IV U1004 ( .A(n913), .Z(n895) );
  XNOR U1005 ( .A(n929), .B(n930), .Z(n913) );
  NANDN U1006 ( .A(n927), .B(n931), .Z(n930) );
  ANDN U1007 ( .B(n924), .A(n932), .Z(n922) );
  IV U1008 ( .A(n902), .Z(n924) );
  XOR U1009 ( .A(n877), .B(n842), .Z(n902) );
  XNOR U1010 ( .A(n933), .B(n929), .Z(n842) );
  NANDN U1011 ( .A(n934), .B(n935), .Z(n929) );
  XOR U1012 ( .A(n931), .B(n936), .Z(n935) );
  ANDN U1013 ( .B(n936), .A(n937), .Z(n933) );
  XOR U1014 ( .A(n938), .B(n925), .Z(n877) );
  NANDN U1015 ( .A(n934), .B(n939), .Z(n925) );
  XOR U1016 ( .A(n940), .B(n928), .Z(n939) );
  XNOR U1017 ( .A(n941), .B(n942), .Z(n927) );
  XOR U1018 ( .A(n943), .B(n944), .Z(n942) );
  XNOR U1019 ( .A(n945), .B(n946), .Z(n941) );
  XNOR U1020 ( .A(n947), .B(n948), .Z(n946) );
  ANDN U1021 ( .B(n940), .A(n944), .Z(n947) );
  ANDN U1022 ( .B(n940), .A(n937), .Z(n938) );
  XNOR U1023 ( .A(n943), .B(n949), .Z(n937) );
  XOR U1024 ( .A(n950), .B(n948), .Z(n949) );
  NAND U1025 ( .A(n951), .B(n952), .Z(n948) );
  XNOR U1026 ( .A(n945), .B(n928), .Z(n952) );
  IV U1027 ( .A(n940), .Z(n945) );
  XNOR U1028 ( .A(n931), .B(n944), .Z(n951) );
  IV U1029 ( .A(n936), .Z(n944) );
  XOR U1030 ( .A(n953), .B(n954), .Z(n936) );
  XNOR U1031 ( .A(n955), .B(n956), .Z(n954) );
  XNOR U1032 ( .A(n957), .B(n958), .Z(n953) );
  NOR U1033 ( .A(n876), .B(n917), .Z(n957) );
  AND U1034 ( .A(n928), .B(n931), .Z(n950) );
  XNOR U1035 ( .A(n928), .B(n931), .Z(n943) );
  XNOR U1036 ( .A(n959), .B(n960), .Z(n931) );
  XNOR U1037 ( .A(n961), .B(n956), .Z(n960) );
  XOR U1038 ( .A(n962), .B(n963), .Z(n959) );
  XNOR U1039 ( .A(n964), .B(n958), .Z(n963) );
  OR U1040 ( .A(n875), .B(n916), .Z(n958) );
  XOR U1041 ( .A(n917), .B(n907), .Z(n916) );
  XNOR U1042 ( .A(n876), .B(n848), .Z(n875) );
  ANDN U1043 ( .B(n907), .A(n848), .Z(n964) );
  XNOR U1044 ( .A(n965), .B(n966), .Z(n928) );
  XNOR U1045 ( .A(n956), .B(n967), .Z(n966) );
  XOR U1046 ( .A(n886), .B(n962), .Z(n967) );
  XNOR U1047 ( .A(n917), .B(n968), .Z(n956) );
  XNOR U1048 ( .A(n969), .B(n970), .Z(n965) );
  XNOR U1049 ( .A(n971), .B(n972), .Z(n970) );
  ANDN U1050 ( .B(n912), .A(n894), .Z(n971) );
  XNOR U1051 ( .A(n973), .B(n974), .Z(n940) );
  XNOR U1052 ( .A(n961), .B(n975), .Z(n974) );
  XNOR U1053 ( .A(n894), .B(n955), .Z(n975) );
  XOR U1054 ( .A(n962), .B(n976), .Z(n955) );
  XNOR U1055 ( .A(n977), .B(n978), .Z(n976) );
  NAND U1056 ( .A(n921), .B(n891), .Z(n978) );
  XNOR U1057 ( .A(n979), .B(n977), .Z(n962) );
  NANDN U1058 ( .A(n923), .B(n900), .Z(n977) );
  XOR U1059 ( .A(n901), .B(n891), .Z(n900) );
  XNOR U1060 ( .A(n980), .B(n848), .Z(n891) );
  XOR U1061 ( .A(n932), .B(n921), .Z(n923) );
  XOR U1062 ( .A(n912), .B(n907), .Z(n921) );
  ANDN U1063 ( .B(n901), .A(n932), .Z(n979) );
  XOR U1064 ( .A(n969), .B(n917), .Z(n932) );
  XOR U1065 ( .A(n981), .B(n982), .Z(n917) );
  XOR U1066 ( .A(n983), .B(n984), .Z(n982) );
  XOR U1067 ( .A(n985), .B(n968), .Z(n901) );
  XNOR U1068 ( .A(n986), .B(n987), .Z(n848) );
  XNOR U1069 ( .A(n988), .B(n984), .Z(n987) );
  XNOR U1070 ( .A(n984), .B(n986), .Z(n907) );
  XNOR U1071 ( .A(n912), .B(n989), .Z(n973) );
  XNOR U1072 ( .A(n990), .B(n972), .Z(n989) );
  OR U1073 ( .A(n897), .B(n911), .Z(n972) );
  XNOR U1074 ( .A(n969), .B(n912), .Z(n911) );
  XOR U1075 ( .A(n886), .B(n980), .Z(n897) );
  IV U1076 ( .A(n894), .Z(n980) );
  XOR U1077 ( .A(n968), .B(n991), .Z(n894) );
  XNOR U1078 ( .A(n988), .B(n981), .Z(n991) );
  XOR U1079 ( .A(key[186]), .B(\w0[1][58] ), .Z(n981) );
  XOR U1080 ( .A(n992), .B(n993), .Z(\w0[1][58] ) );
  XOR U1081 ( .A(n415), .B(n994), .Z(n993) );
  IV U1082 ( .A(n995), .Z(n415) );
  XOR U1083 ( .A(n996), .B(n997), .Z(n992) );
  IV U1084 ( .A(n876), .Z(n968) );
  XNOR U1085 ( .A(n986), .B(n998), .Z(n876) );
  XNOR U1086 ( .A(n984), .B(n999), .Z(n998) );
  ANDN U1087 ( .B(n985), .A(n841), .Z(n990) );
  IV U1088 ( .A(n886), .Z(n985) );
  XNOR U1089 ( .A(n986), .B(n1000), .Z(n886) );
  XNOR U1090 ( .A(n984), .B(n1001), .Z(n1000) );
  XOR U1091 ( .A(n841), .B(n1002), .Z(n984) );
  XOR U1092 ( .A(key[190]), .B(\w0[1][62] ), .Z(n1002) );
  XNOR U1093 ( .A(n389), .B(n1003), .Z(\w0[1][62] ) );
  XNOR U1094 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U1095 ( .A(n1006), .B(n398), .Z(n389) );
  IV U1096 ( .A(n969), .Z(n841) );
  XOR U1097 ( .A(key[189]), .B(\w0[1][61] ), .Z(n986) );
  XOR U1098 ( .A(n1007), .B(n1008), .Z(\w0[1][61] ) );
  XOR U1099 ( .A(n1009), .B(n1010), .Z(n1008) );
  XOR U1100 ( .A(n1011), .B(n1012), .Z(n1007) );
  XOR U1101 ( .A(n1013), .B(n1014), .Z(n912) );
  XNOR U1102 ( .A(n1001), .B(n999), .Z(n1014) );
  XOR U1103 ( .A(key[191]), .B(\w0[1][63] ), .Z(n999) );
  XNOR U1104 ( .A(n1015), .B(n1016), .Z(\w0[1][63] ) );
  XNOR U1105 ( .A(n1017), .B(n1018), .Z(n1016) );
  XOR U1106 ( .A(key[188]), .B(\w0[1][60] ), .Z(n1001) );
  XOR U1107 ( .A(n1019), .B(n1020), .Z(\w0[1][60] ) );
  XNOR U1108 ( .A(n1021), .B(n1022), .Z(n1020) );
  XOR U1109 ( .A(n1023), .B(n404), .Z(n1019) );
  XNOR U1110 ( .A(n398), .B(n1024), .Z(n404) );
  XNOR U1111 ( .A(n969), .B(n983), .Z(n1013) );
  XOR U1112 ( .A(n988), .B(n1025), .Z(n983) );
  XOR U1113 ( .A(key[187]), .B(\w0[1][59] ), .Z(n1025) );
  XOR U1114 ( .A(n1026), .B(n1027), .Z(\w0[1][59] ) );
  XOR U1115 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U1116 ( .A(n1030), .B(n411), .Z(n1026) );
  XOR U1117 ( .A(n398), .B(n1031), .Z(n411) );
  XOR U1118 ( .A(key[185]), .B(\w0[1][57] ), .Z(n988) );
  XOR U1119 ( .A(n1032), .B(n1033), .Z(\w0[1][57] ) );
  XOR U1120 ( .A(n1034), .B(n420), .Z(n1033) );
  XOR U1121 ( .A(key[184]), .B(\w0[1][56] ), .Z(n969) );
  XOR U1122 ( .A(n1037), .B(n1038), .Z(\w0[1][56] ) );
  XOR U1123 ( .A(n417), .B(n1039), .Z(n1038) );
  XNOR U1124 ( .A(n398), .B(n1040), .Z(n1037) );
  XOR U1125 ( .A(n1041), .B(n1042), .Z(out[55]) );
  XOR U1126 ( .A(n1043), .B(n1044), .Z(n1041) );
  XOR U1127 ( .A(key[183]), .B(n1045), .Z(n1044) );
  XNOR U1128 ( .A(n1046), .B(n1047), .Z(out[54]) );
  XNOR U1129 ( .A(key[182]), .B(n1048), .Z(n1047) );
  XOR U1130 ( .A(n1049), .B(n1050), .Z(out[53]) );
  XNOR U1131 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U1132 ( .A(n1043), .B(n1053), .Z(n1052) );
  XNOR U1133 ( .A(n1055), .B(n1056), .Z(n1054) );
  NANDN U1134 ( .A(n1057), .B(n1058), .Z(n1056) );
  XOR U1135 ( .A(n1060), .B(n1061), .Z(n1049) );
  XOR U1136 ( .A(key[181]), .B(n1062), .Z(n1061) );
  ANDN U1137 ( .B(n1063), .A(n1064), .Z(n1060) );
  XNOR U1138 ( .A(n1065), .B(n1066), .Z(out[52]) );
  XNOR U1139 ( .A(key[180]), .B(n1067), .Z(n1066) );
  XOR U1140 ( .A(n1068), .B(n1069), .Z(out[51]) );
  XNOR U1141 ( .A(n1070), .B(n1046), .Z(n1069) );
  XNOR U1142 ( .A(n1071), .B(n1072), .Z(n1046) );
  XNOR U1143 ( .A(n1073), .B(n1062), .Z(n1072) );
  ANDN U1144 ( .B(n1074), .A(n1075), .Z(n1062) );
  NOR U1145 ( .A(n1076), .B(n1077), .Z(n1073) );
  XNOR U1146 ( .A(n1078), .B(n1079), .Z(n1068) );
  XOR U1147 ( .A(key[179]), .B(n1045), .Z(n1079) );
  XOR U1148 ( .A(key[178]), .B(n1065), .Z(out[50]) );
  XNOR U1149 ( .A(n1080), .B(n1081), .Z(n1065) );
  XNOR U1150 ( .A(n1082), .B(n1083), .Z(out[4]) );
  XNOR U1151 ( .A(key[132]), .B(n1084), .Z(n1083) );
  XOR U1152 ( .A(n1085), .B(n1042), .Z(out[49]) );
  XNOR U1153 ( .A(n1071), .B(n1086), .Z(n1070) );
  XNOR U1154 ( .A(n1087), .B(n1088), .Z(n1086) );
  NANDN U1155 ( .A(n1089), .B(n1058), .Z(n1088) );
  XNOR U1156 ( .A(n1053), .B(n1090), .Z(n1071) );
  XNOR U1157 ( .A(n1091), .B(n1092), .Z(n1090) );
  NANDN U1158 ( .A(n1093), .B(n1094), .Z(n1092) );
  XOR U1159 ( .A(n1081), .B(n1078), .Z(n1048) );
  XNOR U1160 ( .A(n1053), .B(n1095), .Z(n1078) );
  XNOR U1161 ( .A(n1087), .B(n1096), .Z(n1095) );
  NANDN U1162 ( .A(n1097), .B(n1098), .Z(n1096) );
  OR U1163 ( .A(n1099), .B(n1100), .Z(n1087) );
  XOR U1164 ( .A(n1101), .B(n1091), .Z(n1053) );
  NANDN U1165 ( .A(n1102), .B(n1103), .Z(n1091) );
  ANDN U1166 ( .B(n1104), .A(n1105), .Z(n1101) );
  XNOR U1167 ( .A(key[177]), .B(n1080), .Z(n1085) );
  IV U1168 ( .A(n1045), .Z(n1080) );
  XOR U1169 ( .A(n1106), .B(n1107), .Z(n1045) );
  XNOR U1170 ( .A(n1108), .B(n1109), .Z(n1107) );
  NAND U1171 ( .A(n1063), .B(n1110), .Z(n1109) );
  XNOR U1172 ( .A(n1051), .B(n1111), .Z(out[48]) );
  XOR U1173 ( .A(key[176]), .B(n1081), .Z(n1111) );
  XNOR U1174 ( .A(n1106), .B(n1112), .Z(n1081) );
  XOR U1175 ( .A(n1113), .B(n1055), .Z(n1112) );
  OR U1176 ( .A(n1114), .B(n1099), .Z(n1055) );
  XNOR U1177 ( .A(n1058), .B(n1098), .Z(n1099) );
  ANDN U1178 ( .B(n1115), .A(n1116), .Z(n1113) );
  IV U1179 ( .A(n1067), .Z(n1051) );
  XOR U1180 ( .A(n1059), .B(n1117), .Z(n1067) );
  XOR U1181 ( .A(n1118), .B(n1108), .Z(n1117) );
  XNOR U1182 ( .A(n1077), .B(n1063), .Z(n1074) );
  NOR U1183 ( .A(n1120), .B(n1077), .Z(n1118) );
  XNOR U1184 ( .A(n1106), .B(n1121), .Z(n1059) );
  XNOR U1185 ( .A(n1122), .B(n1123), .Z(n1121) );
  NANDN U1186 ( .A(n1093), .B(n1124), .Z(n1123) );
  XOR U1187 ( .A(n1125), .B(n1122), .Z(n1106) );
  OR U1188 ( .A(n1102), .B(n1126), .Z(n1122) );
  XOR U1189 ( .A(n1127), .B(n1093), .Z(n1102) );
  XNOR U1190 ( .A(n1098), .B(n1063), .Z(n1093) );
  XOR U1191 ( .A(n1128), .B(n1129), .Z(n1063) );
  NANDN U1192 ( .A(n1130), .B(n1131), .Z(n1129) );
  IV U1193 ( .A(n1116), .Z(n1098) );
  XNOR U1194 ( .A(n1132), .B(n1133), .Z(n1116) );
  NANDN U1195 ( .A(n1130), .B(n1134), .Z(n1133) );
  ANDN U1196 ( .B(n1127), .A(n1135), .Z(n1125) );
  IV U1197 ( .A(n1105), .Z(n1127) );
  XOR U1198 ( .A(n1077), .B(n1058), .Z(n1105) );
  XNOR U1199 ( .A(n1136), .B(n1132), .Z(n1058) );
  NANDN U1200 ( .A(n1137), .B(n1138), .Z(n1132) );
  XOR U1201 ( .A(n1134), .B(n1139), .Z(n1138) );
  ANDN U1202 ( .B(n1139), .A(n1140), .Z(n1136) );
  XOR U1203 ( .A(n1141), .B(n1128), .Z(n1077) );
  NANDN U1204 ( .A(n1137), .B(n1142), .Z(n1128) );
  XOR U1205 ( .A(n1143), .B(n1131), .Z(n1142) );
  XNOR U1206 ( .A(n1144), .B(n1145), .Z(n1130) );
  XOR U1207 ( .A(n1146), .B(n1147), .Z(n1145) );
  XNOR U1208 ( .A(n1148), .B(n1149), .Z(n1144) );
  XNOR U1209 ( .A(n1150), .B(n1151), .Z(n1149) );
  ANDN U1210 ( .B(n1143), .A(n1147), .Z(n1150) );
  ANDN U1211 ( .B(n1143), .A(n1140), .Z(n1141) );
  XNOR U1212 ( .A(n1146), .B(n1152), .Z(n1140) );
  XOR U1213 ( .A(n1153), .B(n1151), .Z(n1152) );
  NAND U1214 ( .A(n1154), .B(n1155), .Z(n1151) );
  XNOR U1215 ( .A(n1148), .B(n1131), .Z(n1155) );
  IV U1216 ( .A(n1143), .Z(n1148) );
  XNOR U1217 ( .A(n1134), .B(n1147), .Z(n1154) );
  IV U1218 ( .A(n1139), .Z(n1147) );
  XOR U1219 ( .A(n1156), .B(n1157), .Z(n1139) );
  XNOR U1220 ( .A(n1158), .B(n1159), .Z(n1157) );
  XNOR U1221 ( .A(n1160), .B(n1161), .Z(n1156) );
  NOR U1222 ( .A(n1076), .B(n1120), .Z(n1160) );
  AND U1223 ( .A(n1131), .B(n1134), .Z(n1153) );
  XNOR U1224 ( .A(n1131), .B(n1134), .Z(n1146) );
  XNOR U1225 ( .A(n1162), .B(n1163), .Z(n1134) );
  XNOR U1226 ( .A(n1164), .B(n1159), .Z(n1163) );
  XOR U1227 ( .A(n1165), .B(n1166), .Z(n1162) );
  XNOR U1228 ( .A(n1167), .B(n1161), .Z(n1166) );
  OR U1229 ( .A(n1075), .B(n1119), .Z(n1161) );
  XOR U1230 ( .A(n1120), .B(n1110), .Z(n1119) );
  XNOR U1231 ( .A(n1076), .B(n1064), .Z(n1075) );
  ANDN U1232 ( .B(n1110), .A(n1064), .Z(n1167) );
  XNOR U1233 ( .A(n1168), .B(n1169), .Z(n1131) );
  XNOR U1234 ( .A(n1159), .B(n1170), .Z(n1169) );
  XOR U1235 ( .A(n1089), .B(n1165), .Z(n1170) );
  XNOR U1236 ( .A(n1120), .B(n1171), .Z(n1159) );
  XNOR U1237 ( .A(n1172), .B(n1173), .Z(n1168) );
  XNOR U1238 ( .A(n1174), .B(n1175), .Z(n1173) );
  ANDN U1239 ( .B(n1115), .A(n1097), .Z(n1174) );
  XNOR U1240 ( .A(n1176), .B(n1177), .Z(n1143) );
  XNOR U1241 ( .A(n1164), .B(n1178), .Z(n1177) );
  XNOR U1242 ( .A(n1097), .B(n1158), .Z(n1178) );
  XOR U1243 ( .A(n1165), .B(n1179), .Z(n1158) );
  XNOR U1244 ( .A(n1180), .B(n1181), .Z(n1179) );
  NAND U1245 ( .A(n1124), .B(n1094), .Z(n1181) );
  XNOR U1246 ( .A(n1182), .B(n1180), .Z(n1165) );
  NANDN U1247 ( .A(n1126), .B(n1103), .Z(n1180) );
  XOR U1248 ( .A(n1104), .B(n1094), .Z(n1103) );
  XNOR U1249 ( .A(n1183), .B(n1064), .Z(n1094) );
  XOR U1250 ( .A(n1135), .B(n1124), .Z(n1126) );
  XOR U1251 ( .A(n1115), .B(n1110), .Z(n1124) );
  ANDN U1252 ( .B(n1104), .A(n1135), .Z(n1182) );
  XOR U1253 ( .A(n1172), .B(n1120), .Z(n1135) );
  XOR U1254 ( .A(n1184), .B(n1185), .Z(n1120) );
  XOR U1255 ( .A(n1186), .B(n1187), .Z(n1185) );
  XOR U1256 ( .A(n1188), .B(n1171), .Z(n1104) );
  XNOR U1257 ( .A(n1189), .B(n1190), .Z(n1064) );
  XNOR U1258 ( .A(n1191), .B(n1187), .Z(n1190) );
  XNOR U1259 ( .A(n1187), .B(n1189), .Z(n1110) );
  XNOR U1260 ( .A(n1115), .B(n1192), .Z(n1176) );
  XNOR U1261 ( .A(n1193), .B(n1175), .Z(n1192) );
  OR U1262 ( .A(n1100), .B(n1114), .Z(n1175) );
  XNOR U1263 ( .A(n1172), .B(n1115), .Z(n1114) );
  XOR U1264 ( .A(n1089), .B(n1183), .Z(n1100) );
  IV U1265 ( .A(n1097), .Z(n1183) );
  XOR U1266 ( .A(n1171), .B(n1194), .Z(n1097) );
  XNOR U1267 ( .A(n1191), .B(n1184), .Z(n1194) );
  XOR U1268 ( .A(key[146]), .B(\w0[1][18] ), .Z(n1184) );
  XNOR U1269 ( .A(n625), .B(n1195), .Z(\w0[1][18] ) );
  XOR U1270 ( .A(n621), .B(n1196), .Z(n1195) );
  IV U1271 ( .A(n1076), .Z(n1171) );
  XNOR U1272 ( .A(n1189), .B(n1197), .Z(n1076) );
  XNOR U1273 ( .A(n1187), .B(n1198), .Z(n1197) );
  ANDN U1274 ( .B(n1188), .A(n1057), .Z(n1193) );
  IV U1275 ( .A(n1089), .Z(n1188) );
  XNOR U1276 ( .A(n1189), .B(n1199), .Z(n1089) );
  XNOR U1277 ( .A(n1187), .B(n1200), .Z(n1199) );
  XOR U1278 ( .A(n1057), .B(n1201), .Z(n1187) );
  XOR U1279 ( .A(key[150]), .B(\w0[1][22] ), .Z(n1201) );
  XNOR U1280 ( .A(n599), .B(n1202), .Z(\w0[1][22] ) );
  XNOR U1281 ( .A(n595), .B(n1203), .Z(n1202) );
  XNOR U1282 ( .A(n1204), .B(n1205), .Z(n599) );
  IV U1283 ( .A(n1172), .Z(n1057) );
  XOR U1284 ( .A(key[149]), .B(\w0[1][21] ), .Z(n1189) );
  XNOR U1285 ( .A(n594), .B(n1206), .Z(\w0[1][21] ) );
  XOR U1286 ( .A(n1207), .B(n1208), .Z(n1206) );
  XOR U1287 ( .A(n1209), .B(n1210), .Z(n594) );
  XOR U1288 ( .A(n1211), .B(n1212), .Z(n1115) );
  XNOR U1289 ( .A(n1200), .B(n1198), .Z(n1212) );
  XOR U1290 ( .A(key[151]), .B(\w0[1][23] ), .Z(n1198) );
  XNOR U1291 ( .A(n587), .B(n1213), .Z(\w0[1][23] ) );
  XOR U1292 ( .A(n1214), .B(n1205), .Z(n1213) );
  XOR U1293 ( .A(n1215), .B(n1216), .Z(n1205) );
  XNOR U1294 ( .A(n1217), .B(n1218), .Z(n587) );
  XOR U1295 ( .A(key[148]), .B(\w0[1][20] ), .Z(n1200) );
  XNOR U1296 ( .A(n578), .B(n1219), .Z(\w0[1][20] ) );
  XNOR U1297 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U1298 ( .A(n1222), .B(n1223), .Z(n578) );
  XNOR U1299 ( .A(n1224), .B(n1216), .Z(n1223) );
  XNOR U1300 ( .A(n1225), .B(n1226), .Z(n1222) );
  XNOR U1301 ( .A(n1172), .B(n1186), .Z(n1211) );
  XOR U1302 ( .A(n1191), .B(n1227), .Z(n1186) );
  XOR U1303 ( .A(key[147]), .B(\w0[1][19] ), .Z(n1227) );
  XOR U1304 ( .A(n1228), .B(n1229), .Z(\w0[1][19] ) );
  XNOR U1305 ( .A(n1230), .B(n613), .Z(n1229) );
  XOR U1306 ( .A(n1220), .B(n1216), .Z(n613) );
  XOR U1307 ( .A(n627), .B(n1231), .Z(n1228) );
  XOR U1308 ( .A(key[145]), .B(\w0[1][17] ), .Z(n1191) );
  XOR U1309 ( .A(n1232), .B(n1233), .Z(\w0[1][17] ) );
  XOR U1310 ( .A(n620), .B(n606), .Z(n1233) );
  XOR U1311 ( .A(key[144]), .B(\w0[1][16] ), .Z(n1172) );
  XNOR U1312 ( .A(n590), .B(n1234), .Z(\w0[1][16] ) );
  XOR U1313 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U1314 ( .A(n1237), .B(n1238), .Z(out[47]) );
  XOR U1315 ( .A(n1239), .B(n1240), .Z(n1237) );
  XNOR U1316 ( .A(key[175]), .B(n1241), .Z(n1240) );
  XNOR U1317 ( .A(n1242), .B(n1243), .Z(out[46]) );
  XNOR U1318 ( .A(key[174]), .B(n1244), .Z(n1243) );
  XOR U1319 ( .A(n1245), .B(n1246), .Z(out[45]) );
  XNOR U1320 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U1321 ( .A(n1239), .B(n1249), .Z(n1248) );
  XNOR U1322 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1323 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U1324 ( .A(n1256), .B(n1257), .Z(n1245) );
  XOR U1325 ( .A(key[173]), .B(n1258), .Z(n1257) );
  ANDN U1326 ( .B(n1259), .A(n1260), .Z(n1256) );
  XNOR U1327 ( .A(n1261), .B(n1262), .Z(out[44]) );
  XNOR U1328 ( .A(key[172]), .B(n1263), .Z(n1262) );
  XOR U1329 ( .A(n1264), .B(n1265), .Z(out[43]) );
  XNOR U1330 ( .A(n1266), .B(n1242), .Z(n1265) );
  XNOR U1331 ( .A(n1267), .B(n1268), .Z(n1242) );
  XNOR U1332 ( .A(n1269), .B(n1258), .Z(n1268) );
  ANDN U1333 ( .B(n1270), .A(n1271), .Z(n1258) );
  NOR U1334 ( .A(n1272), .B(n1273), .Z(n1269) );
  XNOR U1335 ( .A(n1274), .B(n1275), .Z(n1264) );
  XOR U1336 ( .A(key[171]), .B(n1276), .Z(n1275) );
  XOR U1337 ( .A(key[170]), .B(n1261), .Z(out[42]) );
  XNOR U1338 ( .A(n1241), .B(n1277), .Z(n1261) );
  IV U1339 ( .A(n1276), .Z(n1241) );
  XOR U1340 ( .A(n1278), .B(n1238), .Z(out[41]) );
  XNOR U1341 ( .A(n1267), .B(n1279), .Z(n1266) );
  XNOR U1342 ( .A(n1280), .B(n1281), .Z(n1279) );
  NANDN U1343 ( .A(n1282), .B(n1254), .Z(n1281) );
  XNOR U1344 ( .A(n1249), .B(n1283), .Z(n1267) );
  XNOR U1345 ( .A(n1284), .B(n1285), .Z(n1283) );
  NANDN U1346 ( .A(n1286), .B(n1287), .Z(n1285) );
  XOR U1347 ( .A(n1277), .B(n1274), .Z(n1244) );
  XNOR U1348 ( .A(n1249), .B(n1288), .Z(n1274) );
  XNOR U1349 ( .A(n1280), .B(n1289), .Z(n1288) );
  NANDN U1350 ( .A(n1290), .B(n1291), .Z(n1289) );
  OR U1351 ( .A(n1292), .B(n1293), .Z(n1280) );
  XOR U1352 ( .A(n1294), .B(n1284), .Z(n1249) );
  NANDN U1353 ( .A(n1295), .B(n1296), .Z(n1284) );
  ANDN U1354 ( .B(n1297), .A(n1298), .Z(n1294) );
  XOR U1355 ( .A(key[169]), .B(n1276), .Z(n1278) );
  XOR U1356 ( .A(n1299), .B(n1300), .Z(n1276) );
  XNOR U1357 ( .A(n1301), .B(n1302), .Z(n1300) );
  NAND U1358 ( .A(n1259), .B(n1303), .Z(n1302) );
  XNOR U1359 ( .A(n1247), .B(n1304), .Z(out[40]) );
  XOR U1360 ( .A(key[168]), .B(n1277), .Z(n1304) );
  XNOR U1361 ( .A(n1299), .B(n1305), .Z(n1277) );
  XOR U1362 ( .A(n1306), .B(n1251), .Z(n1305) );
  OR U1363 ( .A(n1307), .B(n1292), .Z(n1251) );
  XNOR U1364 ( .A(n1254), .B(n1291), .Z(n1292) );
  ANDN U1365 ( .B(n1308), .A(n1309), .Z(n1306) );
  IV U1366 ( .A(n1263), .Z(n1247) );
  XOR U1367 ( .A(n1255), .B(n1310), .Z(n1263) );
  XOR U1368 ( .A(n1311), .B(n1301), .Z(n1310) );
  XNOR U1369 ( .A(n1273), .B(n1259), .Z(n1270) );
  NOR U1370 ( .A(n1313), .B(n1273), .Z(n1311) );
  XNOR U1371 ( .A(n1299), .B(n1314), .Z(n1255) );
  XNOR U1372 ( .A(n1315), .B(n1316), .Z(n1314) );
  NANDN U1373 ( .A(n1286), .B(n1317), .Z(n1316) );
  XOR U1374 ( .A(n1318), .B(n1315), .Z(n1299) );
  OR U1375 ( .A(n1295), .B(n1319), .Z(n1315) );
  XOR U1376 ( .A(n1320), .B(n1286), .Z(n1295) );
  XNOR U1377 ( .A(n1291), .B(n1259), .Z(n1286) );
  XOR U1378 ( .A(n1321), .B(n1322), .Z(n1259) );
  NANDN U1379 ( .A(n1323), .B(n1324), .Z(n1322) );
  IV U1380 ( .A(n1309), .Z(n1291) );
  XNOR U1381 ( .A(n1325), .B(n1326), .Z(n1309) );
  NANDN U1382 ( .A(n1323), .B(n1327), .Z(n1326) );
  ANDN U1383 ( .B(n1320), .A(n1328), .Z(n1318) );
  IV U1384 ( .A(n1298), .Z(n1320) );
  XOR U1385 ( .A(n1273), .B(n1254), .Z(n1298) );
  XNOR U1386 ( .A(n1329), .B(n1325), .Z(n1254) );
  NANDN U1387 ( .A(n1330), .B(n1331), .Z(n1325) );
  XOR U1388 ( .A(n1327), .B(n1332), .Z(n1331) );
  ANDN U1389 ( .B(n1332), .A(n1333), .Z(n1329) );
  XOR U1390 ( .A(n1334), .B(n1321), .Z(n1273) );
  NANDN U1391 ( .A(n1330), .B(n1335), .Z(n1321) );
  XOR U1392 ( .A(n1336), .B(n1324), .Z(n1335) );
  XNOR U1393 ( .A(n1337), .B(n1338), .Z(n1323) );
  XOR U1394 ( .A(n1339), .B(n1340), .Z(n1338) );
  XNOR U1395 ( .A(n1341), .B(n1342), .Z(n1337) );
  XNOR U1396 ( .A(n1343), .B(n1344), .Z(n1342) );
  ANDN U1397 ( .B(n1336), .A(n1340), .Z(n1343) );
  ANDN U1398 ( .B(n1336), .A(n1333), .Z(n1334) );
  XNOR U1399 ( .A(n1339), .B(n1345), .Z(n1333) );
  XOR U1400 ( .A(n1346), .B(n1344), .Z(n1345) );
  NAND U1401 ( .A(n1347), .B(n1348), .Z(n1344) );
  XNOR U1402 ( .A(n1341), .B(n1324), .Z(n1348) );
  IV U1403 ( .A(n1336), .Z(n1341) );
  XNOR U1404 ( .A(n1327), .B(n1340), .Z(n1347) );
  IV U1405 ( .A(n1332), .Z(n1340) );
  XOR U1406 ( .A(n1349), .B(n1350), .Z(n1332) );
  XNOR U1407 ( .A(n1351), .B(n1352), .Z(n1350) );
  XNOR U1408 ( .A(n1353), .B(n1354), .Z(n1349) );
  NOR U1409 ( .A(n1272), .B(n1313), .Z(n1353) );
  AND U1410 ( .A(n1324), .B(n1327), .Z(n1346) );
  XNOR U1411 ( .A(n1324), .B(n1327), .Z(n1339) );
  XNOR U1412 ( .A(n1355), .B(n1356), .Z(n1327) );
  XNOR U1413 ( .A(n1357), .B(n1352), .Z(n1356) );
  XOR U1414 ( .A(n1358), .B(n1359), .Z(n1355) );
  XNOR U1415 ( .A(n1360), .B(n1354), .Z(n1359) );
  OR U1416 ( .A(n1271), .B(n1312), .Z(n1354) );
  XOR U1417 ( .A(n1313), .B(n1303), .Z(n1312) );
  XNOR U1418 ( .A(n1272), .B(n1260), .Z(n1271) );
  ANDN U1419 ( .B(n1303), .A(n1260), .Z(n1360) );
  XNOR U1420 ( .A(n1361), .B(n1362), .Z(n1324) );
  XNOR U1421 ( .A(n1352), .B(n1363), .Z(n1362) );
  XOR U1422 ( .A(n1282), .B(n1358), .Z(n1363) );
  XNOR U1423 ( .A(n1313), .B(n1364), .Z(n1352) );
  XNOR U1424 ( .A(n1365), .B(n1366), .Z(n1361) );
  XNOR U1425 ( .A(n1367), .B(n1368), .Z(n1366) );
  ANDN U1426 ( .B(n1308), .A(n1290), .Z(n1367) );
  XNOR U1427 ( .A(n1369), .B(n1370), .Z(n1336) );
  XNOR U1428 ( .A(n1357), .B(n1371), .Z(n1370) );
  XNOR U1429 ( .A(n1290), .B(n1351), .Z(n1371) );
  XOR U1430 ( .A(n1358), .B(n1372), .Z(n1351) );
  XNOR U1431 ( .A(n1373), .B(n1374), .Z(n1372) );
  NAND U1432 ( .A(n1317), .B(n1287), .Z(n1374) );
  XNOR U1433 ( .A(n1375), .B(n1373), .Z(n1358) );
  NANDN U1434 ( .A(n1319), .B(n1296), .Z(n1373) );
  XOR U1435 ( .A(n1297), .B(n1287), .Z(n1296) );
  XNOR U1436 ( .A(n1376), .B(n1260), .Z(n1287) );
  XOR U1437 ( .A(n1328), .B(n1317), .Z(n1319) );
  XOR U1438 ( .A(n1308), .B(n1303), .Z(n1317) );
  ANDN U1439 ( .B(n1297), .A(n1328), .Z(n1375) );
  XOR U1440 ( .A(n1365), .B(n1313), .Z(n1328) );
  XOR U1441 ( .A(n1377), .B(n1378), .Z(n1313) );
  XOR U1442 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U1443 ( .A(n1381), .B(n1364), .Z(n1297) );
  XNOR U1444 ( .A(n1382), .B(n1383), .Z(n1260) );
  XNOR U1445 ( .A(n1384), .B(n1380), .Z(n1383) );
  XNOR U1446 ( .A(n1380), .B(n1382), .Z(n1303) );
  XNOR U1447 ( .A(n1308), .B(n1385), .Z(n1369) );
  XNOR U1448 ( .A(n1386), .B(n1368), .Z(n1385) );
  OR U1449 ( .A(n1293), .B(n1307), .Z(n1368) );
  XNOR U1450 ( .A(n1365), .B(n1308), .Z(n1307) );
  XOR U1451 ( .A(n1282), .B(n1376), .Z(n1293) );
  IV U1452 ( .A(n1290), .Z(n1376) );
  XOR U1453 ( .A(n1364), .B(n1387), .Z(n1290) );
  XNOR U1454 ( .A(n1384), .B(n1377), .Z(n1387) );
  XOR U1455 ( .A(key[234]), .B(\w0[1][106] ), .Z(n1377) );
  XOR U1456 ( .A(n1388), .B(n1389), .Z(\w0[1][106] ) );
  XNOR U1457 ( .A(n1390), .B(n811), .Z(n1389) );
  XNOR U1458 ( .A(n1391), .B(n1392), .Z(n1388) );
  IV U1459 ( .A(n1272), .Z(n1364) );
  XNOR U1460 ( .A(n1382), .B(n1393), .Z(n1272) );
  XOR U1461 ( .A(n1380), .B(n1394), .Z(n1393) );
  ANDN U1462 ( .B(n1381), .A(n1253), .Z(n1386) );
  IV U1463 ( .A(n1282), .Z(n1381) );
  XNOR U1464 ( .A(n1382), .B(n1395), .Z(n1282) );
  XNOR U1465 ( .A(n1380), .B(n1396), .Z(n1395) );
  XOR U1466 ( .A(n1253), .B(n1397), .Z(n1380) );
  XOR U1467 ( .A(key[238]), .B(\w0[1][110] ), .Z(n1397) );
  XNOR U1468 ( .A(n817), .B(n1398), .Z(\w0[1][110] ) );
  XNOR U1469 ( .A(n1399), .B(n1400), .Z(n1398) );
  XNOR U1470 ( .A(n1401), .B(n1402), .Z(n817) );
  IV U1471 ( .A(n1365), .Z(n1253) );
  XOR U1472 ( .A(key[237]), .B(\w0[1][109] ), .Z(n1382) );
  XOR U1473 ( .A(n1403), .B(n1404), .Z(\w0[1][109] ) );
  XOR U1474 ( .A(n1405), .B(n1406), .Z(n1404) );
  XNOR U1475 ( .A(n1407), .B(n1408), .Z(n1403) );
  XOR U1476 ( .A(n1409), .B(n1410), .Z(n1308) );
  XOR U1477 ( .A(n1396), .B(n1394), .Z(n1410) );
  XNOR U1478 ( .A(key[239]), .B(\w0[1][111] ), .Z(n1394) );
  XNOR U1479 ( .A(n1411), .B(n1412), .Z(\w0[1][111] ) );
  XOR U1480 ( .A(n1413), .B(n1414), .Z(n1412) );
  XOR U1481 ( .A(key[236]), .B(\w0[1][108] ), .Z(n1396) );
  XOR U1482 ( .A(n1415), .B(n1416), .Z(\w0[1][108] ) );
  XOR U1483 ( .A(n1417), .B(n784), .Z(n1416) );
  XOR U1484 ( .A(n794), .B(n1418), .Z(n784) );
  XOR U1485 ( .A(n1419), .B(n1420), .Z(n1415) );
  XNOR U1486 ( .A(n1365), .B(n1379), .Z(n1409) );
  XOR U1487 ( .A(n1384), .B(n1421), .Z(n1379) );
  XOR U1488 ( .A(key[235]), .B(\w0[1][107] ), .Z(n1421) );
  XOR U1489 ( .A(n1422), .B(n1423), .Z(\w0[1][107] ) );
  XOR U1490 ( .A(n812), .B(n1424), .Z(n1423) );
  XOR U1491 ( .A(n806), .B(n1425), .Z(n1422) );
  XOR U1492 ( .A(n1426), .B(n794), .Z(n806) );
  IV U1493 ( .A(n1401), .Z(n794) );
  XOR U1494 ( .A(key[233]), .B(\w0[1][105] ), .Z(n1384) );
  XOR U1495 ( .A(n1427), .B(n1428), .Z(\w0[1][105] ) );
  XOR U1496 ( .A(n1429), .B(n824), .Z(n1428) );
  XOR U1497 ( .A(n1430), .B(n1431), .Z(n1427) );
  XOR U1498 ( .A(key[232]), .B(\w0[1][104] ), .Z(n1365) );
  XOR U1499 ( .A(n1432), .B(n1433), .Z(\w0[1][104] ) );
  XOR U1500 ( .A(n1434), .B(n821), .Z(n1433) );
  XNOR U1501 ( .A(n1401), .B(n1435), .Z(n1432) );
  XOR U1502 ( .A(n1436), .B(n1437), .Z(out[3]) );
  XNOR U1503 ( .A(n1438), .B(n638), .Z(n1437) );
  XNOR U1504 ( .A(n1439), .B(n1440), .Z(n638) );
  XNOR U1505 ( .A(n1441), .B(n865), .Z(n1440) );
  ANDN U1506 ( .B(n1442), .A(n1443), .Z(n865) );
  NOR U1507 ( .A(n1444), .B(n1445), .Z(n1441) );
  XNOR U1508 ( .A(n1446), .B(n1447), .Z(n1436) );
  XOR U1509 ( .A(key[131]), .B(n425), .Z(n1447) );
  XOR U1510 ( .A(n1448), .B(n1449), .Z(out[39]) );
  XOR U1511 ( .A(n1450), .B(n1451), .Z(n1448) );
  XOR U1512 ( .A(key[167]), .B(n1452), .Z(n1451) );
  XNOR U1513 ( .A(n1453), .B(n1454), .Z(out[38]) );
  XNOR U1514 ( .A(key[166]), .B(n1455), .Z(n1454) );
  XOR U1515 ( .A(n1456), .B(n1457), .Z(out[37]) );
  XNOR U1516 ( .A(n1458), .B(n1459), .Z(n1457) );
  XOR U1517 ( .A(n1450), .B(n1460), .Z(n1459) );
  XNOR U1518 ( .A(n1462), .B(n1463), .Z(n1461) );
  NANDN U1519 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U1520 ( .A(n1467), .B(n1468), .Z(n1456) );
  XOR U1521 ( .A(key[165]), .B(n1469), .Z(n1468) );
  ANDN U1522 ( .B(n1470), .A(n1471), .Z(n1467) );
  XNOR U1523 ( .A(n1472), .B(n1473), .Z(out[36]) );
  XNOR U1524 ( .A(key[164]), .B(n1474), .Z(n1473) );
  XOR U1525 ( .A(n1475), .B(n1476), .Z(out[35]) );
  XNOR U1526 ( .A(n1477), .B(n1453), .Z(n1476) );
  XNOR U1527 ( .A(n1478), .B(n1479), .Z(n1453) );
  XNOR U1528 ( .A(n1480), .B(n1469), .Z(n1479) );
  ANDN U1529 ( .B(n1481), .A(n1482), .Z(n1469) );
  NOR U1530 ( .A(n1483), .B(n1484), .Z(n1480) );
  XNOR U1531 ( .A(n1485), .B(n1486), .Z(n1475) );
  XOR U1532 ( .A(key[163]), .B(n1452), .Z(n1486) );
  XOR U1533 ( .A(key[162]), .B(n1472), .Z(out[34]) );
  XNOR U1534 ( .A(n1487), .B(n1488), .Z(n1472) );
  XOR U1535 ( .A(n1489), .B(n1449), .Z(out[33]) );
  XNOR U1536 ( .A(n1478), .B(n1490), .Z(n1477) );
  XNOR U1537 ( .A(n1491), .B(n1492), .Z(n1490) );
  NANDN U1538 ( .A(n1493), .B(n1465), .Z(n1492) );
  XNOR U1539 ( .A(n1460), .B(n1494), .Z(n1478) );
  XNOR U1540 ( .A(n1495), .B(n1496), .Z(n1494) );
  NANDN U1541 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR U1542 ( .A(n1488), .B(n1485), .Z(n1455) );
  XNOR U1543 ( .A(n1460), .B(n1499), .Z(n1485) );
  XNOR U1544 ( .A(n1491), .B(n1500), .Z(n1499) );
  NANDN U1545 ( .A(n1501), .B(n1502), .Z(n1500) );
  OR U1546 ( .A(n1503), .B(n1504), .Z(n1491) );
  XOR U1547 ( .A(n1505), .B(n1495), .Z(n1460) );
  NANDN U1548 ( .A(n1506), .B(n1507), .Z(n1495) );
  ANDN U1549 ( .B(n1508), .A(n1509), .Z(n1505) );
  XNOR U1550 ( .A(key[161]), .B(n1487), .Z(n1489) );
  IV U1551 ( .A(n1452), .Z(n1487) );
  XOR U1552 ( .A(n1510), .B(n1511), .Z(n1452) );
  XNOR U1553 ( .A(n1512), .B(n1513), .Z(n1511) );
  NANDN U1554 ( .A(n1514), .B(n1470), .Z(n1513) );
  XNOR U1555 ( .A(n1458), .B(n1515), .Z(out[32]) );
  XOR U1556 ( .A(key[160]), .B(n1488), .Z(n1515) );
  XNOR U1557 ( .A(n1510), .B(n1516), .Z(n1488) );
  XOR U1558 ( .A(n1517), .B(n1462), .Z(n1516) );
  OR U1559 ( .A(n1518), .B(n1503), .Z(n1462) );
  XNOR U1560 ( .A(n1465), .B(n1502), .Z(n1503) );
  ANDN U1561 ( .B(n1519), .A(n1520), .Z(n1517) );
  IV U1562 ( .A(n1474), .Z(n1458) );
  XOR U1563 ( .A(n1466), .B(n1521), .Z(n1474) );
  XOR U1564 ( .A(n1522), .B(n1512), .Z(n1521) );
  XNOR U1565 ( .A(n1484), .B(n1470), .Z(n1481) );
  NOR U1566 ( .A(n1524), .B(n1484), .Z(n1522) );
  XNOR U1567 ( .A(n1510), .B(n1525), .Z(n1466) );
  XNOR U1568 ( .A(n1526), .B(n1527), .Z(n1525) );
  NANDN U1569 ( .A(n1497), .B(n1528), .Z(n1527) );
  XOR U1570 ( .A(n1529), .B(n1526), .Z(n1510) );
  OR U1571 ( .A(n1506), .B(n1530), .Z(n1526) );
  XOR U1572 ( .A(n1531), .B(n1497), .Z(n1506) );
  XNOR U1573 ( .A(n1502), .B(n1470), .Z(n1497) );
  XOR U1574 ( .A(n1532), .B(n1533), .Z(n1470) );
  NANDN U1575 ( .A(n1534), .B(n1535), .Z(n1533) );
  IV U1576 ( .A(n1520), .Z(n1502) );
  XNOR U1577 ( .A(n1536), .B(n1537), .Z(n1520) );
  NANDN U1578 ( .A(n1534), .B(n1538), .Z(n1537) );
  ANDN U1579 ( .B(n1531), .A(n1539), .Z(n1529) );
  IV U1580 ( .A(n1509), .Z(n1531) );
  XOR U1581 ( .A(n1484), .B(n1465), .Z(n1509) );
  XNOR U1582 ( .A(n1540), .B(n1536), .Z(n1465) );
  NANDN U1583 ( .A(n1541), .B(n1542), .Z(n1536) );
  XOR U1584 ( .A(n1538), .B(n1543), .Z(n1542) );
  ANDN U1585 ( .B(n1543), .A(n1544), .Z(n1540) );
  XOR U1586 ( .A(n1545), .B(n1532), .Z(n1484) );
  NANDN U1587 ( .A(n1541), .B(n1546), .Z(n1532) );
  XOR U1588 ( .A(n1547), .B(n1535), .Z(n1546) );
  XNOR U1589 ( .A(n1548), .B(n1549), .Z(n1534) );
  XOR U1590 ( .A(n1550), .B(n1551), .Z(n1549) );
  XNOR U1591 ( .A(n1552), .B(n1553), .Z(n1548) );
  XNOR U1592 ( .A(n1554), .B(n1555), .Z(n1553) );
  ANDN U1593 ( .B(n1547), .A(n1551), .Z(n1554) );
  ANDN U1594 ( .B(n1547), .A(n1544), .Z(n1545) );
  XNOR U1595 ( .A(n1550), .B(n1556), .Z(n1544) );
  XOR U1596 ( .A(n1557), .B(n1555), .Z(n1556) );
  NAND U1597 ( .A(n1558), .B(n1559), .Z(n1555) );
  XNOR U1598 ( .A(n1552), .B(n1535), .Z(n1559) );
  IV U1599 ( .A(n1547), .Z(n1552) );
  XNOR U1600 ( .A(n1538), .B(n1551), .Z(n1558) );
  IV U1601 ( .A(n1543), .Z(n1551) );
  XOR U1602 ( .A(n1560), .B(n1561), .Z(n1543) );
  XNOR U1603 ( .A(n1562), .B(n1563), .Z(n1561) );
  XNOR U1604 ( .A(n1564), .B(n1565), .Z(n1560) );
  NOR U1605 ( .A(n1483), .B(n1524), .Z(n1564) );
  AND U1606 ( .A(n1535), .B(n1538), .Z(n1557) );
  XNOR U1607 ( .A(n1535), .B(n1538), .Z(n1550) );
  XNOR U1608 ( .A(n1566), .B(n1567), .Z(n1538) );
  XNOR U1609 ( .A(n1568), .B(n1563), .Z(n1567) );
  XOR U1610 ( .A(n1569), .B(n1570), .Z(n1566) );
  XNOR U1611 ( .A(n1571), .B(n1565), .Z(n1570) );
  OR U1612 ( .A(n1482), .B(n1523), .Z(n1565) );
  XNOR U1613 ( .A(n1524), .B(n1514), .Z(n1523) );
  XNOR U1614 ( .A(n1483), .B(n1471), .Z(n1482) );
  ANDN U1615 ( .B(n1572), .A(n1514), .Z(n1571) );
  XNOR U1616 ( .A(n1573), .B(n1574), .Z(n1535) );
  XNOR U1617 ( .A(n1563), .B(n1575), .Z(n1574) );
  XOR U1618 ( .A(n1493), .B(n1569), .Z(n1575) );
  XNOR U1619 ( .A(n1524), .B(n1576), .Z(n1563) );
  XNOR U1620 ( .A(n1577), .B(n1578), .Z(n1573) );
  XNOR U1621 ( .A(n1579), .B(n1580), .Z(n1578) );
  ANDN U1622 ( .B(n1519), .A(n1501), .Z(n1579) );
  XNOR U1623 ( .A(n1581), .B(n1582), .Z(n1547) );
  XNOR U1624 ( .A(n1568), .B(n1583), .Z(n1582) );
  XNOR U1625 ( .A(n1501), .B(n1562), .Z(n1583) );
  XOR U1626 ( .A(n1569), .B(n1584), .Z(n1562) );
  XNOR U1627 ( .A(n1585), .B(n1586), .Z(n1584) );
  NAND U1628 ( .A(n1528), .B(n1498), .Z(n1586) );
  XNOR U1629 ( .A(n1587), .B(n1585), .Z(n1569) );
  NANDN U1630 ( .A(n1530), .B(n1507), .Z(n1585) );
  XOR U1631 ( .A(n1508), .B(n1498), .Z(n1507) );
  XNOR U1632 ( .A(n1588), .B(n1471), .Z(n1498) );
  XOR U1633 ( .A(n1539), .B(n1528), .Z(n1530) );
  XOR U1634 ( .A(n1519), .B(n1589), .Z(n1528) );
  ANDN U1635 ( .B(n1508), .A(n1539), .Z(n1587) );
  XOR U1636 ( .A(n1577), .B(n1524), .Z(n1539) );
  XOR U1637 ( .A(n1590), .B(n1591), .Z(n1524) );
  XOR U1638 ( .A(n1592), .B(n1593), .Z(n1591) );
  XOR U1639 ( .A(n1594), .B(n1576), .Z(n1508) );
  XOR U1640 ( .A(n1589), .B(n1572), .Z(n1568) );
  IV U1641 ( .A(n1471), .Z(n1572) );
  XOR U1642 ( .A(n1595), .B(n1596), .Z(n1471) );
  XNOR U1643 ( .A(n1597), .B(n1593), .Z(n1596) );
  IV U1644 ( .A(n1514), .Z(n1589) );
  XOR U1645 ( .A(n1593), .B(n1598), .Z(n1514) );
  XNOR U1646 ( .A(n1519), .B(n1599), .Z(n1581) );
  XNOR U1647 ( .A(n1600), .B(n1580), .Z(n1599) );
  OR U1648 ( .A(n1504), .B(n1518), .Z(n1580) );
  XNOR U1649 ( .A(n1577), .B(n1519), .Z(n1518) );
  XOR U1650 ( .A(n1493), .B(n1588), .Z(n1504) );
  IV U1651 ( .A(n1501), .Z(n1588) );
  XOR U1652 ( .A(n1576), .B(n1601), .Z(n1501) );
  XNOR U1653 ( .A(n1597), .B(n1590), .Z(n1601) );
  XOR U1654 ( .A(key[194]), .B(\w0[1][66] ), .Z(n1590) );
  XOR U1655 ( .A(n1602), .B(n1603), .Z(\w0[1][66] ) );
  XNOR U1656 ( .A(n219), .B(n1604), .Z(n1603) );
  IV U1657 ( .A(n1483), .Z(n1576) );
  XOR U1658 ( .A(n1595), .B(n1605), .Z(n1483) );
  XOR U1659 ( .A(n1593), .B(n1606), .Z(n1605) );
  ANDN U1660 ( .B(n1594), .A(n1464), .Z(n1600) );
  IV U1661 ( .A(n1493), .Z(n1594) );
  XOR U1662 ( .A(n1595), .B(n1607), .Z(n1493) );
  XOR U1663 ( .A(n1593), .B(n1608), .Z(n1607) );
  XOR U1664 ( .A(n1464), .B(n1609), .Z(n1593) );
  XOR U1665 ( .A(key[198]), .B(\w0[1][70] ), .Z(n1609) );
  XNOR U1666 ( .A(n1610), .B(n1611), .Z(\w0[1][70] ) );
  XOR U1667 ( .A(n187), .B(n192), .Z(n1611) );
  XNOR U1668 ( .A(n1612), .B(n1613), .Z(n187) );
  IV U1669 ( .A(n1577), .Z(n1464) );
  IV U1670 ( .A(n1598), .Z(n1595) );
  XOR U1671 ( .A(key[197]), .B(\w0[1][69] ), .Z(n1598) );
  XOR U1672 ( .A(n1614), .B(n1615), .Z(\w0[1][69] ) );
  XOR U1673 ( .A(n191), .B(n1616), .Z(n1615) );
  XNOR U1674 ( .A(n1617), .B(n1618), .Z(n191) );
  XOR U1675 ( .A(n1619), .B(n1620), .Z(n1519) );
  XNOR U1676 ( .A(n1608), .B(n1606), .Z(n1620) );
  XNOR U1677 ( .A(key[199]), .B(\w0[1][71] ), .Z(n1606) );
  XOR U1678 ( .A(n1621), .B(n1622), .Z(\w0[1][71] ) );
  XOR U1679 ( .A(n200), .B(n1613), .Z(n1622) );
  XNOR U1680 ( .A(n1623), .B(n1624), .Z(n1613) );
  XOR U1681 ( .A(n1625), .B(n1626), .Z(n200) );
  XNOR U1682 ( .A(key[196]), .B(\w0[1][68] ), .Z(n1608) );
  XOR U1683 ( .A(n1627), .B(n1628), .Z(\w0[1][68] ) );
  XNOR U1684 ( .A(n1629), .B(n1630), .Z(n1628) );
  XNOR U1685 ( .A(n205), .B(n204), .Z(n1627) );
  XNOR U1686 ( .A(n1631), .B(n1632), .Z(n204) );
  XOR U1687 ( .A(n1633), .B(n1616), .Z(n205) );
  XNOR U1688 ( .A(n1577), .B(n1592), .Z(n1619) );
  XOR U1689 ( .A(n1597), .B(n1634), .Z(n1592) );
  XOR U1690 ( .A(key[195]), .B(\w0[1][67] ), .Z(n1634) );
  XOR U1691 ( .A(n1635), .B(n1636), .Z(\w0[1][67] ) );
  XNOR U1692 ( .A(n177), .B(n1637), .Z(n1636) );
  XNOR U1693 ( .A(n212), .B(n211), .Z(n1635) );
  XOR U1694 ( .A(n1633), .B(n1629), .Z(n212) );
  XOR U1695 ( .A(key[193]), .B(\w0[1][65] ), .Z(n1597) );
  XNOR U1696 ( .A(n1638), .B(n1639), .Z(\w0[1][65] ) );
  XOR U1697 ( .A(n217), .B(n223), .Z(n1639) );
  XOR U1698 ( .A(key[192]), .B(\w0[1][64] ), .Z(n1577) );
  XNOR U1699 ( .A(n1640), .B(n1641), .Z(\w0[1][64] ) );
  XNOR U1700 ( .A(n197), .B(n1642), .Z(n1641) );
  XOR U1701 ( .A(n1643), .B(n1644), .Z(out[31]) );
  XOR U1702 ( .A(n1645), .B(n1646), .Z(n1643) );
  XOR U1703 ( .A(key[159]), .B(n1647), .Z(n1646) );
  XNOR U1704 ( .A(n1648), .B(n1649), .Z(out[30]) );
  XNOR U1705 ( .A(key[158]), .B(n1650), .Z(n1649) );
  XOR U1706 ( .A(key[130]), .B(n1082), .Z(out[2]) );
  XOR U1707 ( .A(n1652), .B(n1653), .Z(out[29]) );
  XNOR U1708 ( .A(n1654), .B(n1655), .Z(n1653) );
  XOR U1709 ( .A(n1645), .B(n1656), .Z(n1655) );
  XNOR U1710 ( .A(n1658), .B(n1659), .Z(n1657) );
  NANDN U1711 ( .A(n1660), .B(n1661), .Z(n1659) );
  XOR U1712 ( .A(n1663), .B(n1664), .Z(n1652) );
  XOR U1713 ( .A(key[157]), .B(n1665), .Z(n1664) );
  ANDN U1714 ( .B(n1666), .A(n1667), .Z(n1663) );
  XNOR U1715 ( .A(n1668), .B(n1669), .Z(out[28]) );
  XNOR U1716 ( .A(key[156]), .B(n1670), .Z(n1669) );
  XOR U1717 ( .A(n1671), .B(n1672), .Z(out[27]) );
  XNOR U1718 ( .A(n1673), .B(n1648), .Z(n1672) );
  XNOR U1719 ( .A(n1674), .B(n1675), .Z(n1648) );
  XNOR U1720 ( .A(n1676), .B(n1665), .Z(n1675) );
  ANDN U1721 ( .B(n1677), .A(n1678), .Z(n1665) );
  NOR U1722 ( .A(n1679), .B(n1680), .Z(n1676) );
  XNOR U1723 ( .A(n1681), .B(n1682), .Z(n1671) );
  XOR U1724 ( .A(key[155]), .B(n1647), .Z(n1682) );
  XOR U1725 ( .A(key[154]), .B(n1668), .Z(out[26]) );
  XNOR U1726 ( .A(n1683), .B(n1684), .Z(n1668) );
  XOR U1727 ( .A(n1685), .B(n1644), .Z(out[25]) );
  XNOR U1728 ( .A(n1674), .B(n1686), .Z(n1673) );
  XNOR U1729 ( .A(n1687), .B(n1688), .Z(n1686) );
  NANDN U1730 ( .A(n1689), .B(n1661), .Z(n1688) );
  XNOR U1731 ( .A(n1656), .B(n1690), .Z(n1674) );
  XNOR U1732 ( .A(n1691), .B(n1692), .Z(n1690) );
  NANDN U1733 ( .A(n1693), .B(n1694), .Z(n1692) );
  XOR U1734 ( .A(n1684), .B(n1681), .Z(n1650) );
  XNOR U1735 ( .A(n1656), .B(n1695), .Z(n1681) );
  XNOR U1736 ( .A(n1687), .B(n1696), .Z(n1695) );
  NANDN U1737 ( .A(n1697), .B(n1698), .Z(n1696) );
  OR U1738 ( .A(n1699), .B(n1700), .Z(n1687) );
  XOR U1739 ( .A(n1701), .B(n1691), .Z(n1656) );
  NANDN U1740 ( .A(n1702), .B(n1703), .Z(n1691) );
  ANDN U1741 ( .B(n1704), .A(n1705), .Z(n1701) );
  XNOR U1742 ( .A(key[153]), .B(n1683), .Z(n1685) );
  IV U1743 ( .A(n1647), .Z(n1683) );
  XOR U1744 ( .A(n1706), .B(n1707), .Z(n1647) );
  XNOR U1745 ( .A(n1708), .B(n1709), .Z(n1707) );
  NAND U1746 ( .A(n1666), .B(n1710), .Z(n1709) );
  XNOR U1747 ( .A(n1654), .B(n1711), .Z(out[24]) );
  XOR U1748 ( .A(key[152]), .B(n1684), .Z(n1711) );
  XNOR U1749 ( .A(n1706), .B(n1712), .Z(n1684) );
  XOR U1750 ( .A(n1713), .B(n1658), .Z(n1712) );
  OR U1751 ( .A(n1714), .B(n1699), .Z(n1658) );
  XNOR U1752 ( .A(n1661), .B(n1698), .Z(n1699) );
  ANDN U1753 ( .B(n1715), .A(n1716), .Z(n1713) );
  IV U1754 ( .A(n1670), .Z(n1654) );
  XOR U1755 ( .A(n1662), .B(n1717), .Z(n1670) );
  XOR U1756 ( .A(n1718), .B(n1708), .Z(n1717) );
  XNOR U1757 ( .A(n1680), .B(n1666), .Z(n1677) );
  NOR U1758 ( .A(n1720), .B(n1680), .Z(n1718) );
  XNOR U1759 ( .A(n1706), .B(n1721), .Z(n1662) );
  XNOR U1760 ( .A(n1722), .B(n1723), .Z(n1721) );
  NANDN U1761 ( .A(n1693), .B(n1724), .Z(n1723) );
  XOR U1762 ( .A(n1725), .B(n1722), .Z(n1706) );
  OR U1763 ( .A(n1702), .B(n1726), .Z(n1722) );
  XOR U1764 ( .A(n1727), .B(n1693), .Z(n1702) );
  XNOR U1765 ( .A(n1698), .B(n1666), .Z(n1693) );
  XOR U1766 ( .A(n1728), .B(n1729), .Z(n1666) );
  NANDN U1767 ( .A(n1730), .B(n1731), .Z(n1729) );
  IV U1768 ( .A(n1716), .Z(n1698) );
  XNOR U1769 ( .A(n1732), .B(n1733), .Z(n1716) );
  NANDN U1770 ( .A(n1730), .B(n1734), .Z(n1733) );
  ANDN U1771 ( .B(n1727), .A(n1735), .Z(n1725) );
  IV U1772 ( .A(n1705), .Z(n1727) );
  XOR U1773 ( .A(n1680), .B(n1661), .Z(n1705) );
  XNOR U1774 ( .A(n1736), .B(n1732), .Z(n1661) );
  NANDN U1775 ( .A(n1737), .B(n1738), .Z(n1732) );
  XOR U1776 ( .A(n1734), .B(n1739), .Z(n1738) );
  ANDN U1777 ( .B(n1739), .A(n1740), .Z(n1736) );
  XOR U1778 ( .A(n1741), .B(n1728), .Z(n1680) );
  NANDN U1779 ( .A(n1737), .B(n1742), .Z(n1728) );
  XOR U1780 ( .A(n1743), .B(n1731), .Z(n1742) );
  XNOR U1781 ( .A(n1744), .B(n1745), .Z(n1730) );
  XOR U1782 ( .A(n1746), .B(n1747), .Z(n1745) );
  XNOR U1783 ( .A(n1748), .B(n1749), .Z(n1744) );
  XNOR U1784 ( .A(n1750), .B(n1751), .Z(n1749) );
  ANDN U1785 ( .B(n1743), .A(n1747), .Z(n1750) );
  ANDN U1786 ( .B(n1743), .A(n1740), .Z(n1741) );
  XNOR U1787 ( .A(n1746), .B(n1752), .Z(n1740) );
  XOR U1788 ( .A(n1753), .B(n1751), .Z(n1752) );
  NAND U1789 ( .A(n1754), .B(n1755), .Z(n1751) );
  XNOR U1790 ( .A(n1748), .B(n1731), .Z(n1755) );
  IV U1791 ( .A(n1743), .Z(n1748) );
  XNOR U1792 ( .A(n1734), .B(n1747), .Z(n1754) );
  IV U1793 ( .A(n1739), .Z(n1747) );
  XOR U1794 ( .A(n1756), .B(n1757), .Z(n1739) );
  XNOR U1795 ( .A(n1758), .B(n1759), .Z(n1757) );
  XNOR U1796 ( .A(n1760), .B(n1761), .Z(n1756) );
  NOR U1797 ( .A(n1679), .B(n1720), .Z(n1760) );
  AND U1798 ( .A(n1731), .B(n1734), .Z(n1753) );
  XNOR U1799 ( .A(n1731), .B(n1734), .Z(n1746) );
  XNOR U1800 ( .A(n1762), .B(n1763), .Z(n1734) );
  XNOR U1801 ( .A(n1764), .B(n1759), .Z(n1763) );
  XOR U1802 ( .A(n1765), .B(n1766), .Z(n1762) );
  XNOR U1803 ( .A(n1767), .B(n1761), .Z(n1766) );
  OR U1804 ( .A(n1678), .B(n1719), .Z(n1761) );
  XOR U1805 ( .A(n1720), .B(n1710), .Z(n1719) );
  XNOR U1806 ( .A(n1679), .B(n1667), .Z(n1678) );
  ANDN U1807 ( .B(n1710), .A(n1667), .Z(n1767) );
  XNOR U1808 ( .A(n1768), .B(n1769), .Z(n1731) );
  XNOR U1809 ( .A(n1759), .B(n1770), .Z(n1769) );
  XOR U1810 ( .A(n1689), .B(n1765), .Z(n1770) );
  XNOR U1811 ( .A(n1720), .B(n1771), .Z(n1759) );
  XNOR U1812 ( .A(n1772), .B(n1773), .Z(n1768) );
  XNOR U1813 ( .A(n1774), .B(n1775), .Z(n1773) );
  ANDN U1814 ( .B(n1715), .A(n1697), .Z(n1774) );
  XNOR U1815 ( .A(n1776), .B(n1777), .Z(n1743) );
  XNOR U1816 ( .A(n1764), .B(n1778), .Z(n1777) );
  XNOR U1817 ( .A(n1697), .B(n1758), .Z(n1778) );
  XOR U1818 ( .A(n1765), .B(n1779), .Z(n1758) );
  XNOR U1819 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1820 ( .A(n1724), .B(n1694), .Z(n1781) );
  XNOR U1821 ( .A(n1782), .B(n1780), .Z(n1765) );
  NANDN U1822 ( .A(n1726), .B(n1703), .Z(n1780) );
  XOR U1823 ( .A(n1704), .B(n1694), .Z(n1703) );
  XNOR U1824 ( .A(n1783), .B(n1667), .Z(n1694) );
  XOR U1825 ( .A(n1735), .B(n1724), .Z(n1726) );
  XOR U1826 ( .A(n1715), .B(n1710), .Z(n1724) );
  ANDN U1827 ( .B(n1704), .A(n1735), .Z(n1782) );
  XOR U1828 ( .A(n1772), .B(n1720), .Z(n1735) );
  XOR U1829 ( .A(n1784), .B(n1785), .Z(n1720) );
  XOR U1830 ( .A(n1786), .B(n1787), .Z(n1785) );
  XOR U1831 ( .A(n1788), .B(n1771), .Z(n1704) );
  XNOR U1832 ( .A(n1789), .B(n1790), .Z(n1667) );
  XNOR U1833 ( .A(n1791), .B(n1787), .Z(n1790) );
  XNOR U1834 ( .A(n1787), .B(n1789), .Z(n1710) );
  XNOR U1835 ( .A(n1715), .B(n1792), .Z(n1776) );
  XNOR U1836 ( .A(n1793), .B(n1775), .Z(n1792) );
  OR U1837 ( .A(n1700), .B(n1714), .Z(n1775) );
  XNOR U1838 ( .A(n1772), .B(n1715), .Z(n1714) );
  XOR U1839 ( .A(n1689), .B(n1783), .Z(n1700) );
  IV U1840 ( .A(n1697), .Z(n1783) );
  XOR U1841 ( .A(n1771), .B(n1794), .Z(n1697) );
  XNOR U1842 ( .A(n1791), .B(n1784), .Z(n1794) );
  XOR U1843 ( .A(key[154]), .B(\w0[1][26] ), .Z(n1784) );
  XOR U1844 ( .A(n1795), .B(n1796), .Z(\w0[1][26] ) );
  XOR U1845 ( .A(n615), .B(n1232), .Z(n1796) );
  XNOR U1846 ( .A(n619), .B(n1797), .Z(n1795) );
  IV U1847 ( .A(n1679), .Z(n1771) );
  XNOR U1848 ( .A(n1789), .B(n1798), .Z(n1679) );
  XNOR U1849 ( .A(n1787), .B(n1799), .Z(n1798) );
  ANDN U1850 ( .B(n1788), .A(n1660), .Z(n1793) );
  IV U1851 ( .A(n1689), .Z(n1788) );
  XNOR U1852 ( .A(n1789), .B(n1800), .Z(n1689) );
  XNOR U1853 ( .A(n1787), .B(n1801), .Z(n1800) );
  XOR U1854 ( .A(n1660), .B(n1802), .Z(n1787) );
  XOR U1855 ( .A(key[158]), .B(\w0[1][30] ), .Z(n1802) );
  XNOR U1856 ( .A(n1203), .B(n1803), .Z(\w0[1][30] ) );
  XNOR U1857 ( .A(n1804), .B(n596), .Z(n1803) );
  XOR U1858 ( .A(n1805), .B(n589), .Z(n1203) );
  IV U1859 ( .A(n1772), .Z(n1660) );
  XOR U1860 ( .A(key[157]), .B(\w0[1][29] ), .Z(n1789) );
  XOR U1861 ( .A(n1806), .B(n1807), .Z(\w0[1][29] ) );
  XOR U1862 ( .A(n1808), .B(n1210), .Z(n1807) );
  XOR U1863 ( .A(n602), .B(n1809), .Z(n1806) );
  XOR U1864 ( .A(n1810), .B(n1811), .Z(n1715) );
  XNOR U1865 ( .A(n1801), .B(n1799), .Z(n1811) );
  XOR U1866 ( .A(key[159]), .B(\w0[1][31] ), .Z(n1799) );
  XNOR U1867 ( .A(n1218), .B(n1812), .Z(\w0[1][31] ) );
  XOR U1868 ( .A(n608), .B(n1813), .Z(n1812) );
  XOR U1869 ( .A(key[156]), .B(\w0[1][28] ), .Z(n1801) );
  XOR U1870 ( .A(n1814), .B(n1815), .Z(\w0[1][28] ) );
  XNOR U1871 ( .A(n1805), .B(n593), .Z(n1221) );
  XNOR U1872 ( .A(n1816), .B(n1817), .Z(n1814) );
  XNOR U1873 ( .A(n1772), .B(n1786), .Z(n1810) );
  XOR U1874 ( .A(n1791), .B(n1818), .Z(n1786) );
  XOR U1875 ( .A(key[155]), .B(\w0[1][27] ), .Z(n1818) );
  XOR U1876 ( .A(n1819), .B(n1820), .Z(\w0[1][27] ) );
  XOR U1877 ( .A(n624), .B(n1230), .Z(n1820) );
  XOR U1878 ( .A(n1214), .B(n581), .Z(n1230) );
  XOR U1879 ( .A(n1821), .B(n1196), .Z(n1819) );
  XOR U1880 ( .A(key[153]), .B(\w0[1][25] ), .Z(n1791) );
  XOR U1881 ( .A(n1822), .B(n1823), .Z(\w0[1][25] ) );
  XOR U1882 ( .A(n626), .B(n1236), .Z(n1823) );
  XOR U1883 ( .A(n607), .B(n1824), .Z(n1822) );
  XOR U1884 ( .A(key[152]), .B(\w0[1][24] ), .Z(n1772) );
  XOR U1885 ( .A(n1825), .B(n1826), .Z(\w0[1][24] ) );
  XNOR U1886 ( .A(n1805), .B(n590), .Z(n1826) );
  XNOR U1887 ( .A(n605), .B(n1216), .Z(n590) );
  XOR U1888 ( .A(n1827), .B(n618), .Z(n1825) );
  XOR U1889 ( .A(n1828), .B(n1829), .Z(out[23]) );
  XOR U1890 ( .A(n1830), .B(n1831), .Z(n1828) );
  XOR U1891 ( .A(key[151]), .B(n1832), .Z(n1831) );
  XNOR U1892 ( .A(n1833), .B(n1834), .Z(out[22]) );
  XNOR U1893 ( .A(key[150]), .B(n1835), .Z(n1834) );
  XOR U1894 ( .A(n1836), .B(n1837), .Z(out[21]) );
  XNOR U1895 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U1896 ( .A(n1830), .B(n1840), .Z(n1839) );
  XNOR U1897 ( .A(n1842), .B(n1843), .Z(n1841) );
  NANDN U1898 ( .A(n1844), .B(n1845), .Z(n1843) );
  XOR U1899 ( .A(n1847), .B(n1848), .Z(n1836) );
  XOR U1900 ( .A(key[149]), .B(n1849), .Z(n1848) );
  ANDN U1901 ( .B(n1850), .A(n1851), .Z(n1847) );
  XNOR U1902 ( .A(n1852), .B(n1853), .Z(out[20]) );
  XNOR U1903 ( .A(key[148]), .B(n1854), .Z(n1853) );
  XOR U1904 ( .A(n1855), .B(n422), .Z(out[1]) );
  XNOR U1905 ( .A(n1439), .B(n1856), .Z(n1438) );
  XNOR U1906 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1907 ( .A(n1859), .B(n861), .Z(n1858) );
  XNOR U1908 ( .A(n856), .B(n1860), .Z(n1439) );
  XNOR U1909 ( .A(n1861), .B(n1862), .Z(n1860) );
  NANDN U1910 ( .A(n1863), .B(n1864), .Z(n1862) );
  XOR U1911 ( .A(n1651), .B(n1446), .Z(n640) );
  XNOR U1912 ( .A(n856), .B(n1865), .Z(n1446) );
  XNOR U1913 ( .A(n1857), .B(n1866), .Z(n1865) );
  NANDN U1914 ( .A(n1867), .B(n1868), .Z(n1866) );
  OR U1915 ( .A(n1869), .B(n1870), .Z(n1857) );
  XOR U1916 ( .A(n1871), .B(n1861), .Z(n856) );
  NANDN U1917 ( .A(n1872), .B(n1873), .Z(n1861) );
  ANDN U1918 ( .B(n1874), .A(n1875), .Z(n1871) );
  XOR U1919 ( .A(key[129]), .B(n425), .Z(n1855) );
  XOR U1920 ( .A(n1876), .B(n1877), .Z(n425) );
  XNOR U1921 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1922 ( .A(n866), .B(n1880), .Z(n1879) );
  XOR U1923 ( .A(n1881), .B(n1882), .Z(out[19]) );
  XNOR U1924 ( .A(n1883), .B(n1833), .Z(n1882) );
  XNOR U1925 ( .A(n1884), .B(n1885), .Z(n1833) );
  XNOR U1926 ( .A(n1886), .B(n1849), .Z(n1885) );
  ANDN U1927 ( .B(n1887), .A(n1888), .Z(n1849) );
  NOR U1928 ( .A(n1889), .B(n1890), .Z(n1886) );
  XNOR U1929 ( .A(n1891), .B(n1892), .Z(n1881) );
  XOR U1930 ( .A(key[147]), .B(n1832), .Z(n1892) );
  XOR U1931 ( .A(key[146]), .B(n1852), .Z(out[18]) );
  XNOR U1932 ( .A(n1893), .B(n1894), .Z(n1852) );
  XOR U1933 ( .A(n1895), .B(n1829), .Z(out[17]) );
  XNOR U1934 ( .A(n1884), .B(n1896), .Z(n1883) );
  XNOR U1935 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1936 ( .A(n1899), .B(n1845), .Z(n1898) );
  XNOR U1937 ( .A(n1840), .B(n1900), .Z(n1884) );
  XNOR U1938 ( .A(n1901), .B(n1902), .Z(n1900) );
  NANDN U1939 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U1940 ( .A(n1894), .B(n1891), .Z(n1835) );
  XNOR U1941 ( .A(n1840), .B(n1905), .Z(n1891) );
  XNOR U1942 ( .A(n1897), .B(n1906), .Z(n1905) );
  NANDN U1943 ( .A(n1907), .B(n1908), .Z(n1906) );
  OR U1944 ( .A(n1909), .B(n1910), .Z(n1897) );
  XOR U1945 ( .A(n1911), .B(n1901), .Z(n1840) );
  NANDN U1946 ( .A(n1912), .B(n1913), .Z(n1901) );
  ANDN U1947 ( .B(n1914), .A(n1915), .Z(n1911) );
  XNOR U1948 ( .A(key[145]), .B(n1893), .Z(n1895) );
  IV U1949 ( .A(n1832), .Z(n1893) );
  XOR U1950 ( .A(n1916), .B(n1917), .Z(n1832) );
  XNOR U1951 ( .A(n1918), .B(n1919), .Z(n1917) );
  NAND U1952 ( .A(n1850), .B(n1920), .Z(n1919) );
  XNOR U1953 ( .A(n1838), .B(n1921), .Z(out[16]) );
  XOR U1954 ( .A(key[144]), .B(n1894), .Z(n1921) );
  XNOR U1955 ( .A(n1916), .B(n1922), .Z(n1894) );
  XOR U1956 ( .A(n1923), .B(n1842), .Z(n1922) );
  OR U1957 ( .A(n1924), .B(n1909), .Z(n1842) );
  XNOR U1958 ( .A(n1845), .B(n1908), .Z(n1909) );
  ANDN U1959 ( .B(n1925), .A(n1926), .Z(n1923) );
  IV U1960 ( .A(n1854), .Z(n1838) );
  XOR U1961 ( .A(n1846), .B(n1927), .Z(n1854) );
  XOR U1962 ( .A(n1928), .B(n1918), .Z(n1927) );
  XNOR U1963 ( .A(n1890), .B(n1850), .Z(n1887) );
  NOR U1964 ( .A(n1930), .B(n1890), .Z(n1928) );
  XNOR U1965 ( .A(n1916), .B(n1931), .Z(n1846) );
  XNOR U1966 ( .A(n1932), .B(n1933), .Z(n1931) );
  NANDN U1967 ( .A(n1903), .B(n1934), .Z(n1933) );
  XOR U1968 ( .A(n1935), .B(n1932), .Z(n1916) );
  OR U1969 ( .A(n1912), .B(n1936), .Z(n1932) );
  XOR U1970 ( .A(n1937), .B(n1903), .Z(n1912) );
  XNOR U1971 ( .A(n1908), .B(n1850), .Z(n1903) );
  XOR U1972 ( .A(n1938), .B(n1939), .Z(n1850) );
  NANDN U1973 ( .A(n1940), .B(n1941), .Z(n1939) );
  IV U1974 ( .A(n1926), .Z(n1908) );
  XNOR U1975 ( .A(n1942), .B(n1943), .Z(n1926) );
  NANDN U1976 ( .A(n1940), .B(n1944), .Z(n1943) );
  ANDN U1977 ( .B(n1937), .A(n1945), .Z(n1935) );
  IV U1978 ( .A(n1915), .Z(n1937) );
  XOR U1979 ( .A(n1890), .B(n1845), .Z(n1915) );
  XNOR U1980 ( .A(n1946), .B(n1942), .Z(n1845) );
  NANDN U1981 ( .A(n1947), .B(n1948), .Z(n1942) );
  XOR U1982 ( .A(n1944), .B(n1949), .Z(n1948) );
  ANDN U1983 ( .B(n1949), .A(n1950), .Z(n1946) );
  XOR U1984 ( .A(n1951), .B(n1938), .Z(n1890) );
  NANDN U1985 ( .A(n1947), .B(n1952), .Z(n1938) );
  XOR U1986 ( .A(n1953), .B(n1941), .Z(n1952) );
  XNOR U1987 ( .A(n1954), .B(n1955), .Z(n1940) );
  XOR U1988 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U1989 ( .A(n1958), .B(n1959), .Z(n1954) );
  XNOR U1990 ( .A(n1960), .B(n1961), .Z(n1959) );
  ANDN U1991 ( .B(n1953), .A(n1957), .Z(n1960) );
  ANDN U1992 ( .B(n1953), .A(n1950), .Z(n1951) );
  XNOR U1993 ( .A(n1956), .B(n1962), .Z(n1950) );
  XOR U1994 ( .A(n1963), .B(n1961), .Z(n1962) );
  NAND U1995 ( .A(n1964), .B(n1965), .Z(n1961) );
  XNOR U1996 ( .A(n1958), .B(n1941), .Z(n1965) );
  IV U1997 ( .A(n1953), .Z(n1958) );
  XNOR U1998 ( .A(n1944), .B(n1957), .Z(n1964) );
  IV U1999 ( .A(n1949), .Z(n1957) );
  XOR U2000 ( .A(n1966), .B(n1967), .Z(n1949) );
  XNOR U2001 ( .A(n1968), .B(n1969), .Z(n1967) );
  XNOR U2002 ( .A(n1970), .B(n1971), .Z(n1966) );
  NOR U2003 ( .A(n1889), .B(n1930), .Z(n1970) );
  AND U2004 ( .A(n1941), .B(n1944), .Z(n1963) );
  XNOR U2005 ( .A(n1941), .B(n1944), .Z(n1956) );
  XNOR U2006 ( .A(n1972), .B(n1973), .Z(n1944) );
  XNOR U2007 ( .A(n1974), .B(n1969), .Z(n1973) );
  XOR U2008 ( .A(n1975), .B(n1976), .Z(n1972) );
  XNOR U2009 ( .A(n1977), .B(n1971), .Z(n1976) );
  OR U2010 ( .A(n1888), .B(n1929), .Z(n1971) );
  XOR U2011 ( .A(n1930), .B(n1920), .Z(n1929) );
  XNOR U2012 ( .A(n1889), .B(n1851), .Z(n1888) );
  ANDN U2013 ( .B(n1920), .A(n1851), .Z(n1977) );
  XNOR U2014 ( .A(n1978), .B(n1979), .Z(n1941) );
  XNOR U2015 ( .A(n1969), .B(n1980), .Z(n1979) );
  XOR U2016 ( .A(n1899), .B(n1975), .Z(n1980) );
  XNOR U2017 ( .A(n1930), .B(n1981), .Z(n1969) );
  XNOR U2018 ( .A(n1982), .B(n1983), .Z(n1978) );
  XNOR U2019 ( .A(n1984), .B(n1985), .Z(n1983) );
  ANDN U2020 ( .B(n1925), .A(n1907), .Z(n1984) );
  XNOR U2021 ( .A(n1986), .B(n1987), .Z(n1953) );
  XNOR U2022 ( .A(n1974), .B(n1988), .Z(n1987) );
  XNOR U2023 ( .A(n1907), .B(n1968), .Z(n1988) );
  XOR U2024 ( .A(n1975), .B(n1989), .Z(n1968) );
  XNOR U2025 ( .A(n1990), .B(n1991), .Z(n1989) );
  NAND U2026 ( .A(n1934), .B(n1904), .Z(n1991) );
  XNOR U2027 ( .A(n1992), .B(n1990), .Z(n1975) );
  NANDN U2028 ( .A(n1936), .B(n1913), .Z(n1990) );
  XOR U2029 ( .A(n1914), .B(n1904), .Z(n1913) );
  XNOR U2030 ( .A(n1993), .B(n1851), .Z(n1904) );
  XOR U2031 ( .A(n1945), .B(n1934), .Z(n1936) );
  XOR U2032 ( .A(n1925), .B(n1920), .Z(n1934) );
  ANDN U2033 ( .B(n1914), .A(n1945), .Z(n1992) );
  XOR U2034 ( .A(n1982), .B(n1930), .Z(n1945) );
  XOR U2035 ( .A(n1994), .B(n1995), .Z(n1930) );
  XOR U2036 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U2037 ( .A(n1998), .B(n1981), .Z(n1914) );
  XNOR U2038 ( .A(n1999), .B(n2000), .Z(n1851) );
  XNOR U2039 ( .A(n2001), .B(n1997), .Z(n2000) );
  XNOR U2040 ( .A(n1997), .B(n1999), .Z(n1920) );
  XNOR U2041 ( .A(n1925), .B(n2002), .Z(n1986) );
  XNOR U2042 ( .A(n2003), .B(n1985), .Z(n2002) );
  OR U2043 ( .A(n1910), .B(n1924), .Z(n1985) );
  XNOR U2044 ( .A(n1982), .B(n1925), .Z(n1924) );
  XOR U2045 ( .A(n1899), .B(n1993), .Z(n1910) );
  IV U2046 ( .A(n1907), .Z(n1993) );
  XOR U2047 ( .A(n1981), .B(n2004), .Z(n1907) );
  XNOR U2048 ( .A(n2001), .B(n1994), .Z(n2004) );
  XOR U2049 ( .A(key[242]), .B(\w0[1][114] ), .Z(n1994) );
  XNOR U2050 ( .A(n811), .B(n2005), .Z(\w0[1][114] ) );
  XOR U2051 ( .A(n2006), .B(n2007), .Z(n2005) );
  XOR U2052 ( .A(n2008), .B(n814), .Z(n811) );
  IV U2053 ( .A(n1889), .Z(n1981) );
  XNOR U2054 ( .A(n1999), .B(n2009), .Z(n1889) );
  XNOR U2055 ( .A(n1997), .B(n2010), .Z(n2009) );
  ANDN U2056 ( .B(n1998), .A(n1844), .Z(n2003) );
  IV U2057 ( .A(n1899), .Z(n1998) );
  XNOR U2058 ( .A(n1999), .B(n2011), .Z(n1899) );
  XNOR U2059 ( .A(n1997), .B(n2012), .Z(n2011) );
  XOR U2060 ( .A(n1844), .B(n2013), .Z(n1997) );
  XOR U2061 ( .A(key[246]), .B(\w0[1][118] ), .Z(n2013) );
  XNOR U2062 ( .A(n1400), .B(n2014), .Z(\w0[1][118] ) );
  XNOR U2063 ( .A(n1407), .B(n2015), .Z(n2014) );
  XNOR U2064 ( .A(n2016), .B(n796), .Z(n1400) );
  XOR U2065 ( .A(n1408), .B(n820), .Z(n796) );
  IV U2066 ( .A(n1982), .Z(n1844) );
  XOR U2067 ( .A(key[245]), .B(\w0[1][117] ), .Z(n1999) );
  XNOR U2068 ( .A(n1406), .B(n2017), .Z(\w0[1][117] ) );
  XOR U2069 ( .A(n2018), .B(n2019), .Z(n2017) );
  XNOR U2070 ( .A(n1418), .B(n799), .Z(n1406) );
  XOR U2071 ( .A(n2020), .B(n2021), .Z(n1925) );
  XNOR U2072 ( .A(n2012), .B(n2010), .Z(n2021) );
  XOR U2073 ( .A(key[247]), .B(\w0[1][119] ), .Z(n2010) );
  XNOR U2074 ( .A(n1411), .B(n2022), .Z(\w0[1][119] ) );
  XOR U2075 ( .A(n2023), .B(n2016), .Z(n2022) );
  XNOR U2076 ( .A(n823), .B(n2024), .Z(n2016) );
  XOR U2077 ( .A(n1402), .B(n2025), .Z(n1411) );
  XOR U2078 ( .A(key[244]), .B(\w0[1][116] ), .Z(n2012) );
  XOR U2079 ( .A(n2026), .B(n2027), .Z(\w0[1][116] ) );
  XOR U2080 ( .A(n1420), .B(n1417), .Z(n2027) );
  XNOR U2081 ( .A(n1426), .B(n785), .Z(n1417) );
  XOR U2082 ( .A(n823), .B(n2019), .Z(n1420) );
  XNOR U2083 ( .A(n2028), .B(n2029), .Z(n2026) );
  XNOR U2084 ( .A(n1982), .B(n1996), .Z(n2020) );
  XOR U2085 ( .A(n2001), .B(n2030), .Z(n1996) );
  XOR U2086 ( .A(key[243]), .B(\w0[1][115] ), .Z(n2030) );
  XOR U2087 ( .A(n2031), .B(n2032), .Z(\w0[1][115] ) );
  XNOR U2088 ( .A(n2033), .B(n1424), .Z(n2032) );
  XOR U2089 ( .A(n823), .B(n2029), .Z(n1424) );
  XOR U2090 ( .A(n1391), .B(n812), .Z(n2031) );
  XOR U2091 ( .A(n805), .B(n1390), .Z(n812) );
  XOR U2092 ( .A(key[241]), .B(\w0[1][113] ), .Z(n2001) );
  XNOR U2093 ( .A(n824), .B(n2034), .Z(\w0[1][113] ) );
  XNOR U2094 ( .A(n815), .B(n1435), .Z(n2034) );
  XOR U2095 ( .A(n808), .B(n1434), .Z(n824) );
  XOR U2096 ( .A(key[240]), .B(\w0[1][112] ), .Z(n1982) );
  XNOR U2097 ( .A(n1414), .B(n2035), .Z(\w0[1][112] ) );
  XNOR U2098 ( .A(n2036), .B(n810), .Z(n2035) );
  XOR U2099 ( .A(n2037), .B(n2038), .Z(out[15]) );
  XNOR U2100 ( .A(n4), .B(n2039), .Z(n2038) );
  XNOR U2101 ( .A(n3), .B(n2040), .Z(n2037) );
  XOR U2102 ( .A(key[143]), .B(n5), .Z(n2040) );
  XNOR U2103 ( .A(n2041), .B(n2042), .Z(out[14]) );
  XOR U2104 ( .A(key[142]), .B(n3), .Z(n2042) );
  XOR U2105 ( .A(n63), .B(n2043), .Z(n3) );
  IV U2106 ( .A(n2044), .Z(n63) );
  XOR U2107 ( .A(n2045), .B(n2046), .Z(out[13]) );
  XNOR U2108 ( .A(n2039), .B(n2047), .Z(n2046) );
  XNOR U2109 ( .A(n2048), .B(n61), .Z(n2047) );
  XNOR U2110 ( .A(n2049), .B(n2050), .Z(n2039) );
  XNOR U2111 ( .A(n2051), .B(n2052), .Z(n2050) );
  OR U2112 ( .A(n2053), .B(n2054), .Z(n2052) );
  XOR U2113 ( .A(n2055), .B(n2056), .Z(n2045) );
  XOR U2114 ( .A(key[141]), .B(n2057), .Z(n2056) );
  AND U2115 ( .A(n2058), .B(n2059), .Z(n2055) );
  XNOR U2116 ( .A(n2060), .B(n2061), .Z(out[12]) );
  XOR U2117 ( .A(key[140]), .B(n61), .Z(n2061) );
  XNOR U2118 ( .A(n2049), .B(n2062), .Z(n61) );
  XOR U2119 ( .A(n2063), .B(n2064), .Z(n2062) );
  ANDN U2120 ( .B(n2065), .A(n2066), .Z(n2063) );
  XNOR U2121 ( .A(n2067), .B(n2068), .Z(n2049) );
  XNOR U2122 ( .A(n2069), .B(n2070), .Z(n2068) );
  NAND U2123 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U2124 ( .A(n2073), .B(n2074), .Z(out[127]) );
  XOR U2125 ( .A(n2075), .B(n2076), .Z(n2073) );
  XOR U2126 ( .A(key[255]), .B(n2077), .Z(n2076) );
  XNOR U2127 ( .A(n2078), .B(n2079), .Z(out[126]) );
  XNOR U2128 ( .A(key[254]), .B(n2080), .Z(n2079) );
  XOR U2129 ( .A(n2081), .B(n2082), .Z(out[125]) );
  XNOR U2130 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U2131 ( .A(n2075), .B(n2085), .Z(n2084) );
  XNOR U2132 ( .A(n2087), .B(n2088), .Z(n2086) );
  NANDN U2133 ( .A(n2089), .B(n2090), .Z(n2088) );
  XOR U2134 ( .A(n2092), .B(n2093), .Z(n2081) );
  XOR U2135 ( .A(key[253]), .B(n2094), .Z(n2093) );
  ANDN U2136 ( .B(n2095), .A(n2096), .Z(n2092) );
  XNOR U2137 ( .A(n2097), .B(n2098), .Z(out[124]) );
  XNOR U2138 ( .A(key[252]), .B(n2099), .Z(n2098) );
  XOR U2139 ( .A(n2100), .B(n2101), .Z(out[123]) );
  XNOR U2140 ( .A(n2102), .B(n2078), .Z(n2101) );
  XNOR U2141 ( .A(n2103), .B(n2104), .Z(n2078) );
  XNOR U2142 ( .A(n2105), .B(n2094), .Z(n2104) );
  ANDN U2143 ( .B(n2106), .A(n2107), .Z(n2094) );
  NOR U2144 ( .A(n2108), .B(n2109), .Z(n2105) );
  XNOR U2145 ( .A(n2110), .B(n2111), .Z(n2100) );
  XOR U2146 ( .A(key[251]), .B(n2077), .Z(n2111) );
  XOR U2147 ( .A(key[250]), .B(n2097), .Z(out[122]) );
  XNOR U2148 ( .A(n2112), .B(n2113), .Z(n2097) );
  XOR U2149 ( .A(n2114), .B(n2074), .Z(out[121]) );
  XNOR U2150 ( .A(n2103), .B(n2115), .Z(n2102) );
  XNOR U2151 ( .A(n2116), .B(n2117), .Z(n2115) );
  NANDN U2152 ( .A(n2118), .B(n2090), .Z(n2117) );
  XNOR U2153 ( .A(n2085), .B(n2119), .Z(n2103) );
  XNOR U2154 ( .A(n2120), .B(n2121), .Z(n2119) );
  NANDN U2155 ( .A(n2122), .B(n2123), .Z(n2121) );
  XOR U2156 ( .A(n2113), .B(n2110), .Z(n2080) );
  XNOR U2157 ( .A(n2085), .B(n2124), .Z(n2110) );
  XNOR U2158 ( .A(n2116), .B(n2125), .Z(n2124) );
  NANDN U2159 ( .A(n2126), .B(n2127), .Z(n2125) );
  OR U2160 ( .A(n2128), .B(n2129), .Z(n2116) );
  XOR U2161 ( .A(n2130), .B(n2120), .Z(n2085) );
  NANDN U2162 ( .A(n2131), .B(n2132), .Z(n2120) );
  ANDN U2163 ( .B(n2133), .A(n2134), .Z(n2130) );
  XNOR U2164 ( .A(key[249]), .B(n2112), .Z(n2114) );
  IV U2165 ( .A(n2077), .Z(n2112) );
  XOR U2166 ( .A(n2135), .B(n2136), .Z(n2077) );
  XNOR U2167 ( .A(n2137), .B(n2138), .Z(n2136) );
  NAND U2168 ( .A(n2095), .B(n2139), .Z(n2138) );
  XNOR U2169 ( .A(n2083), .B(n2140), .Z(out[120]) );
  XOR U2170 ( .A(key[248]), .B(n2113), .Z(n2140) );
  XNOR U2171 ( .A(n2135), .B(n2141), .Z(n2113) );
  XOR U2172 ( .A(n2142), .B(n2087), .Z(n2141) );
  OR U2173 ( .A(n2143), .B(n2128), .Z(n2087) );
  XNOR U2174 ( .A(n2090), .B(n2127), .Z(n2128) );
  ANDN U2175 ( .B(n2144), .A(n2145), .Z(n2142) );
  IV U2176 ( .A(n2099), .Z(n2083) );
  XOR U2177 ( .A(n2091), .B(n2146), .Z(n2099) );
  XOR U2178 ( .A(n2147), .B(n2137), .Z(n2146) );
  XNOR U2179 ( .A(n2109), .B(n2095), .Z(n2106) );
  NOR U2180 ( .A(n2149), .B(n2109), .Z(n2147) );
  XNOR U2181 ( .A(n2135), .B(n2150), .Z(n2091) );
  XNOR U2182 ( .A(n2151), .B(n2152), .Z(n2150) );
  NANDN U2183 ( .A(n2122), .B(n2153), .Z(n2152) );
  XOR U2184 ( .A(n2154), .B(n2151), .Z(n2135) );
  OR U2185 ( .A(n2131), .B(n2155), .Z(n2151) );
  XOR U2186 ( .A(n2156), .B(n2122), .Z(n2131) );
  XNOR U2187 ( .A(n2127), .B(n2095), .Z(n2122) );
  XOR U2188 ( .A(n2157), .B(n2158), .Z(n2095) );
  NANDN U2189 ( .A(n2159), .B(n2160), .Z(n2158) );
  IV U2190 ( .A(n2145), .Z(n2127) );
  XNOR U2191 ( .A(n2161), .B(n2162), .Z(n2145) );
  NANDN U2192 ( .A(n2159), .B(n2163), .Z(n2162) );
  ANDN U2193 ( .B(n2156), .A(n2164), .Z(n2154) );
  IV U2194 ( .A(n2134), .Z(n2156) );
  XOR U2195 ( .A(n2109), .B(n2090), .Z(n2134) );
  XNOR U2196 ( .A(n2165), .B(n2161), .Z(n2090) );
  NANDN U2197 ( .A(n2166), .B(n2167), .Z(n2161) );
  XOR U2198 ( .A(n2163), .B(n2168), .Z(n2167) );
  ANDN U2199 ( .B(n2168), .A(n2169), .Z(n2165) );
  XOR U2200 ( .A(n2170), .B(n2157), .Z(n2109) );
  NANDN U2201 ( .A(n2166), .B(n2171), .Z(n2157) );
  XOR U2202 ( .A(n2172), .B(n2160), .Z(n2171) );
  XNOR U2203 ( .A(n2173), .B(n2174), .Z(n2159) );
  XOR U2204 ( .A(n2175), .B(n2176), .Z(n2174) );
  XNOR U2205 ( .A(n2177), .B(n2178), .Z(n2173) );
  XNOR U2206 ( .A(n2179), .B(n2180), .Z(n2178) );
  ANDN U2207 ( .B(n2172), .A(n2176), .Z(n2179) );
  ANDN U2208 ( .B(n2172), .A(n2169), .Z(n2170) );
  XNOR U2209 ( .A(n2175), .B(n2181), .Z(n2169) );
  XOR U2210 ( .A(n2182), .B(n2180), .Z(n2181) );
  NAND U2211 ( .A(n2183), .B(n2184), .Z(n2180) );
  XNOR U2212 ( .A(n2177), .B(n2160), .Z(n2184) );
  IV U2213 ( .A(n2172), .Z(n2177) );
  XNOR U2214 ( .A(n2163), .B(n2176), .Z(n2183) );
  IV U2215 ( .A(n2168), .Z(n2176) );
  XOR U2216 ( .A(n2185), .B(n2186), .Z(n2168) );
  XNOR U2217 ( .A(n2187), .B(n2188), .Z(n2186) );
  XNOR U2218 ( .A(n2189), .B(n2190), .Z(n2185) );
  NOR U2219 ( .A(n2108), .B(n2149), .Z(n2189) );
  AND U2220 ( .A(n2160), .B(n2163), .Z(n2182) );
  XNOR U2221 ( .A(n2160), .B(n2163), .Z(n2175) );
  XNOR U2222 ( .A(n2191), .B(n2192), .Z(n2163) );
  XNOR U2223 ( .A(n2193), .B(n2188), .Z(n2192) );
  XOR U2224 ( .A(n2194), .B(n2195), .Z(n2191) );
  XNOR U2225 ( .A(n2196), .B(n2190), .Z(n2195) );
  OR U2226 ( .A(n2107), .B(n2148), .Z(n2190) );
  XOR U2227 ( .A(n2149), .B(n2139), .Z(n2148) );
  XNOR U2228 ( .A(n2108), .B(n2096), .Z(n2107) );
  ANDN U2229 ( .B(n2139), .A(n2096), .Z(n2196) );
  XNOR U2230 ( .A(n2197), .B(n2198), .Z(n2160) );
  XNOR U2231 ( .A(n2188), .B(n2199), .Z(n2198) );
  XOR U2232 ( .A(n2118), .B(n2194), .Z(n2199) );
  XNOR U2233 ( .A(n2149), .B(n2200), .Z(n2188) );
  XNOR U2234 ( .A(n2201), .B(n2202), .Z(n2197) );
  XNOR U2235 ( .A(n2203), .B(n2204), .Z(n2202) );
  ANDN U2236 ( .B(n2144), .A(n2126), .Z(n2203) );
  XNOR U2237 ( .A(n2205), .B(n2206), .Z(n2172) );
  XNOR U2238 ( .A(n2193), .B(n2207), .Z(n2206) );
  XNOR U2239 ( .A(n2126), .B(n2187), .Z(n2207) );
  XOR U2240 ( .A(n2194), .B(n2208), .Z(n2187) );
  XNOR U2241 ( .A(n2209), .B(n2210), .Z(n2208) );
  NAND U2242 ( .A(n2153), .B(n2123), .Z(n2210) );
  XNOR U2243 ( .A(n2211), .B(n2209), .Z(n2194) );
  NANDN U2244 ( .A(n2155), .B(n2132), .Z(n2209) );
  XOR U2245 ( .A(n2133), .B(n2123), .Z(n2132) );
  XNOR U2246 ( .A(n2212), .B(n2096), .Z(n2123) );
  XOR U2247 ( .A(n2164), .B(n2153), .Z(n2155) );
  XOR U2248 ( .A(n2144), .B(n2139), .Z(n2153) );
  ANDN U2249 ( .B(n2133), .A(n2164), .Z(n2211) );
  XOR U2250 ( .A(n2201), .B(n2149), .Z(n2164) );
  XOR U2251 ( .A(n2213), .B(n2214), .Z(n2149) );
  XOR U2252 ( .A(n2215), .B(n2216), .Z(n2214) );
  XOR U2253 ( .A(n2217), .B(n2200), .Z(n2133) );
  XNOR U2254 ( .A(n2218), .B(n2219), .Z(n2096) );
  XNOR U2255 ( .A(n2220), .B(n2216), .Z(n2219) );
  XNOR U2256 ( .A(n2216), .B(n2218), .Z(n2139) );
  XNOR U2257 ( .A(n2144), .B(n2221), .Z(n2205) );
  XNOR U2258 ( .A(n2222), .B(n2204), .Z(n2221) );
  OR U2259 ( .A(n2129), .B(n2143), .Z(n2204) );
  XNOR U2260 ( .A(n2201), .B(n2144), .Z(n2143) );
  XOR U2261 ( .A(n2118), .B(n2212), .Z(n2129) );
  IV U2262 ( .A(n2126), .Z(n2212) );
  XOR U2263 ( .A(n2200), .B(n2223), .Z(n2126) );
  XNOR U2264 ( .A(n2220), .B(n2213), .Z(n2223) );
  XOR U2265 ( .A(key[250]), .B(\w0[1][122] ), .Z(n2213) );
  XOR U2266 ( .A(n2224), .B(n2225), .Z(\w0[1][122] ) );
  XNOR U2267 ( .A(n805), .B(n815), .Z(n2225) );
  XNOR U2268 ( .A(n2007), .B(n1392), .Z(n815) );
  IV U2269 ( .A(n1431), .Z(n2007) );
  XNOR U2270 ( .A(n2226), .B(n2227), .Z(n805) );
  XOR U2271 ( .A(n2228), .B(n2229), .Z(n2227) );
  XNOR U2272 ( .A(n2230), .B(n2231), .Z(n2226) );
  XOR U2273 ( .A(n2008), .B(n1425), .Z(n2224) );
  IV U2274 ( .A(n1430), .Z(n2008) );
  IV U2275 ( .A(n2108), .Z(n2200) );
  XNOR U2276 ( .A(n2218), .B(n2232), .Z(n2108) );
  XNOR U2277 ( .A(n2216), .B(n2233), .Z(n2232) );
  ANDN U2278 ( .B(n2217), .A(n2089), .Z(n2222) );
  IV U2279 ( .A(n2118), .Z(n2217) );
  XNOR U2280 ( .A(n2218), .B(n2234), .Z(n2118) );
  XNOR U2281 ( .A(n2216), .B(n2235), .Z(n2234) );
  XOR U2282 ( .A(n2089), .B(n2236), .Z(n2216) );
  XOR U2283 ( .A(key[254]), .B(\w0[1][126] ), .Z(n2236) );
  XNOR U2284 ( .A(n2015), .B(n2237), .Z(\w0[1][126] ) );
  XOR U2285 ( .A(n2238), .B(n2239), .Z(n1408) );
  XNOR U2286 ( .A(n2018), .B(n792), .Z(n819) );
  XOR U2287 ( .A(n2036), .B(n2025), .Z(n792) );
  XNOR U2288 ( .A(n2240), .B(n2241), .Z(n2025) );
  XNOR U2289 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U2290 ( .A(n2230), .B(n2228), .Z(n2240) );
  IV U2291 ( .A(n2244), .Z(n2228) );
  XNOR U2292 ( .A(n1399), .B(n1407), .Z(n2018) );
  XNOR U2293 ( .A(n2245), .B(n2246), .Z(n1407) );
  XOR U2294 ( .A(n2247), .B(n1413), .Z(n2015) );
  IV U2295 ( .A(n2201), .Z(n2089) );
  XOR U2296 ( .A(key[253]), .B(\w0[1][125] ), .Z(n2218) );
  XOR U2297 ( .A(n2248), .B(n2249), .Z(\w0[1][125] ) );
  XNOR U2298 ( .A(n798), .B(n820), .Z(n2249) );
  XOR U2299 ( .A(n2231), .B(n2242), .Z(n820) );
  XOR U2300 ( .A(n2251), .B(n2252), .Z(n2250) );
  NOR U2301 ( .A(n2253), .B(n2254), .Z(n2251) );
  XNOR U2302 ( .A(n1405), .B(n2019), .Z(n798) );
  XNOR U2303 ( .A(n2256), .B(n2257), .Z(n2019) );
  XOR U2304 ( .A(n2258), .B(n2259), .Z(n2257) );
  XNOR U2305 ( .A(n2260), .B(n2261), .Z(n2256) );
  XOR U2306 ( .A(n2262), .B(n2263), .Z(n2261) );
  ANDN U2307 ( .B(n2264), .A(n2265), .Z(n2263) );
  XNOR U2308 ( .A(n1399), .B(n1418), .Z(n2248) );
  XNOR U2309 ( .A(n2266), .B(n2267), .Z(n1418) );
  XNOR U2310 ( .A(n2268), .B(n2269), .Z(n2267) );
  XNOR U2311 ( .A(n2270), .B(n2271), .Z(n2266) );
  XNOR U2312 ( .A(n2272), .B(n2273), .Z(n2271) );
  ANDN U2313 ( .B(n2274), .A(n2275), .Z(n2273) );
  XOR U2314 ( .A(n2276), .B(n2277), .Z(n1399) );
  XOR U2315 ( .A(n2278), .B(n2279), .Z(n2144) );
  XNOR U2316 ( .A(n2235), .B(n2233), .Z(n2279) );
  XOR U2317 ( .A(key[255]), .B(\w0[1][127] ), .Z(n2233) );
  XNOR U2318 ( .A(n795), .B(n2280), .Z(\w0[1][127] ) );
  XNOR U2319 ( .A(n821), .B(n1402), .Z(n2280) );
  XOR U2320 ( .A(n2281), .B(n2282), .Z(n1402) );
  XOR U2321 ( .A(n2239), .B(n2269), .Z(n2282) );
  XNOR U2322 ( .A(n2283), .B(n2284), .Z(n2269) );
  XNOR U2323 ( .A(n2285), .B(n2286), .Z(n2284) );
  OR U2324 ( .A(n2287), .B(n2288), .Z(n2286) );
  XOR U2325 ( .A(n2289), .B(n2290), .Z(n2281) );
  XOR U2326 ( .A(n2036), .B(n2023), .Z(n821) );
  XNOR U2327 ( .A(n1413), .B(n2024), .Z(n795) );
  XNOR U2328 ( .A(n2291), .B(n2292), .Z(n2024) );
  XOR U2329 ( .A(n2246), .B(n2259), .Z(n2292) );
  XNOR U2330 ( .A(n2293), .B(n2294), .Z(n2259) );
  XNOR U2331 ( .A(n2295), .B(n2296), .Z(n2294) );
  OR U2332 ( .A(n2297), .B(n2298), .Z(n2296) );
  XOR U2333 ( .A(n2299), .B(n2300), .Z(n2291) );
  XNOR U2334 ( .A(n2301), .B(n2302), .Z(n1413) );
  XNOR U2335 ( .A(n2277), .B(n2303), .Z(n2302) );
  XOR U2336 ( .A(n2304), .B(n2305), .Z(n2301) );
  XOR U2337 ( .A(key[252]), .B(\w0[1][124] ), .Z(n2235) );
  XOR U2338 ( .A(n2306), .B(n2307), .Z(\w0[1][124] ) );
  XOR U2339 ( .A(n2028), .B(n783), .Z(n2307) );
  XOR U2340 ( .A(n1419), .B(n2029), .Z(n783) );
  XOR U2341 ( .A(n1431), .B(n2258), .Z(n2029) );
  XOR U2342 ( .A(n2299), .B(n2308), .Z(n1431) );
  IV U2343 ( .A(n2309), .Z(n2299) );
  XOR U2344 ( .A(n2247), .B(n1405), .Z(n2028) );
  XNOR U2345 ( .A(n2310), .B(n2311), .Z(n1405) );
  XOR U2346 ( .A(n2312), .B(n2303), .Z(n2311) );
  XNOR U2347 ( .A(n2313), .B(n2314), .Z(n2303) );
  XNOR U2348 ( .A(n2315), .B(n2316), .Z(n2314) );
  OR U2349 ( .A(n2317), .B(n2318), .Z(n2316) );
  XNOR U2350 ( .A(n2319), .B(n2320), .Z(n2310) );
  XOR U2351 ( .A(n2321), .B(n2322), .Z(n2320) );
  ANDN U2352 ( .B(n2323), .A(n2324), .Z(n2322) );
  XOR U2353 ( .A(n1426), .B(n786), .Z(n2306) );
  XOR U2354 ( .A(n2036), .B(n799), .Z(n786) );
  XNOR U2355 ( .A(n2325), .B(n2326), .Z(n799) );
  XNOR U2356 ( .A(n2327), .B(n2243), .Z(n2326) );
  XNOR U2357 ( .A(n2328), .B(n2329), .Z(n2243) );
  XNOR U2358 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2359 ( .A(n2332), .B(n2333), .Z(n2331) );
  XNOR U2360 ( .A(n2334), .B(n2335), .Z(n2325) );
  XNOR U2361 ( .A(n2252), .B(n2336), .Z(n2335) );
  ANDN U2362 ( .B(n2337), .A(n2338), .Z(n2336) );
  NANDN U2363 ( .A(n2339), .B(n2340), .Z(n2252) );
  XOR U2364 ( .A(n2270), .B(n1430), .Z(n1426) );
  XOR U2365 ( .A(n2289), .B(n2341), .Z(n1430) );
  XNOR U2366 ( .A(n2201), .B(n2215), .Z(n2278) );
  XOR U2367 ( .A(n2220), .B(n2342), .Z(n2215) );
  XOR U2368 ( .A(key[251]), .B(\w0[1][123] ), .Z(n2342) );
  XOR U2369 ( .A(n2343), .B(n2344), .Z(\w0[1][123] ) );
  XOR U2370 ( .A(n1390), .B(n2033), .Z(n2344) );
  XOR U2371 ( .A(n2023), .B(n1419), .Z(n2033) );
  XOR U2372 ( .A(n1392), .B(n2312), .Z(n1419) );
  IV U2373 ( .A(n2247), .Z(n2023) );
  XOR U2374 ( .A(n2345), .B(n2346), .Z(n1390) );
  XOR U2375 ( .A(n2290), .B(n2347), .Z(n2346) );
  IV U2376 ( .A(n2348), .Z(n2290) );
  XNOR U2377 ( .A(n2289), .B(n2238), .Z(n2345) );
  XOR U2378 ( .A(n2350), .B(n2272), .Z(n2349) );
  NANDN U2379 ( .A(n2351), .B(n2352), .Z(n2272) );
  NOR U2380 ( .A(n2353), .B(n2354), .Z(n2350) );
  XOR U2381 ( .A(n807), .B(n804), .Z(n2343) );
  IV U2382 ( .A(n2006), .Z(n804) );
  XOR U2383 ( .A(n1391), .B(n1425), .Z(n2006) );
  XOR U2384 ( .A(n2356), .B(n2357), .Z(n1425) );
  XNOR U2385 ( .A(n2358), .B(n2359), .Z(n2357) );
  XNOR U2386 ( .A(n2276), .B(n2360), .Z(n2356) );
  XNOR U2387 ( .A(n2362), .B(n2321), .Z(n2361) );
  ANDN U2388 ( .B(n2363), .A(n2364), .Z(n2321) );
  ANDN U2389 ( .B(n2365), .A(n2366), .Z(n2362) );
  XOR U2390 ( .A(n2368), .B(n2369), .Z(n1391) );
  XNOR U2391 ( .A(n2370), .B(n2371), .Z(n2369) );
  XNOR U2392 ( .A(n2245), .B(n2309), .Z(n2368) );
  XNOR U2393 ( .A(n2373), .B(n2262), .Z(n2372) );
  ANDN U2394 ( .B(n2374), .A(n2375), .Z(n2262) );
  ANDN U2395 ( .B(n2376), .A(n2377), .Z(n2373) );
  XOR U2396 ( .A(n2334), .B(n2379), .Z(n2036) );
  XOR U2397 ( .A(n2334), .B(n814), .Z(n785) );
  XNOR U2398 ( .A(n2328), .B(n2380), .Z(n2334) );
  XNOR U2399 ( .A(n2381), .B(n2382), .Z(n2380) );
  NOR U2400 ( .A(n2383), .B(n2254), .Z(n2381) );
  XNOR U2401 ( .A(n2384), .B(n2385), .Z(n2328) );
  XNOR U2402 ( .A(n2386), .B(n2387), .Z(n2385) );
  NANDN U2403 ( .A(n2388), .B(n2389), .Z(n2387) );
  XOR U2404 ( .A(key[249]), .B(\w0[1][121] ), .Z(n2220) );
  XOR U2405 ( .A(n2390), .B(n2391), .Z(\w0[1][121] ) );
  XOR U2406 ( .A(n810), .B(n1434), .Z(n2391) );
  XNOR U2407 ( .A(n2239), .B(n2392), .Z(n1434) );
  XOR U2408 ( .A(n2289), .B(n2348), .Z(n2392) );
  XOR U2409 ( .A(n2355), .B(n2393), .Z(n2348) );
  XNOR U2410 ( .A(n2394), .B(n2395), .Z(n2393) );
  OR U2411 ( .A(n2287), .B(n2396), .Z(n2395) );
  XNOR U2412 ( .A(n2268), .B(n2397), .Z(n2355) );
  XNOR U2413 ( .A(n2398), .B(n2399), .Z(n2397) );
  OR U2414 ( .A(n2400), .B(n2401), .Z(n2399) );
  XNOR U2415 ( .A(n2402), .B(n2403), .Z(n2289) );
  XOR U2416 ( .A(n2404), .B(n2405), .Z(n2403) );
  OR U2417 ( .A(n2406), .B(n2275), .Z(n2405) );
  XNOR U2418 ( .A(n2341), .B(n2347), .Z(n2239) );
  XOR U2419 ( .A(n2268), .B(n2407), .Z(n2347) );
  XNOR U2420 ( .A(n2394), .B(n2408), .Z(n2407) );
  NANDN U2421 ( .A(n2409), .B(n2410), .Z(n2408) );
  OR U2422 ( .A(n2411), .B(n2412), .Z(n2394) );
  XOR U2423 ( .A(n2413), .B(n2398), .Z(n2268) );
  NANDN U2424 ( .A(n2414), .B(n2415), .Z(n2398) );
  AND U2425 ( .A(n2416), .B(n2417), .Z(n2413) );
  IV U2426 ( .A(n2418), .Z(n2341) );
  XNOR U2427 ( .A(n1429), .B(n1435), .Z(n810) );
  XNOR U2428 ( .A(n2246), .B(n2419), .Z(n1435) );
  XNOR U2429 ( .A(n2309), .B(n2370), .Z(n2419) );
  IV U2430 ( .A(n2300), .Z(n2370) );
  XOR U2431 ( .A(n2378), .B(n2420), .Z(n2300) );
  XNOR U2432 ( .A(n2421), .B(n2422), .Z(n2420) );
  NANDN U2433 ( .A(n2297), .B(n2423), .Z(n2422) );
  XNOR U2434 ( .A(n2260), .B(n2424), .Z(n2378) );
  XNOR U2435 ( .A(n2425), .B(n2426), .Z(n2424) );
  NANDN U2436 ( .A(n2427), .B(n2428), .Z(n2426) );
  XNOR U2437 ( .A(n2429), .B(n2430), .Z(n2309) );
  XNOR U2438 ( .A(n2431), .B(n2432), .Z(n2430) );
  NAND U2439 ( .A(n2433), .B(n2264), .Z(n2432) );
  XNOR U2440 ( .A(n2371), .B(n2308), .Z(n2246) );
  XNOR U2441 ( .A(n2260), .B(n2434), .Z(n2371) );
  XNOR U2442 ( .A(n2421), .B(n2435), .Z(n2434) );
  NANDN U2443 ( .A(n2436), .B(n2437), .Z(n2435) );
  OR U2444 ( .A(n2438), .B(n2439), .Z(n2421) );
  XOR U2445 ( .A(n2440), .B(n2425), .Z(n2260) );
  OR U2446 ( .A(n2441), .B(n2442), .Z(n2425) );
  ANDN U2447 ( .B(n2443), .A(n2444), .Z(n2440) );
  IV U2448 ( .A(n2445), .Z(n1429) );
  XOR U2449 ( .A(n2304), .B(n2446), .Z(n1392) );
  IV U2450 ( .A(n2360), .Z(n2304) );
  XOR U2451 ( .A(key[248]), .B(\w0[1][120] ), .Z(n2201) );
  XOR U2452 ( .A(n2447), .B(n2448), .Z(\w0[1][120] ) );
  XNOR U2453 ( .A(n2247), .B(n1414), .Z(n2448) );
  XOR U2454 ( .A(n1401), .B(n823), .Z(n1414) );
  XOR U2455 ( .A(n2308), .B(n2258), .Z(n823) );
  XOR U2456 ( .A(n2293), .B(n2449), .Z(n2258) );
  XOR U2457 ( .A(n2450), .B(n2431), .Z(n2449) );
  NANDN U2458 ( .A(n2451), .B(n2374), .Z(n2431) );
  XOR U2459 ( .A(n2376), .B(n2264), .Z(n2374) );
  ANDN U2460 ( .B(n2376), .A(n2452), .Z(n2450) );
  XNOR U2461 ( .A(n2429), .B(n2453), .Z(n2293) );
  XNOR U2462 ( .A(n2454), .B(n2455), .Z(n2453) );
  NANDN U2463 ( .A(n2427), .B(n2456), .Z(n2455) );
  XOR U2464 ( .A(n2429), .B(n2457), .Z(n2308) );
  XOR U2465 ( .A(n2458), .B(n2295), .Z(n2457) );
  OR U2466 ( .A(n2438), .B(n2459), .Z(n2295) );
  XOR U2467 ( .A(n2297), .B(n2460), .Z(n2438) );
  ANDN U2468 ( .B(n2461), .A(n2436), .Z(n2458) );
  XOR U2469 ( .A(n2462), .B(n2454), .Z(n2429) );
  NANDN U2470 ( .A(n2442), .B(n2463), .Z(n2454) );
  XOR U2471 ( .A(n2443), .B(n2427), .Z(n2442) );
  XNOR U2472 ( .A(n2460), .B(n2264), .Z(n2427) );
  XOR U2473 ( .A(n2464), .B(n2465), .Z(n2264) );
  NANDN U2474 ( .A(n2466), .B(n2467), .Z(n2465) );
  IV U2475 ( .A(n2436), .Z(n2460) );
  XNOR U2476 ( .A(n2468), .B(n2469), .Z(n2436) );
  NANDN U2477 ( .A(n2466), .B(n2470), .Z(n2469) );
  IV U2478 ( .A(n2471), .Z(n2443) );
  NOR U2479 ( .A(n2471), .B(n2472), .Z(n2462) );
  XOR U2480 ( .A(n2376), .B(n2297), .Z(n2471) );
  XOR U2481 ( .A(n2473), .B(n2468), .Z(n2297) );
  NANDN U2482 ( .A(n2474), .B(n2475), .Z(n2468) );
  NANDN U2483 ( .A(n2474), .B(n2479), .Z(n2464) );
  XOR U2484 ( .A(n2480), .B(n2481), .Z(n2466) );
  XOR U2485 ( .A(n2482), .B(n2477), .Z(n2481) );
  XNOR U2486 ( .A(n2483), .B(n2484), .Z(n2480) );
  XNOR U2487 ( .A(n2485), .B(n2486), .Z(n2484) );
  ANDN U2488 ( .B(n2482), .A(n2477), .Z(n2485) );
  ANDN U2489 ( .B(n2482), .A(n2476), .Z(n2478) );
  XNOR U2490 ( .A(n2483), .B(n2487), .Z(n2476) );
  XOR U2491 ( .A(n2488), .B(n2486), .Z(n2487) );
  NAND U2492 ( .A(n2475), .B(n2479), .Z(n2486) );
  XNOR U2493 ( .A(n2470), .B(n2477), .Z(n2475) );
  XOR U2494 ( .A(n2489), .B(n2490), .Z(n2477) );
  XNOR U2495 ( .A(n2491), .B(n2492), .Z(n2490) );
  XNOR U2496 ( .A(n2493), .B(n2494), .Z(n2489) );
  AND U2497 ( .A(n2467), .B(n2470), .Z(n2488) );
  XNOR U2498 ( .A(n2467), .B(n2470), .Z(n2483) );
  XNOR U2499 ( .A(n2495), .B(n2496), .Z(n2470) );
  XNOR U2500 ( .A(n2497), .B(n2498), .Z(n2496) );
  XNOR U2501 ( .A(n2491), .B(n2499), .Z(n2495) );
  XNOR U2502 ( .A(n2500), .B(n2494), .Z(n2499) );
  OR U2503 ( .A(n2375), .B(n2451), .Z(n2494) );
  XOR U2504 ( .A(n2452), .B(n2433), .Z(n2451) );
  XNOR U2505 ( .A(n2377), .B(n2265), .Z(n2375) );
  ANDN U2506 ( .B(n2433), .A(n2265), .Z(n2500) );
  XNOR U2507 ( .A(n2501), .B(n2502), .Z(n2467) );
  XNOR U2508 ( .A(n2503), .B(n2504), .Z(n2502) );
  XOR U2509 ( .A(n2423), .B(n2491), .Z(n2504) );
  XNOR U2510 ( .A(n2377), .B(n2452), .Z(n2491) );
  XNOR U2511 ( .A(n2298), .B(n2505), .Z(n2501) );
  XNOR U2512 ( .A(n2506), .B(n2507), .Z(n2505) );
  ANDN U2513 ( .B(n2437), .A(n2508), .Z(n2506) );
  XNOR U2514 ( .A(n2509), .B(n2510), .Z(n2482) );
  XNOR U2515 ( .A(n2492), .B(n2511), .Z(n2510) );
  XOR U2516 ( .A(n2508), .B(n2498), .Z(n2511) );
  XOR U2517 ( .A(n2512), .B(n2433), .Z(n2498) );
  XNOR U2518 ( .A(n2503), .B(n2513), .Z(n2492) );
  XNOR U2519 ( .A(n2514), .B(n2515), .Z(n2513) );
  NAND U2520 ( .A(n2456), .B(n2428), .Z(n2515) );
  IV U2521 ( .A(n2497), .Z(n2503) );
  XNOR U2522 ( .A(n2516), .B(n2514), .Z(n2497) );
  NANDN U2523 ( .A(n2441), .B(n2463), .Z(n2514) );
  XNOR U2524 ( .A(n2472), .B(n2456), .Z(n2463) );
  XOR U2525 ( .A(n2461), .B(n2433), .Z(n2456) );
  XOR U2526 ( .A(n2517), .B(n2518), .Z(n2433) );
  XOR U2527 ( .A(n2444), .B(n2428), .Z(n2441) );
  XOR U2528 ( .A(n2512), .B(n2437), .Z(n2428) );
  IV U2529 ( .A(n2265), .Z(n2512) );
  XNOR U2530 ( .A(n2519), .B(n2520), .Z(n2265) );
  NOR U2531 ( .A(n2444), .B(n2472), .Z(n2516) );
  XOR U2532 ( .A(n2521), .B(n2452), .Z(n2472) );
  XOR U2533 ( .A(n2522), .B(n2523), .Z(n2452) );
  XOR U2534 ( .A(n2524), .B(n2525), .Z(n2523) );
  XOR U2535 ( .A(n2377), .B(n2423), .Z(n2444) );
  XOR U2536 ( .A(n2437), .B(n2526), .Z(n2509) );
  XNOR U2537 ( .A(n2527), .B(n2507), .Z(n2526) );
  OR U2538 ( .A(n2439), .B(n2459), .Z(n2507) );
  XOR U2539 ( .A(n2298), .B(n2461), .Z(n2459) );
  IV U2540 ( .A(n2508), .Z(n2461) );
  XOR U2541 ( .A(n2528), .B(n2529), .Z(n2508) );
  XOR U2542 ( .A(n2530), .B(n2522), .Z(n2529) );
  XOR U2543 ( .A(n2519), .B(n2531), .Z(n2522) );
  XNOR U2544 ( .A(state[43]), .B(key[43]), .Z(n2531) );
  XOR U2545 ( .A(n2532), .B(n2298), .Z(n2528) );
  XNOR U2546 ( .A(n2423), .B(n2437), .Z(n2439) );
  ANDN U2547 ( .B(n2423), .A(n2298), .Z(n2527) );
  IV U2548 ( .A(n2521), .Z(n2298) );
  XOR U2549 ( .A(n2530), .B(n2520), .Z(n2423) );
  XNOR U2550 ( .A(state[44]), .B(key[44]), .Z(n2530) );
  XNOR U2551 ( .A(n2525), .B(n2533), .Z(n2437) );
  XNOR U2552 ( .A(n2377), .B(n2519), .Z(n2533) );
  XNOR U2553 ( .A(state[41]), .B(key[41]), .Z(n2519) );
  XOR U2554 ( .A(n2518), .B(n2534), .Z(n2377) );
  XOR U2555 ( .A(n2532), .B(n2517), .Z(n2534) );
  XOR U2556 ( .A(state[45]), .B(key[45]), .Z(n2517) );
  XNOR U2557 ( .A(state[47]), .B(key[47]), .Z(n2532) );
  IV U2558 ( .A(n2524), .Z(n2518) );
  XOR U2559 ( .A(n2521), .B(n2535), .Z(n2524) );
  XNOR U2560 ( .A(state[46]), .B(key[46]), .Z(n2535) );
  XOR U2561 ( .A(state[40]), .B(key[40]), .Z(n2521) );
  XOR U2562 ( .A(state[42]), .B(key[42]), .Z(n2525) );
  XOR U2563 ( .A(n2270), .B(n2418), .Z(n1401) );
  XOR U2564 ( .A(n2402), .B(n2536), .Z(n2418) );
  XOR U2565 ( .A(n2537), .B(n2285), .Z(n2536) );
  OR U2566 ( .A(n2538), .B(n2411), .Z(n2285) );
  XOR U2567 ( .A(n2287), .B(n2539), .Z(n2411) );
  ANDN U2568 ( .B(n2540), .A(n2409), .Z(n2537) );
  XNOR U2569 ( .A(n2283), .B(n2541), .Z(n2270) );
  XNOR U2570 ( .A(n2542), .B(n2404), .Z(n2541) );
  ANDN U2571 ( .B(n2352), .A(n2543), .Z(n2404) );
  XOR U2572 ( .A(n2354), .B(n2275), .Z(n2352) );
  NOR U2573 ( .A(n2544), .B(n2354), .Z(n2542) );
  XNOR U2574 ( .A(n2402), .B(n2545), .Z(n2283) );
  XNOR U2575 ( .A(n2546), .B(n2547), .Z(n2545) );
  NANDN U2576 ( .A(n2400), .B(n2548), .Z(n2547) );
  XOR U2577 ( .A(n2549), .B(n2546), .Z(n2402) );
  OR U2578 ( .A(n2414), .B(n2550), .Z(n2546) );
  XOR U2579 ( .A(n2416), .B(n2400), .Z(n2414) );
  XOR U2580 ( .A(n2539), .B(n2275), .Z(n2400) );
  XNOR U2581 ( .A(n2551), .B(n2552), .Z(n2275) );
  NANDN U2582 ( .A(n2553), .B(n2554), .Z(n2552) );
  IV U2583 ( .A(n2409), .Z(n2539) );
  XNOR U2584 ( .A(n2555), .B(n2556), .Z(n2409) );
  NANDN U2585 ( .A(n2553), .B(n2557), .Z(n2556) );
  ANDN U2586 ( .B(n2416), .A(n2558), .Z(n2549) );
  XOR U2587 ( .A(n2354), .B(n2287), .Z(n2416) );
  XOR U2588 ( .A(n2559), .B(n2555), .Z(n2287) );
  NANDN U2589 ( .A(n2560), .B(n2561), .Z(n2555) );
  NANDN U2590 ( .A(n2560), .B(n2565), .Z(n2551) );
  XOR U2591 ( .A(n2566), .B(n2567), .Z(n2553) );
  XOR U2592 ( .A(n2568), .B(n2563), .Z(n2567) );
  XNOR U2593 ( .A(n2569), .B(n2570), .Z(n2566) );
  XNOR U2594 ( .A(n2571), .B(n2572), .Z(n2570) );
  ANDN U2595 ( .B(n2568), .A(n2563), .Z(n2571) );
  ANDN U2596 ( .B(n2568), .A(n2562), .Z(n2564) );
  XNOR U2597 ( .A(n2569), .B(n2573), .Z(n2562) );
  XOR U2598 ( .A(n2574), .B(n2572), .Z(n2573) );
  NAND U2599 ( .A(n2561), .B(n2565), .Z(n2572) );
  XNOR U2600 ( .A(n2557), .B(n2563), .Z(n2561) );
  XOR U2601 ( .A(n2575), .B(n2576), .Z(n2563) );
  XOR U2602 ( .A(n2577), .B(n2578), .Z(n2576) );
  XNOR U2603 ( .A(n2579), .B(n2580), .Z(n2575) );
  ANDN U2604 ( .B(n2581), .A(n2353), .Z(n2579) );
  AND U2605 ( .A(n2554), .B(n2557), .Z(n2574) );
  XNOR U2606 ( .A(n2554), .B(n2557), .Z(n2569) );
  XNOR U2607 ( .A(n2582), .B(n2583), .Z(n2557) );
  XNOR U2608 ( .A(n2584), .B(n2585), .Z(n2583) );
  XOR U2609 ( .A(n2577), .B(n2586), .Z(n2582) );
  XNOR U2610 ( .A(n2587), .B(n2580), .Z(n2586) );
  OR U2611 ( .A(n2351), .B(n2543), .Z(n2580) );
  XNOR U2612 ( .A(n2544), .B(n2406), .Z(n2543) );
  XNOR U2613 ( .A(n2353), .B(n2588), .Z(n2351) );
  NOR U2614 ( .A(n2588), .B(n2406), .Z(n2587) );
  XNOR U2615 ( .A(n2589), .B(n2590), .Z(n2554) );
  XNOR U2616 ( .A(n2591), .B(n2592), .Z(n2590) );
  XOR U2617 ( .A(n2396), .B(n2577), .Z(n2592) );
  XOR U2618 ( .A(n2581), .B(n2593), .Z(n2577) );
  XNOR U2619 ( .A(n2288), .B(n2594), .Z(n2589) );
  XNOR U2620 ( .A(n2595), .B(n2596), .Z(n2594) );
  ANDN U2621 ( .B(n2410), .A(n2597), .Z(n2595) );
  XNOR U2622 ( .A(n2598), .B(n2599), .Z(n2568) );
  XNOR U2623 ( .A(n2578), .B(n2600), .Z(n2599) );
  XNOR U2624 ( .A(n2410), .B(n2585), .Z(n2600) );
  XOR U2625 ( .A(n2406), .B(n2588), .Z(n2585) );
  XNOR U2626 ( .A(n2591), .B(n2601), .Z(n2578) );
  XNOR U2627 ( .A(n2602), .B(n2603), .Z(n2601) );
  NANDN U2628 ( .A(n2401), .B(n2548), .Z(n2603) );
  IV U2629 ( .A(n2584), .Z(n2591) );
  XNOR U2630 ( .A(n2604), .B(n2602), .Z(n2584) );
  NANDN U2631 ( .A(n2550), .B(n2415), .Z(n2602) );
  XOR U2632 ( .A(n2410), .B(n2588), .Z(n2401) );
  IV U2633 ( .A(n2274), .Z(n2588) );
  XOR U2634 ( .A(n2605), .B(n2606), .Z(n2274) );
  XNOR U2635 ( .A(n2607), .B(n2608), .Z(n2606) );
  XOR U2636 ( .A(n2558), .B(n2548), .Z(n2550) );
  XNOR U2637 ( .A(n2540), .B(n2406), .Z(n2548) );
  XNOR U2638 ( .A(n2608), .B(n2605), .Z(n2406) );
  ANDN U2639 ( .B(n2417), .A(n2558), .Z(n2604) );
  XNOR U2640 ( .A(n2609), .B(n2581), .Z(n2558) );
  IV U2641 ( .A(n2544), .Z(n2581) );
  XNOR U2642 ( .A(n2610), .B(n2611), .Z(n2544) );
  XNOR U2643 ( .A(n2612), .B(n2608), .Z(n2611) );
  XOR U2644 ( .A(n2613), .B(n2593), .Z(n2417) );
  XNOR U2645 ( .A(n2597), .B(n2614), .Z(n2598) );
  XNOR U2646 ( .A(n2615), .B(n2596), .Z(n2614) );
  OR U2647 ( .A(n2412), .B(n2538), .Z(n2596) );
  XOR U2648 ( .A(n2288), .B(n2540), .Z(n2538) );
  IV U2649 ( .A(n2597), .Z(n2540) );
  XOR U2650 ( .A(n2396), .B(n2410), .Z(n2412) );
  XNOR U2651 ( .A(n2593), .B(n2616), .Z(n2410) );
  XNOR U2652 ( .A(n2607), .B(n2610), .Z(n2616) );
  XNOR U2653 ( .A(state[2]), .B(key[2]), .Z(n2610) );
  IV U2654 ( .A(n2353), .Z(n2593) );
  XOR U2655 ( .A(n2617), .B(n2618), .Z(n2353) );
  XOR U2656 ( .A(n2608), .B(n2619), .Z(n2618) );
  IV U2657 ( .A(n2613), .Z(n2396) );
  ANDN U2658 ( .B(n2613), .A(n2288), .Z(n2615) );
  XOR U2659 ( .A(n2605), .B(n2620), .Z(n2613) );
  XNOR U2660 ( .A(n2608), .B(n2621), .Z(n2620) );
  XOR U2661 ( .A(n2609), .B(n2622), .Z(n2608) );
  XNOR U2662 ( .A(state[6]), .B(key[6]), .Z(n2622) );
  IV U2663 ( .A(n2617), .Z(n2605) );
  XOR U2664 ( .A(state[5]), .B(key[5]), .Z(n2617) );
  XOR U2665 ( .A(n2623), .B(n2624), .Z(n2597) );
  XOR U2666 ( .A(n2621), .B(n2619), .Z(n2624) );
  XOR U2667 ( .A(state[7]), .B(key[7]), .Z(n2619) );
  XNOR U2668 ( .A(state[4]), .B(key[4]), .Z(n2621) );
  XOR U2669 ( .A(n2288), .B(n2612), .Z(n2623) );
  XNOR U2670 ( .A(n2607), .B(n2625), .Z(n2612) );
  XNOR U2671 ( .A(state[3]), .B(key[3]), .Z(n2625) );
  XNOR U2672 ( .A(state[1]), .B(key[1]), .Z(n2607) );
  IV U2673 ( .A(n2609), .Z(n2288) );
  XOR U2674 ( .A(state[0]), .B(key[0]), .Z(n2609) );
  XNOR U2675 ( .A(n2446), .B(n2312), .Z(n2247) );
  XOR U2676 ( .A(n2313), .B(n2626), .Z(n2312) );
  XOR U2677 ( .A(n2627), .B(n2628), .Z(n2626) );
  ANDN U2678 ( .B(n2365), .A(n2629), .Z(n2627) );
  XNOR U2679 ( .A(n2630), .B(n2631), .Z(n2313) );
  XNOR U2680 ( .A(n2632), .B(n2633), .Z(n2631) );
  NANDN U2681 ( .A(n2634), .B(n2635), .Z(n2633) );
  XOR U2682 ( .A(n2445), .B(n808), .Z(n2447) );
  XNOR U2683 ( .A(n2242), .B(n2636), .Z(n808) );
  XOR U2684 ( .A(n2230), .B(n2244), .Z(n2636) );
  XOR U2685 ( .A(n2255), .B(n2637), .Z(n2244) );
  XNOR U2686 ( .A(n2638), .B(n2639), .Z(n2637) );
  OR U2687 ( .A(n2332), .B(n2640), .Z(n2639) );
  XNOR U2688 ( .A(n2327), .B(n2641), .Z(n2255) );
  XNOR U2689 ( .A(n2642), .B(n2643), .Z(n2641) );
  OR U2690 ( .A(n2388), .B(n2644), .Z(n2643) );
  XNOR U2691 ( .A(n2384), .B(n2645), .Z(n2230) );
  XOR U2692 ( .A(n2382), .B(n2646), .Z(n2645) );
  OR U2693 ( .A(n2647), .B(n2338), .Z(n2646) );
  ANDN U2694 ( .B(n2340), .A(n2648), .Z(n2382) );
  XOR U2695 ( .A(n2254), .B(n2338), .Z(n2340) );
  XNOR U2696 ( .A(n2379), .B(n2229), .Z(n2242) );
  XOR U2697 ( .A(n2327), .B(n2649), .Z(n2229) );
  XNOR U2698 ( .A(n2638), .B(n2650), .Z(n2649) );
  NANDN U2699 ( .A(n2651), .B(n2652), .Z(n2650) );
  OR U2700 ( .A(n2653), .B(n2654), .Z(n2638) );
  XOR U2701 ( .A(n2655), .B(n2642), .Z(n2327) );
  NANDN U2702 ( .A(n2656), .B(n2657), .Z(n2642) );
  AND U2703 ( .A(n2658), .B(n2659), .Z(n2655) );
  XOR U2704 ( .A(n2384), .B(n2660), .Z(n2379) );
  XOR U2705 ( .A(n2661), .B(n2330), .Z(n2660) );
  OR U2706 ( .A(n2662), .B(n2653), .Z(n2330) );
  XOR U2707 ( .A(n2332), .B(n2663), .Z(n2653) );
  ANDN U2708 ( .B(n2664), .A(n2651), .Z(n2661) );
  XOR U2709 ( .A(n2665), .B(n2386), .Z(n2384) );
  OR U2710 ( .A(n2656), .B(n2666), .Z(n2386) );
  XOR U2711 ( .A(n2658), .B(n2388), .Z(n2656) );
  XOR U2712 ( .A(n2663), .B(n2338), .Z(n2388) );
  XNOR U2713 ( .A(n2667), .B(n2668), .Z(n2338) );
  NANDN U2714 ( .A(n2669), .B(n2670), .Z(n2668) );
  IV U2715 ( .A(n2651), .Z(n2663) );
  XNOR U2716 ( .A(n2671), .B(n2672), .Z(n2651) );
  NANDN U2717 ( .A(n2669), .B(n2673), .Z(n2672) );
  ANDN U2718 ( .B(n2658), .A(n2674), .Z(n2665) );
  XOR U2719 ( .A(n2254), .B(n2332), .Z(n2658) );
  XOR U2720 ( .A(n2675), .B(n2671), .Z(n2332) );
  NANDN U2721 ( .A(n2676), .B(n2677), .Z(n2671) );
  NANDN U2722 ( .A(n2676), .B(n2681), .Z(n2667) );
  XOR U2723 ( .A(n2682), .B(n2683), .Z(n2669) );
  XOR U2724 ( .A(n2684), .B(n2679), .Z(n2683) );
  XNOR U2725 ( .A(n2685), .B(n2686), .Z(n2682) );
  XNOR U2726 ( .A(n2687), .B(n2688), .Z(n2686) );
  ANDN U2727 ( .B(n2684), .A(n2679), .Z(n2687) );
  ANDN U2728 ( .B(n2684), .A(n2678), .Z(n2680) );
  XNOR U2729 ( .A(n2685), .B(n2689), .Z(n2678) );
  XOR U2730 ( .A(n2690), .B(n2688), .Z(n2689) );
  NAND U2731 ( .A(n2677), .B(n2681), .Z(n2688) );
  XNOR U2732 ( .A(n2673), .B(n2679), .Z(n2677) );
  XOR U2733 ( .A(n2691), .B(n2692), .Z(n2679) );
  XOR U2734 ( .A(n2693), .B(n2694), .Z(n2692) );
  XNOR U2735 ( .A(n2695), .B(n2696), .Z(n2691) );
  ANDN U2736 ( .B(n2697), .A(n2253), .Z(n2695) );
  AND U2737 ( .A(n2670), .B(n2673), .Z(n2690) );
  XNOR U2738 ( .A(n2670), .B(n2673), .Z(n2685) );
  XNOR U2739 ( .A(n2698), .B(n2699), .Z(n2673) );
  XNOR U2740 ( .A(n2700), .B(n2701), .Z(n2699) );
  XOR U2741 ( .A(n2693), .B(n2702), .Z(n2698) );
  XNOR U2742 ( .A(n2703), .B(n2696), .Z(n2702) );
  OR U2743 ( .A(n2339), .B(n2648), .Z(n2696) );
  XNOR U2744 ( .A(n2383), .B(n2647), .Z(n2648) );
  XNOR U2745 ( .A(n2253), .B(n2704), .Z(n2339) );
  NOR U2746 ( .A(n2704), .B(n2647), .Z(n2703) );
  XNOR U2747 ( .A(n2705), .B(n2706), .Z(n2670) );
  XNOR U2748 ( .A(n2707), .B(n2708), .Z(n2706) );
  XOR U2749 ( .A(n2640), .B(n2693), .Z(n2708) );
  XOR U2750 ( .A(n2697), .B(n2709), .Z(n2693) );
  XNOR U2751 ( .A(n2333), .B(n2710), .Z(n2705) );
  XNOR U2752 ( .A(n2711), .B(n2712), .Z(n2710) );
  ANDN U2753 ( .B(n2652), .A(n2713), .Z(n2711) );
  XNOR U2754 ( .A(n2714), .B(n2715), .Z(n2684) );
  XNOR U2755 ( .A(n2694), .B(n2716), .Z(n2715) );
  XNOR U2756 ( .A(n2652), .B(n2701), .Z(n2716) );
  XOR U2757 ( .A(n2647), .B(n2704), .Z(n2701) );
  XNOR U2758 ( .A(n2707), .B(n2717), .Z(n2694) );
  XNOR U2759 ( .A(n2718), .B(n2719), .Z(n2717) );
  NANDN U2760 ( .A(n2644), .B(n2389), .Z(n2719) );
  IV U2761 ( .A(n2700), .Z(n2707) );
  XNOR U2762 ( .A(n2720), .B(n2718), .Z(n2700) );
  NANDN U2763 ( .A(n2666), .B(n2657), .Z(n2718) );
  XOR U2764 ( .A(n2652), .B(n2704), .Z(n2644) );
  IV U2765 ( .A(n2337), .Z(n2704) );
  XOR U2766 ( .A(n2721), .B(n2722), .Z(n2337) );
  XNOR U2767 ( .A(n2723), .B(n2724), .Z(n2722) );
  XOR U2768 ( .A(n2674), .B(n2389), .Z(n2666) );
  XNOR U2769 ( .A(n2664), .B(n2647), .Z(n2389) );
  XNOR U2770 ( .A(n2724), .B(n2721), .Z(n2647) );
  ANDN U2771 ( .B(n2659), .A(n2674), .Z(n2720) );
  XNOR U2772 ( .A(n2725), .B(n2697), .Z(n2674) );
  IV U2773 ( .A(n2383), .Z(n2697) );
  XNOR U2774 ( .A(n2726), .B(n2727), .Z(n2383) );
  XNOR U2775 ( .A(n2728), .B(n2724), .Z(n2727) );
  XOR U2776 ( .A(n2729), .B(n2709), .Z(n2659) );
  XNOR U2777 ( .A(n2713), .B(n2730), .Z(n2714) );
  XNOR U2778 ( .A(n2731), .B(n2712), .Z(n2730) );
  OR U2779 ( .A(n2654), .B(n2662), .Z(n2712) );
  XOR U2780 ( .A(n2333), .B(n2664), .Z(n2662) );
  IV U2781 ( .A(n2713), .Z(n2664) );
  XOR U2782 ( .A(n2640), .B(n2652), .Z(n2654) );
  XNOR U2783 ( .A(n2709), .B(n2732), .Z(n2652) );
  XNOR U2784 ( .A(n2723), .B(n2726), .Z(n2732) );
  XNOR U2785 ( .A(state[122]), .B(key[122]), .Z(n2726) );
  IV U2786 ( .A(n2253), .Z(n2709) );
  XOR U2787 ( .A(n2733), .B(n2734), .Z(n2253) );
  XOR U2788 ( .A(n2724), .B(n2735), .Z(n2734) );
  IV U2789 ( .A(n2729), .Z(n2640) );
  ANDN U2790 ( .B(n2729), .A(n2333), .Z(n2731) );
  XOR U2791 ( .A(n2721), .B(n2736), .Z(n2729) );
  XNOR U2792 ( .A(n2724), .B(n2737), .Z(n2736) );
  XOR U2793 ( .A(n2725), .B(n2738), .Z(n2724) );
  XNOR U2794 ( .A(state[126]), .B(key[126]), .Z(n2738) );
  IV U2795 ( .A(n2733), .Z(n2721) );
  XOR U2796 ( .A(state[125]), .B(key[125]), .Z(n2733) );
  XOR U2797 ( .A(n2739), .B(n2740), .Z(n2713) );
  XOR U2798 ( .A(n2737), .B(n2735), .Z(n2740) );
  XOR U2799 ( .A(state[127]), .B(key[127]), .Z(n2735) );
  XNOR U2800 ( .A(state[124]), .B(key[124]), .Z(n2737) );
  XOR U2801 ( .A(n2333), .B(n2728), .Z(n2739) );
  XNOR U2802 ( .A(n2723), .B(n2741), .Z(n2728) );
  XNOR U2803 ( .A(state[123]), .B(key[123]), .Z(n2741) );
  XNOR U2804 ( .A(state[121]), .B(key[121]), .Z(n2723) );
  IV U2805 ( .A(n2725), .Z(n2333) );
  XOR U2806 ( .A(state[120]), .B(key[120]), .Z(n2725) );
  XNOR U2807 ( .A(n2360), .B(n2358), .Z(n2742) );
  IV U2808 ( .A(n2305), .Z(n2358) );
  XOR U2809 ( .A(n2367), .B(n2743), .Z(n2305) );
  XNOR U2810 ( .A(n2744), .B(n2745), .Z(n2743) );
  NANDN U2811 ( .A(n2317), .B(n2746), .Z(n2745) );
  XNOR U2812 ( .A(n2319), .B(n2747), .Z(n2367) );
  XNOR U2813 ( .A(n2748), .B(n2749), .Z(n2747) );
  NANDN U2814 ( .A(n2634), .B(n2750), .Z(n2749) );
  XNOR U2815 ( .A(n2630), .B(n2751), .Z(n2360) );
  XNOR U2816 ( .A(n2628), .B(n2752), .Z(n2751) );
  NAND U2817 ( .A(n2753), .B(n2323), .Z(n2752) );
  NANDN U2818 ( .A(n2754), .B(n2363), .Z(n2628) );
  XOR U2819 ( .A(n2365), .B(n2323), .Z(n2363) );
  XOR U2820 ( .A(n2359), .B(n2446), .Z(n2277) );
  XOR U2821 ( .A(n2630), .B(n2755), .Z(n2446) );
  XOR U2822 ( .A(n2756), .B(n2315), .Z(n2755) );
  OR U2823 ( .A(n2757), .B(n2758), .Z(n2315) );
  ANDN U2824 ( .B(n2759), .A(n2760), .Z(n2756) );
  XOR U2825 ( .A(n2761), .B(n2632), .Z(n2630) );
  NANDN U2826 ( .A(n2762), .B(n2763), .Z(n2632) );
  NOR U2827 ( .A(n2764), .B(n2765), .Z(n2761) );
  XNOR U2828 ( .A(n2319), .B(n2766), .Z(n2359) );
  XNOR U2829 ( .A(n2744), .B(n2767), .Z(n2766) );
  NANDN U2830 ( .A(n2760), .B(n2768), .Z(n2767) );
  OR U2831 ( .A(n2757), .B(n2769), .Z(n2744) );
  XOR U2832 ( .A(n2317), .B(n2770), .Z(n2757) );
  XOR U2833 ( .A(n2771), .B(n2748), .Z(n2319) );
  OR U2834 ( .A(n2772), .B(n2762), .Z(n2748) );
  XOR U2835 ( .A(n2773), .B(n2634), .Z(n2762) );
  XNOR U2836 ( .A(n2770), .B(n2323), .Z(n2634) );
  XOR U2837 ( .A(n2774), .B(n2775), .Z(n2323) );
  NANDN U2838 ( .A(n2776), .B(n2777), .Z(n2775) );
  IV U2839 ( .A(n2760), .Z(n2770) );
  XNOR U2840 ( .A(n2778), .B(n2779), .Z(n2760) );
  NANDN U2841 ( .A(n2776), .B(n2780), .Z(n2779) );
  ANDN U2842 ( .B(n2773), .A(n2781), .Z(n2771) );
  IV U2843 ( .A(n2764), .Z(n2773) );
  XOR U2844 ( .A(n2365), .B(n2317), .Z(n2764) );
  XOR U2845 ( .A(n2782), .B(n2778), .Z(n2317) );
  NANDN U2846 ( .A(n2783), .B(n2784), .Z(n2778) );
  NANDN U2847 ( .A(n2783), .B(n2788), .Z(n2774) );
  XOR U2848 ( .A(n2789), .B(n2790), .Z(n2776) );
  XOR U2849 ( .A(n2791), .B(n2786), .Z(n2790) );
  XNOR U2850 ( .A(n2792), .B(n2793), .Z(n2789) );
  XNOR U2851 ( .A(n2794), .B(n2795), .Z(n2793) );
  ANDN U2852 ( .B(n2791), .A(n2786), .Z(n2794) );
  ANDN U2853 ( .B(n2791), .A(n2785), .Z(n2787) );
  XNOR U2854 ( .A(n2792), .B(n2796), .Z(n2785) );
  XOR U2855 ( .A(n2797), .B(n2795), .Z(n2796) );
  NAND U2856 ( .A(n2784), .B(n2788), .Z(n2795) );
  XNOR U2857 ( .A(n2780), .B(n2786), .Z(n2784) );
  XOR U2858 ( .A(n2798), .B(n2799), .Z(n2786) );
  XNOR U2859 ( .A(n2800), .B(n2801), .Z(n2799) );
  XNOR U2860 ( .A(n2802), .B(n2803), .Z(n2798) );
  AND U2861 ( .A(n2777), .B(n2780), .Z(n2797) );
  XNOR U2862 ( .A(n2777), .B(n2780), .Z(n2792) );
  XNOR U2863 ( .A(n2804), .B(n2805), .Z(n2780) );
  XNOR U2864 ( .A(n2806), .B(n2807), .Z(n2805) );
  XNOR U2865 ( .A(n2800), .B(n2808), .Z(n2804) );
  XNOR U2866 ( .A(n2809), .B(n2803), .Z(n2808) );
  OR U2867 ( .A(n2364), .B(n2754), .Z(n2803) );
  XOR U2868 ( .A(n2629), .B(n2753), .Z(n2754) );
  XNOR U2869 ( .A(n2366), .B(n2324), .Z(n2364) );
  ANDN U2870 ( .B(n2753), .A(n2324), .Z(n2809) );
  XNOR U2871 ( .A(n2810), .B(n2811), .Z(n2777) );
  XNOR U2872 ( .A(n2812), .B(n2813), .Z(n2811) );
  XOR U2873 ( .A(n2746), .B(n2800), .Z(n2813) );
  XNOR U2874 ( .A(n2366), .B(n2629), .Z(n2800) );
  XNOR U2875 ( .A(n2318), .B(n2814), .Z(n2810) );
  XNOR U2876 ( .A(n2815), .B(n2816), .Z(n2814) );
  ANDN U2877 ( .B(n2768), .A(n2817), .Z(n2815) );
  XNOR U2878 ( .A(n2818), .B(n2819), .Z(n2791) );
  XNOR U2879 ( .A(n2801), .B(n2820), .Z(n2819) );
  XOR U2880 ( .A(n2817), .B(n2807), .Z(n2820) );
  XOR U2881 ( .A(n2821), .B(n2753), .Z(n2807) );
  XNOR U2882 ( .A(n2812), .B(n2822), .Z(n2801) );
  XNOR U2883 ( .A(n2823), .B(n2824), .Z(n2822) );
  NAND U2884 ( .A(n2635), .B(n2750), .Z(n2824) );
  IV U2885 ( .A(n2806), .Z(n2812) );
  XNOR U2886 ( .A(n2825), .B(n2823), .Z(n2806) );
  NANDN U2887 ( .A(n2772), .B(n2763), .Z(n2823) );
  XNOR U2888 ( .A(n2765), .B(n2635), .Z(n2763) );
  XOR U2889 ( .A(n2759), .B(n2753), .Z(n2635) );
  XOR U2890 ( .A(n2826), .B(n2827), .Z(n2753) );
  XOR U2891 ( .A(n2781), .B(n2750), .Z(n2772) );
  XOR U2892 ( .A(n2821), .B(n2768), .Z(n2750) );
  IV U2893 ( .A(n2324), .Z(n2821) );
  XNOR U2894 ( .A(n2828), .B(n2829), .Z(n2324) );
  NOR U2895 ( .A(n2781), .B(n2765), .Z(n2825) );
  XOR U2896 ( .A(n2830), .B(n2629), .Z(n2765) );
  XOR U2897 ( .A(n2831), .B(n2832), .Z(n2629) );
  XOR U2898 ( .A(n2833), .B(n2834), .Z(n2832) );
  XOR U2899 ( .A(n2366), .B(n2746), .Z(n2781) );
  XOR U2900 ( .A(n2768), .B(n2835), .Z(n2818) );
  XNOR U2901 ( .A(n2836), .B(n2816), .Z(n2835) );
  OR U2902 ( .A(n2769), .B(n2758), .Z(n2816) );
  XOR U2903 ( .A(n2318), .B(n2759), .Z(n2758) );
  IV U2904 ( .A(n2817), .Z(n2759) );
  XOR U2905 ( .A(n2837), .B(n2838), .Z(n2817) );
  XOR U2906 ( .A(n2839), .B(n2831), .Z(n2838) );
  XOR U2907 ( .A(n2828), .B(n2840), .Z(n2831) );
  XNOR U2908 ( .A(state[83]), .B(key[83]), .Z(n2840) );
  XOR U2909 ( .A(n2841), .B(n2318), .Z(n2837) );
  XNOR U2910 ( .A(n2746), .B(n2768), .Z(n2769) );
  ANDN U2911 ( .B(n2746), .A(n2318), .Z(n2836) );
  IV U2912 ( .A(n2830), .Z(n2318) );
  XOR U2913 ( .A(n2839), .B(n2829), .Z(n2746) );
  XNOR U2914 ( .A(state[84]), .B(key[84]), .Z(n2839) );
  XNOR U2915 ( .A(n2834), .B(n2842), .Z(n2768) );
  XNOR U2916 ( .A(n2366), .B(n2828), .Z(n2842) );
  XNOR U2917 ( .A(state[81]), .B(key[81]), .Z(n2828) );
  XOR U2918 ( .A(n2827), .B(n2843), .Z(n2366) );
  XOR U2919 ( .A(n2841), .B(n2826), .Z(n2843) );
  XOR U2920 ( .A(state[85]), .B(key[85]), .Z(n2826) );
  XNOR U2921 ( .A(state[87]), .B(key[87]), .Z(n2841) );
  IV U2922 ( .A(n2833), .Z(n2827) );
  XOR U2923 ( .A(n2830), .B(n2844), .Z(n2833) );
  XNOR U2924 ( .A(state[86]), .B(key[86]), .Z(n2844) );
  XOR U2925 ( .A(state[80]), .B(key[80]), .Z(n2830) );
  XOR U2926 ( .A(state[82]), .B(key[82]), .Z(n2834) );
  XOR U2927 ( .A(n2845), .B(n2846), .Z(out[11]) );
  XNOR U2928 ( .A(n4), .B(n2041), .Z(n2846) );
  XNOR U2929 ( .A(n2847), .B(n2848), .Z(n2041) );
  XNOR U2930 ( .A(n2849), .B(n2057), .Z(n2848) );
  ANDN U2931 ( .B(n2850), .A(n2851), .Z(n2057) );
  NOR U2932 ( .A(n2066), .B(n2852), .Z(n2849) );
  XNOR U2933 ( .A(n2043), .B(n2853), .Z(n2845) );
  XOR U2934 ( .A(key[139]), .B(n5), .Z(n2853) );
  XOR U2935 ( .A(n2847), .B(n2854), .Z(n5) );
  XNOR U2936 ( .A(n2855), .B(n2856), .Z(n2854) );
  NANDN U2937 ( .A(n2053), .B(n2857), .Z(n2856) );
  XNOR U2938 ( .A(n2048), .B(n2858), .Z(n2847) );
  XNOR U2939 ( .A(n2859), .B(n2860), .Z(n2858) );
  NAND U2940 ( .A(n2861), .B(n2071), .Z(n2860) );
  XNOR U2941 ( .A(n2048), .B(n2862), .Z(n2043) );
  XNOR U2942 ( .A(n2855), .B(n2863), .Z(n2862) );
  NANDN U2943 ( .A(n2864), .B(n2865), .Z(n2863) );
  OR U2944 ( .A(n2866), .B(n2867), .Z(n2855) );
  XOR U2945 ( .A(n2868), .B(n2859), .Z(n2048) );
  OR U2946 ( .A(n2869), .B(n2870), .Z(n2859) );
  ANDN U2947 ( .B(n2871), .A(n2872), .Z(n2868) );
  XOR U2948 ( .A(n2873), .B(n2874), .Z(out[119]) );
  XOR U2949 ( .A(n2875), .B(n2876), .Z(n2873) );
  XOR U2950 ( .A(key[247]), .B(n2877), .Z(n2876) );
  XNOR U2951 ( .A(n2878), .B(n2879), .Z(out[118]) );
  XNOR U2952 ( .A(key[246]), .B(n2880), .Z(n2879) );
  XOR U2953 ( .A(n2881), .B(n2882), .Z(out[117]) );
  XNOR U2954 ( .A(n2883), .B(n2884), .Z(n2882) );
  XOR U2955 ( .A(n2875), .B(n2885), .Z(n2884) );
  XNOR U2956 ( .A(n2887), .B(n2888), .Z(n2886) );
  NANDN U2957 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR U2958 ( .A(n2892), .B(n2893), .Z(n2881) );
  XOR U2959 ( .A(key[245]), .B(n2894), .Z(n2893) );
  ANDN U2960 ( .B(n2895), .A(n2896), .Z(n2892) );
  XNOR U2961 ( .A(n2897), .B(n2898), .Z(out[116]) );
  XNOR U2962 ( .A(key[244]), .B(n2899), .Z(n2898) );
  XOR U2963 ( .A(n2900), .B(n2901), .Z(out[115]) );
  XNOR U2964 ( .A(n2902), .B(n2878), .Z(n2901) );
  XNOR U2965 ( .A(n2903), .B(n2904), .Z(n2878) );
  XNOR U2966 ( .A(n2905), .B(n2894), .Z(n2904) );
  ANDN U2967 ( .B(n2906), .A(n2907), .Z(n2894) );
  NOR U2968 ( .A(n2908), .B(n2909), .Z(n2905) );
  XNOR U2969 ( .A(n2910), .B(n2911), .Z(n2900) );
  XOR U2970 ( .A(key[243]), .B(n2877), .Z(n2911) );
  XOR U2971 ( .A(key[242]), .B(n2897), .Z(out[114]) );
  XNOR U2972 ( .A(n2912), .B(n2913), .Z(n2897) );
  XOR U2973 ( .A(n2914), .B(n2874), .Z(out[113]) );
  XNOR U2974 ( .A(n2903), .B(n2915), .Z(n2902) );
  XNOR U2975 ( .A(n2916), .B(n2917), .Z(n2915) );
  NANDN U2976 ( .A(n2918), .B(n2890), .Z(n2917) );
  XNOR U2977 ( .A(n2885), .B(n2919), .Z(n2903) );
  XNOR U2978 ( .A(n2920), .B(n2921), .Z(n2919) );
  NANDN U2979 ( .A(n2922), .B(n2923), .Z(n2921) );
  XOR U2980 ( .A(n2913), .B(n2910), .Z(n2880) );
  XNOR U2981 ( .A(n2885), .B(n2924), .Z(n2910) );
  XNOR U2982 ( .A(n2916), .B(n2925), .Z(n2924) );
  NANDN U2983 ( .A(n2926), .B(n2927), .Z(n2925) );
  OR U2984 ( .A(n2928), .B(n2929), .Z(n2916) );
  XOR U2985 ( .A(n2930), .B(n2920), .Z(n2885) );
  NANDN U2986 ( .A(n2931), .B(n2932), .Z(n2920) );
  ANDN U2987 ( .B(n2933), .A(n2934), .Z(n2930) );
  XNOR U2988 ( .A(key[241]), .B(n2912), .Z(n2914) );
  IV U2989 ( .A(n2877), .Z(n2912) );
  XOR U2990 ( .A(n2935), .B(n2936), .Z(n2877) );
  XNOR U2991 ( .A(n2937), .B(n2938), .Z(n2936) );
  NANDN U2992 ( .A(n2939), .B(n2895), .Z(n2938) );
  XNOR U2993 ( .A(n2883), .B(n2940), .Z(out[112]) );
  XOR U2994 ( .A(key[240]), .B(n2913), .Z(n2940) );
  XNOR U2995 ( .A(n2935), .B(n2941), .Z(n2913) );
  XOR U2996 ( .A(n2942), .B(n2887), .Z(n2941) );
  OR U2997 ( .A(n2943), .B(n2928), .Z(n2887) );
  XNOR U2998 ( .A(n2890), .B(n2927), .Z(n2928) );
  ANDN U2999 ( .B(n2944), .A(n2945), .Z(n2942) );
  IV U3000 ( .A(n2899), .Z(n2883) );
  XOR U3001 ( .A(n2891), .B(n2946), .Z(n2899) );
  XOR U3002 ( .A(n2947), .B(n2937), .Z(n2946) );
  XNOR U3003 ( .A(n2909), .B(n2895), .Z(n2906) );
  NOR U3004 ( .A(n2949), .B(n2909), .Z(n2947) );
  XNOR U3005 ( .A(n2935), .B(n2950), .Z(n2891) );
  XNOR U3006 ( .A(n2951), .B(n2952), .Z(n2950) );
  NANDN U3007 ( .A(n2922), .B(n2953), .Z(n2952) );
  XOR U3008 ( .A(n2954), .B(n2951), .Z(n2935) );
  OR U3009 ( .A(n2931), .B(n2955), .Z(n2951) );
  XOR U3010 ( .A(n2956), .B(n2922), .Z(n2931) );
  XNOR U3011 ( .A(n2927), .B(n2895), .Z(n2922) );
  XOR U3012 ( .A(n2957), .B(n2958), .Z(n2895) );
  NANDN U3013 ( .A(n2959), .B(n2960), .Z(n2958) );
  IV U3014 ( .A(n2945), .Z(n2927) );
  XNOR U3015 ( .A(n2961), .B(n2962), .Z(n2945) );
  NANDN U3016 ( .A(n2959), .B(n2963), .Z(n2962) );
  ANDN U3017 ( .B(n2956), .A(n2964), .Z(n2954) );
  IV U3018 ( .A(n2934), .Z(n2956) );
  XOR U3019 ( .A(n2909), .B(n2890), .Z(n2934) );
  XNOR U3020 ( .A(n2965), .B(n2961), .Z(n2890) );
  NANDN U3021 ( .A(n2966), .B(n2967), .Z(n2961) );
  XOR U3022 ( .A(n2963), .B(n2968), .Z(n2967) );
  ANDN U3023 ( .B(n2968), .A(n2969), .Z(n2965) );
  XOR U3024 ( .A(n2970), .B(n2957), .Z(n2909) );
  NANDN U3025 ( .A(n2966), .B(n2971), .Z(n2957) );
  XOR U3026 ( .A(n2972), .B(n2960), .Z(n2971) );
  XNOR U3027 ( .A(n2973), .B(n2974), .Z(n2959) );
  XOR U3028 ( .A(n2975), .B(n2976), .Z(n2974) );
  XNOR U3029 ( .A(n2977), .B(n2978), .Z(n2973) );
  XNOR U3030 ( .A(n2979), .B(n2980), .Z(n2978) );
  ANDN U3031 ( .B(n2972), .A(n2976), .Z(n2979) );
  ANDN U3032 ( .B(n2972), .A(n2969), .Z(n2970) );
  XNOR U3033 ( .A(n2975), .B(n2981), .Z(n2969) );
  XOR U3034 ( .A(n2982), .B(n2980), .Z(n2981) );
  NAND U3035 ( .A(n2983), .B(n2984), .Z(n2980) );
  XNOR U3036 ( .A(n2977), .B(n2960), .Z(n2984) );
  IV U3037 ( .A(n2972), .Z(n2977) );
  XNOR U3038 ( .A(n2963), .B(n2976), .Z(n2983) );
  IV U3039 ( .A(n2968), .Z(n2976) );
  XOR U3040 ( .A(n2985), .B(n2986), .Z(n2968) );
  XNOR U3041 ( .A(n2987), .B(n2988), .Z(n2986) );
  XNOR U3042 ( .A(n2989), .B(n2990), .Z(n2985) );
  ANDN U3043 ( .B(n2991), .A(n2949), .Z(n2989) );
  AND U3044 ( .A(n2960), .B(n2963), .Z(n2982) );
  XNOR U3045 ( .A(n2960), .B(n2963), .Z(n2975) );
  XNOR U3046 ( .A(n2992), .B(n2993), .Z(n2963) );
  XNOR U3047 ( .A(n2994), .B(n2988), .Z(n2993) );
  XOR U3048 ( .A(n2995), .B(n2996), .Z(n2992) );
  XNOR U3049 ( .A(n2997), .B(n2990), .Z(n2996) );
  OR U3050 ( .A(n2907), .B(n2948), .Z(n2990) );
  XNOR U3051 ( .A(n2998), .B(n2999), .Z(n2948) );
  XNOR U3052 ( .A(n2908), .B(n2896), .Z(n2907) );
  ANDN U3053 ( .B(n3000), .A(n2939), .Z(n2997) );
  XNOR U3054 ( .A(n3001), .B(n3002), .Z(n2960) );
  XNOR U3055 ( .A(n2988), .B(n3003), .Z(n3002) );
  XOR U3056 ( .A(n2918), .B(n2995), .Z(n3003) );
  XNOR U3057 ( .A(n2998), .B(n2908), .Z(n2988) );
  XNOR U3058 ( .A(n3004), .B(n3005), .Z(n3001) );
  XNOR U3059 ( .A(n3006), .B(n3007), .Z(n3005) );
  ANDN U3060 ( .B(n2944), .A(n2926), .Z(n3006) );
  XNOR U3061 ( .A(n3008), .B(n3009), .Z(n2972) );
  XNOR U3062 ( .A(n2994), .B(n3010), .Z(n3009) );
  XNOR U3063 ( .A(n2926), .B(n2987), .Z(n3010) );
  XOR U3064 ( .A(n2995), .B(n3011), .Z(n2987) );
  XNOR U3065 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U3066 ( .A(n2953), .B(n2923), .Z(n3013) );
  XNOR U3067 ( .A(n3014), .B(n3012), .Z(n2995) );
  NANDN U3068 ( .A(n2955), .B(n2932), .Z(n3012) );
  XOR U3069 ( .A(n2933), .B(n2923), .Z(n2932) );
  XNOR U3070 ( .A(n3015), .B(n2896), .Z(n2923) );
  XOR U3071 ( .A(n2964), .B(n2953), .Z(n2955) );
  XOR U3072 ( .A(n2944), .B(n2999), .Z(n2953) );
  ANDN U3073 ( .B(n2933), .A(n2964), .Z(n3014) );
  XNOR U3074 ( .A(n3004), .B(n2998), .Z(n2964) );
  IV U3075 ( .A(n2949), .Z(n2998) );
  XNOR U3076 ( .A(n3016), .B(n3017), .Z(n2949) );
  XOR U3077 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U3078 ( .A(n3020), .B(n2991), .Z(n2933) );
  XOR U3079 ( .A(n2999), .B(n3000), .Z(n2994) );
  IV U3080 ( .A(n2896), .Z(n3000) );
  XOR U3081 ( .A(n3021), .B(n3022), .Z(n2896) );
  XNOR U3082 ( .A(n3023), .B(n3019), .Z(n3022) );
  IV U3083 ( .A(n2939), .Z(n2999) );
  XOR U3084 ( .A(n3019), .B(n3024), .Z(n2939) );
  XNOR U3085 ( .A(n2944), .B(n3025), .Z(n3008) );
  XNOR U3086 ( .A(n3026), .B(n3007), .Z(n3025) );
  OR U3087 ( .A(n2929), .B(n2943), .Z(n3007) );
  XNOR U3088 ( .A(n3004), .B(n2944), .Z(n2943) );
  XOR U3089 ( .A(n2918), .B(n3015), .Z(n2929) );
  IV U3090 ( .A(n2926), .Z(n3015) );
  XOR U3091 ( .A(n2991), .B(n3027), .Z(n2926) );
  XOR U3092 ( .A(n3023), .B(n3016), .Z(n3027) );
  XNOR U3093 ( .A(key[210]), .B(\w0[1][82] ), .Z(n3016) );
  XNOR U3094 ( .A(n1638), .B(n3028), .Z(\w0[1][82] ) );
  XOR U3095 ( .A(n3029), .B(n211), .Z(n3028) );
  XOR U3096 ( .A(n179), .B(n3030), .Z(n211) );
  IV U3097 ( .A(n2908), .Z(n2991) );
  XOR U3098 ( .A(n3021), .B(n3031), .Z(n2908) );
  XOR U3099 ( .A(n3019), .B(n3032), .Z(n3031) );
  ANDN U3100 ( .B(n3020), .A(n2889), .Z(n3026) );
  IV U3101 ( .A(n2918), .Z(n3020) );
  XOR U3102 ( .A(n3021), .B(n3033), .Z(n2918) );
  XOR U3103 ( .A(n3019), .B(n3034), .Z(n3033) );
  XOR U3104 ( .A(n2889), .B(n3035), .Z(n3019) );
  XOR U3105 ( .A(key[214]), .B(\w0[1][86] ), .Z(n3035) );
  XNOR U3106 ( .A(n3036), .B(n3037), .Z(\w0[1][86] ) );
  XNOR U3107 ( .A(n3038), .B(n185), .Z(n3037) );
  XOR U3108 ( .A(n1626), .B(n3039), .Z(n185) );
  IV U3109 ( .A(n3004), .Z(n2889) );
  IV U3110 ( .A(n3024), .Z(n3021) );
  XOR U3111 ( .A(key[213]), .B(\w0[1][85] ), .Z(n3024) );
  XNOR U3112 ( .A(n3040), .B(n3041), .Z(\w0[1][85] ) );
  XOR U3113 ( .A(n1612), .B(n1618), .Z(n3041) );
  XNOR U3114 ( .A(n193), .B(n3038), .Z(n1612) );
  XOR U3115 ( .A(n3042), .B(n3043), .Z(n2944) );
  XNOR U3116 ( .A(n3034), .B(n3032), .Z(n3043) );
  XNOR U3117 ( .A(key[215]), .B(\w0[1][87] ), .Z(n3032) );
  XNOR U3118 ( .A(n3044), .B(n3045), .Z(\w0[1][87] ) );
  XNOR U3119 ( .A(n224), .B(n3046), .Z(n3045) );
  XNOR U3120 ( .A(key[212]), .B(\w0[1][84] ), .Z(n3034) );
  XOR U3121 ( .A(n3047), .B(n3048), .Z(\w0[1][84] ) );
  XNOR U3122 ( .A(n3049), .B(n3050), .Z(n3048) );
  XOR U3123 ( .A(n206), .B(n1631), .Z(n3047) );
  XOR U3124 ( .A(n224), .B(n1617), .Z(n206) );
  IV U3125 ( .A(n3039), .Z(n224) );
  XNOR U3126 ( .A(n3004), .B(n3018), .Z(n3042) );
  XOR U3127 ( .A(n3023), .B(n3051), .Z(n3018) );
  XOR U3128 ( .A(key[211]), .B(\w0[1][83] ), .Z(n3051) );
  XOR U3129 ( .A(n3052), .B(n3053), .Z(\w0[1][83] ) );
  XOR U3130 ( .A(n1602), .B(n3054), .Z(n3053) );
  XOR U3131 ( .A(n213), .B(n3030), .Z(n3052) );
  IV U3132 ( .A(n3055), .Z(n3030) );
  XNOR U3133 ( .A(n3039), .B(n1632), .Z(n213) );
  XOR U3134 ( .A(key[209]), .B(\w0[1][81] ), .Z(n3023) );
  XNOR U3135 ( .A(n1640), .B(n3056), .Z(\w0[1][81] ) );
  XNOR U3136 ( .A(n176), .B(n3057), .Z(n3056) );
  IV U3137 ( .A(n1604), .Z(n176) );
  XNOR U3138 ( .A(n3029), .B(n218), .Z(n1604) );
  XOR U3139 ( .A(key[208]), .B(\w0[1][80] ), .Z(n3004) );
  XOR U3140 ( .A(n222), .B(n3058), .Z(\w0[1][80] ) );
  XNOR U3141 ( .A(n1623), .B(n217), .Z(n3058) );
  XNOR U3142 ( .A(n3057), .B(n225), .Z(n217) );
  IV U3143 ( .A(n1633), .Z(n1623) );
  XOR U3144 ( .A(n3059), .B(n3060), .Z(out[111]) );
  XOR U3145 ( .A(n3061), .B(n3062), .Z(n3059) );
  XOR U3146 ( .A(key[239]), .B(n3063), .Z(n3062) );
  XNOR U3147 ( .A(n3064), .B(n3065), .Z(out[110]) );
  XNOR U3148 ( .A(key[238]), .B(n3066), .Z(n3065) );
  XOR U3149 ( .A(key[138]), .B(n2060), .Z(out[10]) );
  XNOR U3150 ( .A(n2044), .B(n4), .Z(n2060) );
  XNOR U3151 ( .A(n2067), .B(n3067), .Z(n4) );
  XNOR U3152 ( .A(n2064), .B(n3068), .Z(n3067) );
  NANDN U3153 ( .A(n3069), .B(n2059), .Z(n3068) );
  XNOR U3154 ( .A(n2066), .B(n2059), .Z(n2850) );
  XNOR U3155 ( .A(n2067), .B(n3071), .Z(n2044) );
  XOR U3156 ( .A(n3072), .B(n2051), .Z(n3071) );
  OR U3157 ( .A(n2866), .B(n3073), .Z(n2051) );
  XNOR U3158 ( .A(n2053), .B(n2864), .Z(n2866) );
  NOR U3159 ( .A(n3074), .B(n2864), .Z(n3072) );
  XOR U3160 ( .A(n3075), .B(n2069), .Z(n2067) );
  NANDN U3161 ( .A(n2870), .B(n3076), .Z(n2069) );
  XNOR U3162 ( .A(n2871), .B(n2071), .Z(n2870) );
  XNOR U3163 ( .A(n2864), .B(n2059), .Z(n2071) );
  XOR U3164 ( .A(n3077), .B(n3078), .Z(n2059) );
  NANDN U3165 ( .A(n3079), .B(n3080), .Z(n3078) );
  XNOR U3166 ( .A(n3081), .B(n3082), .Z(n2864) );
  OR U3167 ( .A(n3079), .B(n3083), .Z(n3082) );
  AND U3168 ( .A(n2871), .B(n3084), .Z(n3075) );
  XOR U3169 ( .A(n2053), .B(n2066), .Z(n2871) );
  XOR U3170 ( .A(n3085), .B(n3077), .Z(n2066) );
  NANDN U3171 ( .A(n3086), .B(n3087), .Z(n3077) );
  ANDN U3172 ( .B(n3088), .A(n3089), .Z(n3085) );
  NANDN U3173 ( .A(n3086), .B(n3091), .Z(n3081) );
  XOR U3174 ( .A(n3092), .B(n3079), .Z(n3086) );
  XNOR U3175 ( .A(n3093), .B(n3094), .Z(n3079) );
  XOR U3176 ( .A(n3095), .B(n3088), .Z(n3094) );
  XNOR U3177 ( .A(n3096), .B(n3097), .Z(n3093) );
  XNOR U3178 ( .A(n3098), .B(n3099), .Z(n3097) );
  ANDN U3179 ( .B(n3088), .A(n3100), .Z(n3098) );
  IV U3180 ( .A(n3101), .Z(n3088) );
  ANDN U3181 ( .B(n3092), .A(n3100), .Z(n3090) );
  IV U3182 ( .A(n3096), .Z(n3100) );
  IV U3183 ( .A(n3089), .Z(n3092) );
  XNOR U3184 ( .A(n3095), .B(n3102), .Z(n3089) );
  XOR U3185 ( .A(n3103), .B(n3099), .Z(n3102) );
  NAND U3186 ( .A(n3091), .B(n3087), .Z(n3099) );
  XNOR U3187 ( .A(n3080), .B(n3101), .Z(n3087) );
  XOR U3188 ( .A(n3104), .B(n3105), .Z(n3101) );
  XOR U3189 ( .A(n3106), .B(n3107), .Z(n3105) );
  XOR U3190 ( .A(n3108), .B(n3109), .Z(n3107) );
  XOR U3191 ( .A(n2865), .B(n3110), .Z(n3104) );
  XNOR U3192 ( .A(n3111), .B(n3112), .Z(n3110) );
  ANDN U3193 ( .B(n2857), .A(n2054), .Z(n3111) );
  XNOR U3194 ( .A(n3096), .B(n3083), .Z(n3091) );
  XOR U3195 ( .A(n3113), .B(n3114), .Z(n3096) );
  XNOR U3196 ( .A(n3115), .B(n3109), .Z(n3114) );
  XOR U3197 ( .A(n3116), .B(n3117), .Z(n3109) );
  XNOR U3198 ( .A(n3118), .B(n3119), .Z(n3117) );
  NAND U3199 ( .A(n2072), .B(n2861), .Z(n3119) );
  XNOR U3200 ( .A(n3120), .B(n3121), .Z(n3113) );
  ANDN U3201 ( .B(n2065), .A(n2852), .Z(n3120) );
  ANDN U3202 ( .B(n3080), .A(n3083), .Z(n3103) );
  XOR U3203 ( .A(n3083), .B(n3080), .Z(n3095) );
  XNOR U3204 ( .A(n3122), .B(n3123), .Z(n3080) );
  XNOR U3205 ( .A(n3116), .B(n3124), .Z(n3123) );
  XNOR U3206 ( .A(n2857), .B(n3115), .Z(n3124) );
  XOR U3207 ( .A(n2054), .B(n3125), .Z(n3122) );
  XNOR U3208 ( .A(n3126), .B(n3112), .Z(n3125) );
  OR U3209 ( .A(n2867), .B(n3073), .Z(n3112) );
  XNOR U3210 ( .A(n3127), .B(n3108), .Z(n3073) );
  XNOR U3211 ( .A(n2857), .B(n2865), .Z(n2867) );
  ANDN U3212 ( .B(n2865), .A(n3074), .Z(n3126) );
  IV U3213 ( .A(n3108), .Z(n3074) );
  XOR U3214 ( .A(n3128), .B(n3129), .Z(n3083) );
  XOR U3215 ( .A(n3116), .B(n3106), .Z(n3129) );
  XOR U3216 ( .A(n2058), .B(n3069), .Z(n3106) );
  XOR U3217 ( .A(n3130), .B(n3118), .Z(n3116) );
  NANDN U3218 ( .A(n2869), .B(n3076), .Z(n3118) );
  XOR U3219 ( .A(n3084), .B(n2072), .Z(n3076) );
  XNOR U3220 ( .A(n3069), .B(n3108), .Z(n2072) );
  XOR U3221 ( .A(n3131), .B(n3132), .Z(n3108) );
  XNOR U3222 ( .A(n3133), .B(n3134), .Z(n3132) );
  XOR U3223 ( .A(n3127), .B(n3135), .Z(n3131) );
  XOR U3224 ( .A(n2872), .B(n2861), .Z(n2869) );
  XOR U3225 ( .A(n2058), .B(n2865), .Z(n2861) );
  XOR U3226 ( .A(n3136), .B(n3137), .Z(n2865) );
  XNOR U3227 ( .A(n2852), .B(n3138), .Z(n3137) );
  ANDN U3228 ( .B(n3084), .A(n2872), .Z(n3130) );
  XOR U3229 ( .A(n2852), .B(n2857), .Z(n2872) );
  XOR U3230 ( .A(n3133), .B(n3139), .Z(n2857) );
  XOR U3231 ( .A(key[204]), .B(\w0[1][76] ), .Z(n3133) );
  XOR U3232 ( .A(n3140), .B(n3141), .Z(\w0[1][76] ) );
  XOR U3233 ( .A(n3050), .B(n1630), .Z(n3141) );
  XNOR U3234 ( .A(n194), .B(n1621), .Z(n1630) );
  XOR U3235 ( .A(n203), .B(n1629), .Z(n3050) );
  XNOR U3236 ( .A(n3142), .B(n219), .Z(n1629) );
  XNOR U3237 ( .A(n1632), .B(n3049), .Z(n3140) );
  XNOR U3238 ( .A(n1618), .B(n3143), .Z(n3049) );
  XNOR U3239 ( .A(n3144), .B(n3145), .Z(n1618) );
  XNOR U3240 ( .A(n3146), .B(n3147), .Z(n3145) );
  XOR U3241 ( .A(n3148), .B(n3149), .Z(n3144) );
  XNOR U3242 ( .A(n3150), .B(n3151), .Z(n3149) );
  ANDN U3243 ( .B(n3152), .A(n3153), .Z(n3151) );
  XOR U3244 ( .A(n3154), .B(n218), .Z(n1632) );
  XOR U3245 ( .A(n3127), .B(n2065), .Z(n3084) );
  XOR U3246 ( .A(n3115), .B(n3155), .Z(n3128) );
  XNOR U3247 ( .A(n3156), .B(n3121), .Z(n3155) );
  OR U3248 ( .A(n3070), .B(n2851), .Z(n3121) );
  XOR U3249 ( .A(n2852), .B(n2058), .Z(n2851) );
  XNOR U3250 ( .A(n2065), .B(n3139), .Z(n3070) );
  ANDN U3251 ( .B(n2058), .A(n3069), .Z(n3156) );
  IV U3252 ( .A(n3139), .Z(n3069) );
  XOR U3253 ( .A(n3138), .B(n3139), .Z(n2058) );
  XOR U3254 ( .A(n2852), .B(n2065), .Z(n3115) );
  XNOR U3255 ( .A(n3134), .B(n3157), .Z(n2065) );
  XNOR U3256 ( .A(n3158), .B(n3136), .Z(n3157) );
  XOR U3257 ( .A(key[202]), .B(\w0[1][74] ), .Z(n3136) );
  XOR U3258 ( .A(n3159), .B(n3160), .Z(\w0[1][74] ) );
  XOR U3259 ( .A(n3055), .B(n1638), .Z(n3160) );
  XOR U3260 ( .A(n178), .B(n219), .Z(n1638) );
  XNOR U3261 ( .A(n3161), .B(n3162), .Z(n219) );
  XNOR U3262 ( .A(n3163), .B(n3164), .Z(n3055) );
  XOR U3263 ( .A(n3165), .B(n3166), .Z(n3164) );
  XOR U3264 ( .A(n3167), .B(n3168), .Z(n3163) );
  XNOR U3265 ( .A(n218), .B(n210), .Z(n3159) );
  XOR U3266 ( .A(n3169), .B(n3170), .Z(n218) );
  XNOR U3267 ( .A(n3138), .B(n3171), .Z(n3134) );
  XOR U3268 ( .A(key[203]), .B(\w0[1][75] ), .Z(n3171) );
  XOR U3269 ( .A(n3172), .B(n3173), .Z(\w0[1][75] ) );
  XOR U3270 ( .A(n3054), .B(n1637), .Z(n3173) );
  XNOR U3271 ( .A(n203), .B(n1621), .Z(n1637) );
  XOR U3272 ( .A(n3174), .B(n3175), .Z(n203) );
  XNOR U3273 ( .A(n1631), .B(n1642), .Z(n3054) );
  XNOR U3274 ( .A(n3147), .B(n3029), .Z(n1631) );
  XNOR U3275 ( .A(n179), .B(n1602), .Z(n3172) );
  XNOR U3276 ( .A(n210), .B(n177), .Z(n1602) );
  XNOR U3277 ( .A(n3176), .B(n3177), .Z(n177) );
  XOR U3278 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U3279 ( .A(n3162), .B(n3180), .Z(n3176) );
  XOR U3280 ( .A(n3181), .B(n3182), .Z(n210) );
  XOR U3281 ( .A(n3185), .B(n3186), .Z(n3181) );
  XOR U3282 ( .A(n3187), .B(n3188), .Z(n179) );
  XOR U3283 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U3284 ( .A(n3169), .B(n3191), .Z(n3187) );
  XOR U3285 ( .A(key[201]), .B(\w0[1][73] ), .Z(n3138) );
  XOR U3286 ( .A(n3192), .B(n3193), .Z(\w0[1][73] ) );
  XOR U3287 ( .A(n225), .B(n1640), .Z(n3193) );
  XNOR U3288 ( .A(n216), .B(n223), .Z(n1640) );
  XNOR U3289 ( .A(n3194), .B(n3195), .Z(n223) );
  XNOR U3290 ( .A(n3162), .B(n3180), .Z(n3195) );
  XOR U3291 ( .A(n3196), .B(n3197), .Z(n225) );
  XNOR U3292 ( .A(n3169), .B(n3191), .Z(n3197) );
  XNOR U3293 ( .A(n3175), .B(n3029), .Z(n3192) );
  XOR U3294 ( .A(n3167), .B(n3198), .Z(n3029) );
  IV U3295 ( .A(n178), .Z(n3175) );
  XNOR U3296 ( .A(n3135), .B(n3139), .Z(n2852) );
  XNOR U3297 ( .A(n3200), .B(n3158), .Z(n3139) );
  XOR U3298 ( .A(n2054), .B(n3201), .Z(n3158) );
  XOR U3299 ( .A(key[206]), .B(\w0[1][78] ), .Z(n3201) );
  XNOR U3300 ( .A(n1610), .B(n3202), .Z(\w0[1][78] ) );
  XNOR U3301 ( .A(n193), .B(n3036), .Z(n3202) );
  XOR U3302 ( .A(n3046), .B(n1614), .Z(n3036) );
  XOR U3303 ( .A(n188), .B(n192), .Z(n1614) );
  XOR U3304 ( .A(n3203), .B(n3179), .Z(n192) );
  XNOR U3305 ( .A(n3204), .B(n3205), .Z(n3179) );
  XOR U3306 ( .A(n3206), .B(n3207), .Z(n3205) );
  NOR U3307 ( .A(n3208), .B(n3209), .Z(n3206) );
  XNOR U3308 ( .A(n1625), .B(n1642), .Z(n3046) );
  XOR U3309 ( .A(n3210), .B(n3211), .Z(n1625) );
  XOR U3310 ( .A(n3212), .B(n3165), .Z(n3211) );
  XNOR U3311 ( .A(n3214), .B(n3215), .Z(n3213) );
  NANDN U3312 ( .A(n3216), .B(n3217), .Z(n3215) );
  XOR U3313 ( .A(n3196), .B(n3190), .Z(n193) );
  XNOR U3314 ( .A(n3219), .B(n3220), .Z(n3190) );
  XOR U3315 ( .A(n3221), .B(n3222), .Z(n3220) );
  NOR U3316 ( .A(n3223), .B(n3224), .Z(n3221) );
  XNOR U3317 ( .A(n199), .B(n3225), .Z(n1610) );
  IV U3318 ( .A(n3127), .Z(n2054) );
  XOR U3319 ( .A(key[200]), .B(\w0[1][72] ), .Z(n3127) );
  XOR U3320 ( .A(n3226), .B(n3227), .Z(\w0[1][72] ) );
  XNOR U3321 ( .A(n3057), .B(n3225), .Z(n3227) );
  IV U3322 ( .A(n1621), .Z(n3225) );
  XOR U3323 ( .A(n3165), .B(n3228), .Z(n3057) );
  XOR U3324 ( .A(n3167), .B(n3212), .Z(n3228) );
  XOR U3325 ( .A(n3229), .B(n3230), .Z(n3167) );
  XOR U3326 ( .A(n3231), .B(n3232), .Z(n3230) );
  ANDN U3327 ( .B(n3233), .A(n3153), .Z(n3231) );
  XOR U3328 ( .A(n3234), .B(n3235), .Z(n3165) );
  XOR U3329 ( .A(n3236), .B(n3237), .Z(n3235) );
  ANDN U3330 ( .B(n3238), .A(n3216), .Z(n3236) );
  XOR U3331 ( .A(n197), .B(n216), .Z(n3226) );
  XOR U3332 ( .A(n3184), .B(n3239), .Z(n216) );
  XOR U3333 ( .A(n3240), .B(n3186), .Z(n3239) );
  XOR U3334 ( .A(n1633), .B(n3039), .Z(n197) );
  XOR U3335 ( .A(n3170), .B(n3154), .Z(n3039) );
  XOR U3336 ( .A(key[205]), .B(\w0[1][77] ), .Z(n3200) );
  XOR U3337 ( .A(n3241), .B(n3242), .Z(\w0[1][77] ) );
  XOR U3338 ( .A(n1617), .B(n3040), .Z(n3242) );
  XOR U3339 ( .A(n194), .B(n1616), .Z(n3040) );
  XNOR U3340 ( .A(n3243), .B(n3244), .Z(n1616) );
  XNOR U3341 ( .A(n3245), .B(n3246), .Z(n3244) );
  XNOR U3342 ( .A(n3142), .B(n3247), .Z(n3243) );
  XNOR U3343 ( .A(n3207), .B(n3248), .Z(n3247) );
  ANDN U3344 ( .B(n3249), .A(n3250), .Z(n3248) );
  NANDN U3345 ( .A(n3251), .B(n3252), .Z(n3207) );
  XNOR U3346 ( .A(n3253), .B(n3254), .Z(n3142) );
  XNOR U3347 ( .A(n3255), .B(n3256), .Z(n3254) );
  NOR U3348 ( .A(n3257), .B(n3209), .Z(n3255) );
  XOR U3349 ( .A(n3258), .B(n3259), .Z(n194) );
  XNOR U3350 ( .A(n3260), .B(n3174), .Z(n3259) );
  XNOR U3351 ( .A(n3261), .B(n3262), .Z(n3258) );
  XNOR U3352 ( .A(n3263), .B(n3264), .Z(n3262) );
  ANDN U3353 ( .B(n3265), .A(n3266), .Z(n3263) );
  XNOR U3354 ( .A(n3267), .B(n3268), .Z(n1617) );
  XOR U3355 ( .A(n3269), .B(n3154), .Z(n3268) );
  XOR U3356 ( .A(n3270), .B(n3271), .Z(n3154) );
  XNOR U3357 ( .A(n3272), .B(n3273), .Z(n3271) );
  NOR U3358 ( .A(n3274), .B(n3224), .Z(n3272) );
  XNOR U3359 ( .A(n3275), .B(n3276), .Z(n3267) );
  XNOR U3360 ( .A(n3222), .B(n3277), .Z(n3276) );
  ANDN U3361 ( .B(n3278), .A(n3279), .Z(n3277) );
  NANDN U3362 ( .A(n3280), .B(n3281), .Z(n3222) );
  XNOR U3363 ( .A(n3038), .B(n188), .Z(n3241) );
  XOR U3364 ( .A(n3183), .B(n3240), .Z(n188) );
  XNOR U3365 ( .A(n3282), .B(n3283), .Z(n3183) );
  XNOR U3366 ( .A(n3264), .B(n3284), .Z(n3283) );
  NAND U3367 ( .A(n3285), .B(n3286), .Z(n3284) );
  NANDN U3368 ( .A(n3287), .B(n3288), .Z(n3264) );
  XNOR U3369 ( .A(n3166), .B(n3212), .Z(n3038) );
  XOR U3370 ( .A(n3168), .B(n3198), .Z(n3212) );
  XOR U3371 ( .A(n3146), .B(n3289), .Z(n3168) );
  XNOR U3372 ( .A(n3237), .B(n3290), .Z(n3289) );
  NAND U3373 ( .A(n3291), .B(n3292), .Z(n3290) );
  OR U3374 ( .A(n3293), .B(n3294), .Z(n3237) );
  XNOR U3375 ( .A(n3234), .B(n3295), .Z(n3166) );
  XOR U3376 ( .A(n3296), .B(n3150), .Z(n3295) );
  OR U3377 ( .A(n3297), .B(n3298), .Z(n3150) );
  ANDN U3378 ( .B(n3299), .A(n3300), .Z(n3296) );
  XNOR U3379 ( .A(n3146), .B(n3301), .Z(n3234) );
  XNOR U3380 ( .A(n3302), .B(n3303), .Z(n3301) );
  NAND U3381 ( .A(n3304), .B(n3305), .Z(n3303) );
  XOR U3382 ( .A(n3306), .B(n3302), .Z(n3146) );
  NANDN U3383 ( .A(n3307), .B(n3308), .Z(n3302) );
  ANDN U3384 ( .B(n3309), .A(n3310), .Z(n3306) );
  XOR U3385 ( .A(key[207]), .B(\w0[1][79] ), .Z(n3135) );
  XNOR U3386 ( .A(n3044), .B(n3311), .Z(\w0[1][79] ) );
  XOR U3387 ( .A(n1626), .B(n222), .Z(n3311) );
  XOR U3388 ( .A(n1621), .B(n3143), .Z(n222) );
  IV U3389 ( .A(n1642), .Z(n3143) );
  XNOR U3390 ( .A(n3198), .B(n3147), .Z(n1642) );
  XNOR U3391 ( .A(n3218), .B(n3312), .Z(n3147) );
  XNOR U3392 ( .A(n3232), .B(n3313), .Z(n3312) );
  NANDN U3393 ( .A(n3314), .B(n3299), .Z(n3313) );
  OR U3394 ( .A(n3315), .B(n3297), .Z(n3232) );
  XNOR U3395 ( .A(n3299), .B(n3316), .Z(n3297) );
  XNOR U3396 ( .A(n3229), .B(n3317), .Z(n3218) );
  XNOR U3397 ( .A(n3318), .B(n3319), .Z(n3317) );
  NAND U3398 ( .A(n3305), .B(n3320), .Z(n3319) );
  XNOR U3399 ( .A(n3229), .B(n3321), .Z(n3198) );
  XOR U3400 ( .A(n3322), .B(n3214), .Z(n3321) );
  OR U3401 ( .A(n3323), .B(n3293), .Z(n3214) );
  XOR U3402 ( .A(n3216), .B(n3292), .Z(n3293) );
  ANDN U3403 ( .B(n3292), .A(n3324), .Z(n3322) );
  XOR U3404 ( .A(n3325), .B(n3318), .Z(n3229) );
  OR U3405 ( .A(n3307), .B(n3326), .Z(n3318) );
  XNOR U3406 ( .A(n3327), .B(n3305), .Z(n3307) );
  XNOR U3407 ( .A(n3292), .B(n3153), .Z(n3305) );
  IV U3408 ( .A(n3316), .Z(n3153) );
  XOR U3409 ( .A(n3328), .B(n3329), .Z(n3316) );
  NAND U3410 ( .A(n3330), .B(n3331), .Z(n3329) );
  XOR U3411 ( .A(n3332), .B(n3333), .Z(n3292) );
  NANDN U3412 ( .A(n3334), .B(n3330), .Z(n3333) );
  ANDN U3413 ( .B(n3327), .A(n3335), .Z(n3325) );
  IV U3414 ( .A(n3310), .Z(n3327) );
  XOR U3415 ( .A(n3216), .B(n3299), .Z(n3310) );
  XOR U3416 ( .A(n3328), .B(n3336), .Z(n3299) );
  NANDN U3417 ( .A(n3337), .B(n3338), .Z(n3336) );
  NAND U3418 ( .A(n3339), .B(n3340), .Z(n3328) );
  NANDN U3419 ( .A(n3342), .B(n3340), .Z(n3332) );
  XNOR U3420 ( .A(n3337), .B(n3330), .Z(n3340) );
  XNOR U3421 ( .A(n3343), .B(n3344), .Z(n3330) );
  XOR U3422 ( .A(n3345), .B(n3338), .Z(n3344) );
  IV U3423 ( .A(n3346), .Z(n3338) );
  XNOR U3424 ( .A(n3347), .B(n3348), .Z(n3343) );
  XNOR U3425 ( .A(n3349), .B(n3350), .Z(n3348) );
  NOR U3426 ( .A(n3346), .B(n3347), .Z(n3349) );
  NOR U3427 ( .A(n3337), .B(n3347), .Z(n3341) );
  XNOR U3428 ( .A(n3345), .B(n3351), .Z(n3337) );
  XNOR U3429 ( .A(n3350), .B(n3352), .Z(n3351) );
  NANDN U3430 ( .A(n3334), .B(n3331), .Z(n3352) );
  NANDN U3431 ( .A(n3342), .B(n3339), .Z(n3350) );
  XNOR U3432 ( .A(n3331), .B(n3346), .Z(n3339) );
  XOR U3433 ( .A(n3353), .B(n3354), .Z(n3346) );
  XOR U3434 ( .A(n3355), .B(n3356), .Z(n3354) );
  XOR U3435 ( .A(n3291), .B(n3357), .Z(n3356) );
  XNOR U3436 ( .A(n3324), .B(n3358), .Z(n3353) );
  XNOR U3437 ( .A(n3359), .B(n3360), .Z(n3358) );
  AND U3438 ( .A(n3217), .B(n3238), .Z(n3359) );
  XOR U3439 ( .A(n3361), .B(n3362), .Z(n3347) );
  XNOR U3440 ( .A(n3363), .B(n3357), .Z(n3362) );
  XNOR U3441 ( .A(n3364), .B(n3365), .Z(n3357) );
  XNOR U3442 ( .A(n3366), .B(n3367), .Z(n3365) );
  NAND U3443 ( .A(n3320), .B(n3304), .Z(n3367) );
  XNOR U3444 ( .A(n3368), .B(n3369), .Z(n3361) );
  ANDN U3445 ( .B(n3370), .A(n3300), .Z(n3368) );
  XOR U3446 ( .A(n3334), .B(n3331), .Z(n3345) );
  XNOR U3447 ( .A(n3371), .B(n3372), .Z(n3331) );
  XOR U3448 ( .A(n3373), .B(n3374), .Z(n3372) );
  XOR U3449 ( .A(n3363), .B(n3238), .Z(n3374) );
  XOR U3450 ( .A(n3217), .B(n3375), .Z(n3371) );
  XNOR U3451 ( .A(n3376), .B(n3360), .Z(n3375) );
  OR U3452 ( .A(n3294), .B(n3323), .Z(n3360) );
  XNOR U3453 ( .A(n3217), .B(n3377), .Z(n3323) );
  XNOR U3454 ( .A(n3238), .B(n3291), .Z(n3294) );
  ANDN U3455 ( .B(n3291), .A(n3324), .Z(n3376) );
  XOR U3456 ( .A(n3378), .B(n3379), .Z(n3334) );
  XOR U3457 ( .A(n3364), .B(n3355), .Z(n3379) );
  XOR U3458 ( .A(n3233), .B(n3152), .Z(n3355) );
  IV U3459 ( .A(n3373), .Z(n3364) );
  XNOR U3460 ( .A(n3380), .B(n3366), .Z(n3373) );
  NANDN U3461 ( .A(n3326), .B(n3308), .Z(n3366) );
  XOR U3462 ( .A(n3309), .B(n3304), .Z(n3308) );
  XOR U3463 ( .A(n3152), .B(n3291), .Z(n3304) );
  XNOR U3464 ( .A(n3381), .B(n3382), .Z(n3291) );
  XOR U3465 ( .A(n3383), .B(n3384), .Z(n3382) );
  IV U3466 ( .A(n3385), .Z(n3152) );
  XOR U3467 ( .A(n3335), .B(n3320), .Z(n3326) );
  XNOR U3468 ( .A(n3377), .B(n3386), .Z(n3320) );
  IV U3469 ( .A(n3324), .Z(n3377) );
  XOR U3470 ( .A(n3387), .B(n3388), .Z(n3324) );
  XOR U3471 ( .A(n3389), .B(n3390), .Z(n3388) );
  XOR U3472 ( .A(n3217), .B(n3391), .Z(n3387) );
  ANDN U3473 ( .B(n3309), .A(n3335), .Z(n3380) );
  XNOR U3474 ( .A(n3217), .B(n3370), .Z(n3335) );
  XOR U3475 ( .A(n3381), .B(n3238), .Z(n3309) );
  XNOR U3476 ( .A(n3392), .B(n3393), .Z(n3238) );
  XOR U3477 ( .A(n3394), .B(n3390), .Z(n3393) );
  XOR U3478 ( .A(state[12]), .B(key[12]), .Z(n3390) );
  IV U3479 ( .A(n3300), .Z(n3381) );
  XNOR U3480 ( .A(n3363), .B(n3395), .Z(n3378) );
  XNOR U3481 ( .A(n3396), .B(n3369), .Z(n3395) );
  OR U3482 ( .A(n3298), .B(n3315), .Z(n3369) );
  XNOR U3483 ( .A(n3314), .B(n3386), .Z(n3315) );
  IV U3484 ( .A(n3233), .Z(n3386) );
  IV U3485 ( .A(n3370), .Z(n3314) );
  XNOR U3486 ( .A(n3300), .B(n3385), .Z(n3298) );
  ANDN U3487 ( .B(n3233), .A(n3385), .Z(n3396) );
  XOR U3488 ( .A(n3392), .B(n3397), .Z(n3385) );
  XOR U3489 ( .A(n3383), .B(n3398), .Z(n3397) );
  XOR U3490 ( .A(n3370), .B(n3300), .Z(n3363) );
  XOR U3491 ( .A(n3392), .B(n3399), .Z(n3300) );
  XNOR U3492 ( .A(n3394), .B(n3389), .Z(n3399) );
  XNOR U3493 ( .A(state[15]), .B(key[15]), .Z(n3389) );
  XOR U3494 ( .A(state[13]), .B(key[13]), .Z(n3392) );
  XNOR U3495 ( .A(n3384), .B(n3400), .Z(n3370) );
  XNOR U3496 ( .A(n3391), .B(n3398), .Z(n3400) );
  IV U3497 ( .A(n3394), .Z(n3398) );
  XOR U3498 ( .A(n3217), .B(n3401), .Z(n3394) );
  XNOR U3499 ( .A(state[14]), .B(key[14]), .Z(n3401) );
  XOR U3500 ( .A(state[8]), .B(key[8]), .Z(n3217) );
  XOR U3501 ( .A(n3383), .B(n3402), .Z(n3391) );
  XNOR U3502 ( .A(state[11]), .B(key[11]), .Z(n3402) );
  XNOR U3503 ( .A(state[9]), .B(key[9]), .Z(n3383) );
  XOR U3504 ( .A(state[10]), .B(key[10]), .Z(n3384) );
  XOR U3505 ( .A(n3199), .B(n3174), .Z(n1621) );
  XNOR U3506 ( .A(n3403), .B(n3404), .Z(n3174) );
  XOR U3507 ( .A(n3405), .B(n3406), .Z(n3404) );
  ANDN U3508 ( .B(n3286), .A(n3407), .Z(n3405) );
  XOR U3509 ( .A(n3408), .B(n3409), .Z(n1626) );
  XOR U3510 ( .A(n3191), .B(n3196), .Z(n3409) );
  XOR U3511 ( .A(n3170), .B(n3189), .Z(n3196) );
  XNOR U3512 ( .A(n3269), .B(n3410), .Z(n3189) );
  XNOR U3513 ( .A(n3411), .B(n3412), .Z(n3410) );
  NANDN U3514 ( .A(n3413), .B(n3414), .Z(n3412) );
  XOR U3515 ( .A(n3415), .B(n3416), .Z(n3170) );
  XOR U3516 ( .A(n3417), .B(n3418), .Z(n3416) );
  ANDN U3517 ( .B(n3419), .A(n3413), .Z(n3417) );
  XNOR U3518 ( .A(n3219), .B(n3420), .Z(n3191) );
  XNOR U3519 ( .A(n3411), .B(n3421), .Z(n3420) );
  OR U3520 ( .A(n3422), .B(n3423), .Z(n3421) );
  OR U3521 ( .A(n3424), .B(n3425), .Z(n3411) );
  XOR U3522 ( .A(n3269), .B(n3426), .Z(n3219) );
  XNOR U3523 ( .A(n3427), .B(n3428), .Z(n3426) );
  OR U3524 ( .A(n3429), .B(n3430), .Z(n3428) );
  XOR U3525 ( .A(n3431), .B(n3427), .Z(n3269) );
  NANDN U3526 ( .A(n3432), .B(n3433), .Z(n3427) );
  AND U3527 ( .A(n3434), .B(n3435), .Z(n3431) );
  XOR U3528 ( .A(n3415), .B(n3436), .Z(n3169) );
  XOR U3529 ( .A(n3273), .B(n3437), .Z(n3436) );
  OR U3530 ( .A(n3438), .B(n3279), .Z(n3437) );
  ANDN U3531 ( .B(n3281), .A(n3439), .Z(n3273) );
  XOR U3532 ( .A(n3224), .B(n3279), .Z(n3281) );
  XNOR U3533 ( .A(n3270), .B(n3440), .Z(n3275) );
  XNOR U3534 ( .A(n3418), .B(n3441), .Z(n3440) );
  OR U3535 ( .A(n3422), .B(n3442), .Z(n3441) );
  OR U3536 ( .A(n3443), .B(n3424), .Z(n3418) );
  XOR U3537 ( .A(n3422), .B(n3444), .Z(n3424) );
  XNOR U3538 ( .A(n3415), .B(n3445), .Z(n3270) );
  XNOR U3539 ( .A(n3446), .B(n3447), .Z(n3445) );
  NANDN U3540 ( .A(n3429), .B(n3448), .Z(n3447) );
  XOR U3541 ( .A(n3449), .B(n3446), .Z(n3415) );
  OR U3542 ( .A(n3432), .B(n3450), .Z(n3446) );
  XOR U3543 ( .A(n3434), .B(n3429), .Z(n3432) );
  XOR U3544 ( .A(n3444), .B(n3279), .Z(n3429) );
  XNOR U3545 ( .A(n3451), .B(n3452), .Z(n3279) );
  NANDN U3546 ( .A(n3453), .B(n3454), .Z(n3452) );
  IV U3547 ( .A(n3413), .Z(n3444) );
  XNOR U3548 ( .A(n3455), .B(n3456), .Z(n3413) );
  NANDN U3549 ( .A(n3453), .B(n3457), .Z(n3456) );
  ANDN U3550 ( .B(n3434), .A(n3458), .Z(n3449) );
  XOR U3551 ( .A(n3224), .B(n3422), .Z(n3434) );
  XOR U3552 ( .A(n3459), .B(n3455), .Z(n3422) );
  NANDN U3553 ( .A(n3460), .B(n3461), .Z(n3455) );
  NANDN U3554 ( .A(n3460), .B(n3465), .Z(n3451) );
  XOR U3555 ( .A(n3466), .B(n3467), .Z(n3453) );
  XOR U3556 ( .A(n3468), .B(n3463), .Z(n3467) );
  XNOR U3557 ( .A(n3469), .B(n3470), .Z(n3466) );
  XNOR U3558 ( .A(n3471), .B(n3472), .Z(n3470) );
  ANDN U3559 ( .B(n3468), .A(n3463), .Z(n3471) );
  ANDN U3560 ( .B(n3468), .A(n3462), .Z(n3464) );
  XNOR U3561 ( .A(n3469), .B(n3473), .Z(n3462) );
  XOR U3562 ( .A(n3474), .B(n3472), .Z(n3473) );
  NAND U3563 ( .A(n3461), .B(n3465), .Z(n3472) );
  XNOR U3564 ( .A(n3457), .B(n3463), .Z(n3461) );
  XOR U3565 ( .A(n3475), .B(n3476), .Z(n3463) );
  XOR U3566 ( .A(n3477), .B(n3478), .Z(n3476) );
  XNOR U3567 ( .A(n3479), .B(n3480), .Z(n3475) );
  ANDN U3568 ( .B(n3481), .A(n3223), .Z(n3479) );
  AND U3569 ( .A(n3454), .B(n3457), .Z(n3474) );
  XNOR U3570 ( .A(n3454), .B(n3457), .Z(n3469) );
  XNOR U3571 ( .A(n3482), .B(n3483), .Z(n3457) );
  XNOR U3572 ( .A(n3484), .B(n3485), .Z(n3483) );
  XOR U3573 ( .A(n3477), .B(n3486), .Z(n3482) );
  XNOR U3574 ( .A(n3487), .B(n3480), .Z(n3486) );
  OR U3575 ( .A(n3280), .B(n3439), .Z(n3480) );
  XNOR U3576 ( .A(n3274), .B(n3438), .Z(n3439) );
  XNOR U3577 ( .A(n3223), .B(n3488), .Z(n3280) );
  NOR U3578 ( .A(n3488), .B(n3438), .Z(n3487) );
  XNOR U3579 ( .A(n3489), .B(n3490), .Z(n3454) );
  XNOR U3580 ( .A(n3491), .B(n3492), .Z(n3490) );
  XOR U3581 ( .A(n3423), .B(n3477), .Z(n3492) );
  XOR U3582 ( .A(n3481), .B(n3493), .Z(n3477) );
  XNOR U3583 ( .A(n3442), .B(n3494), .Z(n3489) );
  XNOR U3584 ( .A(n3495), .B(n3496), .Z(n3494) );
  ANDN U3585 ( .B(n3414), .A(n3497), .Z(n3495) );
  XNOR U3586 ( .A(n3498), .B(n3499), .Z(n3468) );
  XNOR U3587 ( .A(n3478), .B(n3500), .Z(n3499) );
  XNOR U3588 ( .A(n3414), .B(n3485), .Z(n3500) );
  XOR U3589 ( .A(n3438), .B(n3488), .Z(n3485) );
  XNOR U3590 ( .A(n3491), .B(n3501), .Z(n3478) );
  XNOR U3591 ( .A(n3502), .B(n3503), .Z(n3501) );
  NANDN U3592 ( .A(n3430), .B(n3448), .Z(n3503) );
  IV U3593 ( .A(n3484), .Z(n3491) );
  XNOR U3594 ( .A(n3504), .B(n3502), .Z(n3484) );
  NANDN U3595 ( .A(n3450), .B(n3433), .Z(n3502) );
  XOR U3596 ( .A(n3414), .B(n3488), .Z(n3430) );
  IV U3597 ( .A(n3278), .Z(n3488) );
  XOR U3598 ( .A(n3505), .B(n3506), .Z(n3278) );
  XNOR U3599 ( .A(n3507), .B(n3508), .Z(n3506) );
  XOR U3600 ( .A(n3458), .B(n3448), .Z(n3450) );
  XNOR U3601 ( .A(n3419), .B(n3438), .Z(n3448) );
  XNOR U3602 ( .A(n3508), .B(n3505), .Z(n3438) );
  ANDN U3603 ( .B(n3435), .A(n3458), .Z(n3504) );
  XNOR U3604 ( .A(n3509), .B(n3481), .Z(n3458) );
  IV U3605 ( .A(n3274), .Z(n3481) );
  XNOR U3606 ( .A(n3510), .B(n3511), .Z(n3274) );
  XNOR U3607 ( .A(n3512), .B(n3508), .Z(n3511) );
  XOR U3608 ( .A(n3513), .B(n3493), .Z(n3435) );
  XNOR U3609 ( .A(n3497), .B(n3514), .Z(n3498) );
  XNOR U3610 ( .A(n3515), .B(n3496), .Z(n3514) );
  OR U3611 ( .A(n3425), .B(n3443), .Z(n3496) );
  XOR U3612 ( .A(n3442), .B(n3419), .Z(n3443) );
  IV U3613 ( .A(n3497), .Z(n3419) );
  XOR U3614 ( .A(n3423), .B(n3414), .Z(n3425) );
  XNOR U3615 ( .A(n3493), .B(n3516), .Z(n3414) );
  XNOR U3616 ( .A(n3507), .B(n3510), .Z(n3516) );
  XNOR U3617 ( .A(state[50]), .B(key[50]), .Z(n3510) );
  IV U3618 ( .A(n3223), .Z(n3493) );
  XOR U3619 ( .A(n3517), .B(n3518), .Z(n3223) );
  XOR U3620 ( .A(n3508), .B(n3519), .Z(n3518) );
  IV U3621 ( .A(n3513), .Z(n3423) );
  ANDN U3622 ( .B(n3513), .A(n3442), .Z(n3515) );
  XOR U3623 ( .A(n3505), .B(n3520), .Z(n3513) );
  XNOR U3624 ( .A(n3508), .B(n3521), .Z(n3520) );
  XOR U3625 ( .A(n3509), .B(n3522), .Z(n3508) );
  XNOR U3626 ( .A(state[54]), .B(key[54]), .Z(n3522) );
  IV U3627 ( .A(n3517), .Z(n3505) );
  XOR U3628 ( .A(state[53]), .B(key[53]), .Z(n3517) );
  XOR U3629 ( .A(n3523), .B(n3524), .Z(n3497) );
  XOR U3630 ( .A(n3521), .B(n3519), .Z(n3524) );
  XOR U3631 ( .A(state[55]), .B(key[55]), .Z(n3519) );
  XNOR U3632 ( .A(state[52]), .B(key[52]), .Z(n3521) );
  XOR U3633 ( .A(n3442), .B(n3512), .Z(n3523) );
  XNOR U3634 ( .A(n3507), .B(n3525), .Z(n3512) );
  XNOR U3635 ( .A(state[51]), .B(key[51]), .Z(n3525) );
  XNOR U3636 ( .A(state[49]), .B(key[49]), .Z(n3507) );
  IV U3637 ( .A(n3509), .Z(n3442) );
  XOR U3638 ( .A(state[48]), .B(key[48]), .Z(n3509) );
  XOR U3639 ( .A(n199), .B(n1624), .Z(n3044) );
  XNOR U3640 ( .A(n3526), .B(n3527), .Z(n1624) );
  XOR U3641 ( .A(n3180), .B(n3194), .Z(n3527) );
  IV U3642 ( .A(n3203), .Z(n3194) );
  XOR U3643 ( .A(n3161), .B(n3178), .Z(n3203) );
  XNOR U3644 ( .A(n3246), .B(n3528), .Z(n3178) );
  XNOR U3645 ( .A(n3529), .B(n3530), .Z(n3528) );
  NANDN U3646 ( .A(n3531), .B(n3532), .Z(n3530) );
  XNOR U3647 ( .A(n3533), .B(n3534), .Z(n3161) );
  XOR U3648 ( .A(n3535), .B(n3536), .Z(n3534) );
  ANDN U3649 ( .B(n3537), .A(n3531), .Z(n3535) );
  XNOR U3650 ( .A(n3204), .B(n3538), .Z(n3180) );
  XNOR U3651 ( .A(n3529), .B(n3539), .Z(n3538) );
  OR U3652 ( .A(n3540), .B(n3541), .Z(n3539) );
  OR U3653 ( .A(n3542), .B(n3543), .Z(n3529) );
  XOR U3654 ( .A(n3246), .B(n3544), .Z(n3204) );
  XNOR U3655 ( .A(n3545), .B(n3546), .Z(n3544) );
  OR U3656 ( .A(n3547), .B(n3548), .Z(n3546) );
  XOR U3657 ( .A(n3549), .B(n3545), .Z(n3246) );
  NANDN U3658 ( .A(n3550), .B(n3551), .Z(n3545) );
  AND U3659 ( .A(n3552), .B(n3553), .Z(n3549) );
  XNOR U3660 ( .A(n3245), .B(n3162), .Z(n3526) );
  XOR U3661 ( .A(n3533), .B(n3554), .Z(n3162) );
  XOR U3662 ( .A(n3256), .B(n3555), .Z(n3554) );
  OR U3663 ( .A(n3556), .B(n3250), .Z(n3555) );
  ANDN U3664 ( .B(n3252), .A(n3557), .Z(n3256) );
  XOR U3665 ( .A(n3209), .B(n3250), .Z(n3252) );
  XNOR U3666 ( .A(n3253), .B(n3558), .Z(n3245) );
  XNOR U3667 ( .A(n3536), .B(n3559), .Z(n3558) );
  OR U3668 ( .A(n3540), .B(n3560), .Z(n3559) );
  OR U3669 ( .A(n3561), .B(n3542), .Z(n3536) );
  XOR U3670 ( .A(n3540), .B(n3562), .Z(n3542) );
  XNOR U3671 ( .A(n3533), .B(n3563), .Z(n3253) );
  XNOR U3672 ( .A(n3564), .B(n3565), .Z(n3563) );
  NANDN U3673 ( .A(n3547), .B(n3566), .Z(n3565) );
  XOR U3674 ( .A(n3567), .B(n3564), .Z(n3533) );
  OR U3675 ( .A(n3550), .B(n3568), .Z(n3564) );
  XOR U3676 ( .A(n3552), .B(n3547), .Z(n3550) );
  XOR U3677 ( .A(n3562), .B(n3250), .Z(n3547) );
  XNOR U3678 ( .A(n3569), .B(n3570), .Z(n3250) );
  NANDN U3679 ( .A(n3571), .B(n3572), .Z(n3570) );
  IV U3680 ( .A(n3531), .Z(n3562) );
  XNOR U3681 ( .A(n3573), .B(n3574), .Z(n3531) );
  NANDN U3682 ( .A(n3571), .B(n3575), .Z(n3574) );
  ANDN U3683 ( .B(n3552), .A(n3576), .Z(n3567) );
  XOR U3684 ( .A(n3209), .B(n3540), .Z(n3552) );
  XOR U3685 ( .A(n3577), .B(n3573), .Z(n3540) );
  NANDN U3686 ( .A(n3578), .B(n3579), .Z(n3573) );
  NANDN U3687 ( .A(n3578), .B(n3583), .Z(n3569) );
  XOR U3688 ( .A(n3584), .B(n3585), .Z(n3571) );
  XOR U3689 ( .A(n3586), .B(n3581), .Z(n3585) );
  XNOR U3690 ( .A(n3587), .B(n3588), .Z(n3584) );
  XNOR U3691 ( .A(n3589), .B(n3590), .Z(n3588) );
  ANDN U3692 ( .B(n3586), .A(n3581), .Z(n3589) );
  ANDN U3693 ( .B(n3586), .A(n3580), .Z(n3582) );
  XNOR U3694 ( .A(n3587), .B(n3591), .Z(n3580) );
  XOR U3695 ( .A(n3592), .B(n3590), .Z(n3591) );
  NAND U3696 ( .A(n3579), .B(n3583), .Z(n3590) );
  XNOR U3697 ( .A(n3575), .B(n3581), .Z(n3579) );
  XOR U3698 ( .A(n3593), .B(n3594), .Z(n3581) );
  XOR U3699 ( .A(n3595), .B(n3596), .Z(n3594) );
  XNOR U3700 ( .A(n3597), .B(n3598), .Z(n3593) );
  ANDN U3701 ( .B(n3599), .A(n3208), .Z(n3597) );
  AND U3702 ( .A(n3572), .B(n3575), .Z(n3592) );
  XNOR U3703 ( .A(n3572), .B(n3575), .Z(n3587) );
  XNOR U3704 ( .A(n3600), .B(n3601), .Z(n3575) );
  XNOR U3705 ( .A(n3602), .B(n3603), .Z(n3601) );
  XOR U3706 ( .A(n3595), .B(n3604), .Z(n3600) );
  XNOR U3707 ( .A(n3605), .B(n3598), .Z(n3604) );
  OR U3708 ( .A(n3251), .B(n3557), .Z(n3598) );
  XNOR U3709 ( .A(n3257), .B(n3556), .Z(n3557) );
  XNOR U3710 ( .A(n3208), .B(n3606), .Z(n3251) );
  NOR U3711 ( .A(n3606), .B(n3556), .Z(n3605) );
  XNOR U3712 ( .A(n3607), .B(n3608), .Z(n3572) );
  XNOR U3713 ( .A(n3609), .B(n3610), .Z(n3608) );
  XOR U3714 ( .A(n3541), .B(n3595), .Z(n3610) );
  XOR U3715 ( .A(n3599), .B(n3611), .Z(n3595) );
  XNOR U3716 ( .A(n3560), .B(n3612), .Z(n3607) );
  XNOR U3717 ( .A(n3613), .B(n3614), .Z(n3612) );
  ANDN U3718 ( .B(n3532), .A(n3615), .Z(n3613) );
  XNOR U3719 ( .A(n3616), .B(n3617), .Z(n3586) );
  XNOR U3720 ( .A(n3596), .B(n3618), .Z(n3617) );
  XNOR U3721 ( .A(n3532), .B(n3603), .Z(n3618) );
  XOR U3722 ( .A(n3556), .B(n3606), .Z(n3603) );
  XNOR U3723 ( .A(n3609), .B(n3619), .Z(n3596) );
  XNOR U3724 ( .A(n3620), .B(n3621), .Z(n3619) );
  NANDN U3725 ( .A(n3548), .B(n3566), .Z(n3621) );
  IV U3726 ( .A(n3602), .Z(n3609) );
  XNOR U3727 ( .A(n3622), .B(n3620), .Z(n3602) );
  NANDN U3728 ( .A(n3568), .B(n3551), .Z(n3620) );
  XOR U3729 ( .A(n3532), .B(n3606), .Z(n3548) );
  IV U3730 ( .A(n3249), .Z(n3606) );
  XOR U3731 ( .A(n3623), .B(n3624), .Z(n3249) );
  XNOR U3732 ( .A(n3625), .B(n3626), .Z(n3624) );
  XOR U3733 ( .A(n3576), .B(n3566), .Z(n3568) );
  XNOR U3734 ( .A(n3537), .B(n3556), .Z(n3566) );
  XNOR U3735 ( .A(n3626), .B(n3623), .Z(n3556) );
  ANDN U3736 ( .B(n3553), .A(n3576), .Z(n3622) );
  XNOR U3737 ( .A(n3627), .B(n3599), .Z(n3576) );
  IV U3738 ( .A(n3257), .Z(n3599) );
  XNOR U3739 ( .A(n3628), .B(n3629), .Z(n3257) );
  XNOR U3740 ( .A(n3630), .B(n3626), .Z(n3629) );
  XOR U3741 ( .A(n3631), .B(n3611), .Z(n3553) );
  XNOR U3742 ( .A(n3615), .B(n3632), .Z(n3616) );
  XNOR U3743 ( .A(n3633), .B(n3614), .Z(n3632) );
  OR U3744 ( .A(n3543), .B(n3561), .Z(n3614) );
  XOR U3745 ( .A(n3560), .B(n3537), .Z(n3561) );
  IV U3746 ( .A(n3615), .Z(n3537) );
  XOR U3747 ( .A(n3541), .B(n3532), .Z(n3543) );
  XNOR U3748 ( .A(n3611), .B(n3634), .Z(n3532) );
  XNOR U3749 ( .A(n3625), .B(n3628), .Z(n3634) );
  XNOR U3750 ( .A(state[90]), .B(key[90]), .Z(n3628) );
  IV U3751 ( .A(n3208), .Z(n3611) );
  XOR U3752 ( .A(n3635), .B(n3636), .Z(n3208) );
  XOR U3753 ( .A(n3626), .B(n3637), .Z(n3636) );
  IV U3754 ( .A(n3631), .Z(n3541) );
  ANDN U3755 ( .B(n3631), .A(n3560), .Z(n3633) );
  XOR U3756 ( .A(n3623), .B(n3638), .Z(n3631) );
  XNOR U3757 ( .A(n3626), .B(n3639), .Z(n3638) );
  XOR U3758 ( .A(n3627), .B(n3640), .Z(n3626) );
  XNOR U3759 ( .A(state[94]), .B(key[94]), .Z(n3640) );
  IV U3760 ( .A(n3635), .Z(n3623) );
  XOR U3761 ( .A(state[93]), .B(key[93]), .Z(n3635) );
  XOR U3762 ( .A(n3641), .B(n3642), .Z(n3615) );
  XOR U3763 ( .A(n3639), .B(n3637), .Z(n3642) );
  XOR U3764 ( .A(state[95]), .B(key[95]), .Z(n3637) );
  XNOR U3765 ( .A(state[92]), .B(key[92]), .Z(n3639) );
  XOR U3766 ( .A(n3560), .B(n3630), .Z(n3641) );
  XNOR U3767 ( .A(n3625), .B(n3643), .Z(n3630) );
  XNOR U3768 ( .A(state[91]), .B(key[91]), .Z(n3643) );
  XNOR U3769 ( .A(state[89]), .B(key[89]), .Z(n3625) );
  IV U3770 ( .A(n3627), .Z(n3560) );
  XOR U3771 ( .A(state[88]), .B(key[88]), .Z(n3627) );
  XOR U3772 ( .A(n3644), .B(n3645), .Z(n199) );
  XNOR U3773 ( .A(n3186), .B(n3184), .Z(n3645) );
  XOR U3774 ( .A(n3646), .B(n3647), .Z(n3184) );
  XNOR U3775 ( .A(n3406), .B(n3648), .Z(n3647) );
  NANDN U3776 ( .A(n3650), .B(n3288), .Z(n3406) );
  XNOR U3777 ( .A(n3286), .B(n3266), .Z(n3288) );
  XOR U3778 ( .A(n3282), .B(n3651), .Z(n3186) );
  XNOR U3779 ( .A(n3652), .B(n3653), .Z(n3651) );
  NANDN U3780 ( .A(n3654), .B(n3655), .Z(n3653) );
  XNOR U3781 ( .A(n3261), .B(n3656), .Z(n3282) );
  XNOR U3782 ( .A(n3657), .B(n3658), .Z(n3656) );
  NANDN U3783 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U3784 ( .A(n3240), .B(n3260), .Z(n3644) );
  XNOR U3785 ( .A(n3403), .B(n3661), .Z(n3260) );
  XNOR U3786 ( .A(n3662), .B(n3663), .Z(n3661) );
  NANDN U3787 ( .A(n3654), .B(n3664), .Z(n3663) );
  XNOR U3788 ( .A(n3646), .B(n3665), .Z(n3403) );
  XNOR U3789 ( .A(n3666), .B(n3667), .Z(n3665) );
  NANDN U3790 ( .A(n3659), .B(n3668), .Z(n3667) );
  XOR U3791 ( .A(n3199), .B(n3185), .Z(n3240) );
  XOR U3792 ( .A(n3261), .B(n3669), .Z(n3185) );
  XOR U3793 ( .A(n3670), .B(n3652), .Z(n3669) );
  OR U3794 ( .A(n3671), .B(n3672), .Z(n3652) );
  ANDN U3795 ( .B(n3673), .A(n3674), .Z(n3670) );
  XOR U3796 ( .A(n3675), .B(n3657), .Z(n3261) );
  NANDN U3797 ( .A(n3676), .B(n3677), .Z(n3657) );
  ANDN U3798 ( .B(n3678), .A(n3679), .Z(n3675) );
  XNOR U3799 ( .A(n3646), .B(n3680), .Z(n3199) );
  XOR U3800 ( .A(n3681), .B(n3662), .Z(n3680) );
  OR U3801 ( .A(n3682), .B(n3671), .Z(n3662) );
  XOR U3802 ( .A(n3654), .B(n3683), .Z(n3671) );
  ANDN U3803 ( .B(n3684), .A(n3674), .Z(n3681) );
  IV U3804 ( .A(n3683), .Z(n3674) );
  XOR U3805 ( .A(n3685), .B(n3666), .Z(n3646) );
  OR U3806 ( .A(n3676), .B(n3686), .Z(n3666) );
  XOR U3807 ( .A(n3687), .B(n3659), .Z(n3676) );
  XOR U3808 ( .A(n3683), .B(n3266), .Z(n3659) );
  XNOR U3809 ( .A(n3688), .B(n3689), .Z(n3266) );
  NANDN U3810 ( .A(n3690), .B(n3691), .Z(n3689) );
  XOR U3811 ( .A(n3692), .B(n3693), .Z(n3683) );
  NANDN U3812 ( .A(n3690), .B(n3694), .Z(n3693) );
  ANDN U3813 ( .B(n3687), .A(n3695), .Z(n3685) );
  IV U3814 ( .A(n3679), .Z(n3687) );
  XOR U3815 ( .A(n3654), .B(n3286), .Z(n3679) );
  XNOR U3816 ( .A(n3696), .B(n3688), .Z(n3286) );
  NANDN U3817 ( .A(n3697), .B(n3698), .Z(n3688) );
  XOR U3818 ( .A(n3691), .B(n3699), .Z(n3698) );
  ANDN U3819 ( .B(n3699), .A(n3700), .Z(n3696) );
  NANDN U3820 ( .A(n3697), .B(n3702), .Z(n3692) );
  XOR U3821 ( .A(n3703), .B(n3704), .Z(n3690) );
  XOR U3822 ( .A(n3705), .B(n3706), .Z(n3704) );
  XNOR U3823 ( .A(n3707), .B(n3708), .Z(n3703) );
  XNOR U3824 ( .A(n3709), .B(n3710), .Z(n3708) );
  ANDN U3825 ( .B(n3706), .A(n3705), .Z(n3709) );
  ANDN U3826 ( .B(n3706), .A(n3700), .Z(n3701) );
  XNOR U3827 ( .A(n3707), .B(n3711), .Z(n3700) );
  XOR U3828 ( .A(n3712), .B(n3710), .Z(n3711) );
  NAND U3829 ( .A(n3702), .B(n3713), .Z(n3710) );
  XNOR U3830 ( .A(n3691), .B(n3705), .Z(n3713) );
  IV U3831 ( .A(n3699), .Z(n3705) );
  XNOR U3832 ( .A(n3714), .B(n3715), .Z(n3699) );
  XNOR U3833 ( .A(n3716), .B(n3717), .Z(n3715) );
  XOR U3834 ( .A(n3718), .B(n3719), .Z(n3717) );
  XNOR U3835 ( .A(n3720), .B(n3721), .Z(n3714) );
  XNOR U3836 ( .A(n3722), .B(n3723), .Z(n3721) );
  AND U3837 ( .A(n3655), .B(n3664), .Z(n3722) );
  XOR U3838 ( .A(n3694), .B(n3706), .Z(n3702) );
  AND U3839 ( .A(n3691), .B(n3694), .Z(n3712) );
  XNOR U3840 ( .A(n3691), .B(n3694), .Z(n3707) );
  XNOR U3841 ( .A(n3724), .B(n3725), .Z(n3694) );
  XNOR U3842 ( .A(n3726), .B(n3719), .Z(n3725) );
  XOR U3843 ( .A(n3727), .B(n3728), .Z(n3724) );
  XNOR U3844 ( .A(n3729), .B(n3730), .Z(n3728) );
  ANDN U3845 ( .B(n3265), .A(n3649), .Z(n3729) );
  XNOR U3846 ( .A(n3731), .B(n3732), .Z(n3691) );
  XNOR U3847 ( .A(n3655), .B(n3727), .Z(n3733) );
  XOR U3848 ( .A(n3664), .B(n3734), .Z(n3731) );
  XNOR U3849 ( .A(n3735), .B(n3723), .Z(n3734) );
  OR U3850 ( .A(n3672), .B(n3682), .Z(n3723) );
  XOR U3851 ( .A(n3664), .B(n3720), .Z(n3682) );
  XNOR U3852 ( .A(n3655), .B(n3673), .Z(n3672) );
  ANDN U3853 ( .B(n3684), .A(n3718), .Z(n3735) );
  XNOR U3854 ( .A(n3736), .B(n3737), .Z(n3706) );
  XOR U3855 ( .A(n3726), .B(n3716), .Z(n3737) );
  XOR U3856 ( .A(n3727), .B(n3738), .Z(n3716) );
  XNOR U3857 ( .A(n3739), .B(n3740), .Z(n3738) );
  NAND U3858 ( .A(n3668), .B(n3660), .Z(n3740) );
  XNOR U3859 ( .A(n3741), .B(n3739), .Z(n3727) );
  NANDN U3860 ( .A(n3686), .B(n3677), .Z(n3739) );
  XOR U3861 ( .A(n3678), .B(n3660), .Z(n3677) );
  XOR U3862 ( .A(n3673), .B(n3265), .Z(n3660) );
  IV U3863 ( .A(n3718), .Z(n3673) );
  XOR U3864 ( .A(n3285), .B(n3742), .Z(n3718) );
  XNOR U3865 ( .A(n3743), .B(n3744), .Z(n3742) );
  XOR U3866 ( .A(n3695), .B(n3668), .Z(n3686) );
  XNOR U3867 ( .A(n3684), .B(n3649), .Z(n3668) );
  IV U3868 ( .A(n3720), .Z(n3684) );
  XOR U3869 ( .A(n3745), .B(n3746), .Z(n3720) );
  XOR U3870 ( .A(n3747), .B(n3748), .Z(n3746) );
  XOR U3871 ( .A(n3664), .B(n3749), .Z(n3745) );
  ANDN U3872 ( .B(n3678), .A(n3695), .Z(n3741) );
  XNOR U3873 ( .A(n3664), .B(n3750), .Z(n3695) );
  XOR U3874 ( .A(n3655), .B(n3285), .Z(n3678) );
  XOR U3875 ( .A(n3751), .B(n3752), .Z(n3655) );
  XOR U3876 ( .A(n3753), .B(n3748), .Z(n3752) );
  XOR U3877 ( .A(state[100]), .B(key[100]), .Z(n3748) );
  XOR U3878 ( .A(n3750), .B(n3285), .Z(n3726) );
  IV U3879 ( .A(n3407), .Z(n3750) );
  XNOR U3880 ( .A(n3754), .B(n3730), .Z(n3736) );
  OR U3881 ( .A(n3287), .B(n3650), .Z(n3730) );
  XNOR U3882 ( .A(n3407), .B(n3649), .Z(n3650) );
  XOR U3883 ( .A(n3755), .B(n3751), .Z(n3649) );
  XNOR U3884 ( .A(n3285), .B(n3265), .Z(n3287) );
  XOR U3885 ( .A(n3751), .B(n3756), .Z(n3265) );
  XOR U3886 ( .A(n3744), .B(n3755), .Z(n3756) );
  ANDN U3887 ( .B(n3285), .A(n3407), .Z(n3754) );
  XOR U3888 ( .A(n3755), .B(n3757), .Z(n3407) );
  XOR U3889 ( .A(n3743), .B(n3749), .Z(n3757) );
  XOR U3890 ( .A(n3744), .B(n3758), .Z(n3749) );
  XNOR U3891 ( .A(state[99]), .B(key[99]), .Z(n3758) );
  XNOR U3892 ( .A(state[97]), .B(key[97]), .Z(n3744) );
  XNOR U3893 ( .A(state[98]), .B(key[98]), .Z(n3743) );
  IV U3894 ( .A(n3753), .Z(n3755) );
  XOR U3895 ( .A(n3751), .B(n3759), .Z(n3285) );
  XNOR U3896 ( .A(n3753), .B(n3747), .Z(n3759) );
  XNOR U3897 ( .A(state[103]), .B(key[103]), .Z(n3747) );
  XOR U3898 ( .A(n3664), .B(n3760), .Z(n3753) );
  XNOR U3899 ( .A(state[102]), .B(key[102]), .Z(n3760) );
  XOR U3900 ( .A(state[96]), .B(key[96]), .Z(n3664) );
  XNOR U3901 ( .A(state[101]), .B(key[101]), .Z(n3751) );
  XOR U3902 ( .A(n3761), .B(n3762), .Z(out[109]) );
  XNOR U3903 ( .A(n3763), .B(n3764), .Z(n3762) );
  XOR U3904 ( .A(n3061), .B(n3765), .Z(n3764) );
  XNOR U3905 ( .A(n3767), .B(n3768), .Z(n3766) );
  NANDN U3906 ( .A(n3769), .B(n3770), .Z(n3768) );
  XOR U3907 ( .A(n3772), .B(n3773), .Z(n3761) );
  XOR U3908 ( .A(key[237]), .B(n3774), .Z(n3773) );
  ANDN U3909 ( .B(n3775), .A(n3776), .Z(n3772) );
  XNOR U3910 ( .A(n3777), .B(n3778), .Z(out[108]) );
  XNOR U3911 ( .A(key[236]), .B(n3779), .Z(n3778) );
  XOR U3912 ( .A(n3780), .B(n3781), .Z(out[107]) );
  XNOR U3913 ( .A(n3782), .B(n3064), .Z(n3781) );
  XNOR U3914 ( .A(n3783), .B(n3784), .Z(n3064) );
  XNOR U3915 ( .A(n3785), .B(n3774), .Z(n3784) );
  ANDN U3916 ( .B(n3786), .A(n3787), .Z(n3774) );
  NOR U3917 ( .A(n3788), .B(n3789), .Z(n3785) );
  XNOR U3918 ( .A(n3790), .B(n3791), .Z(n3780) );
  XOR U3919 ( .A(key[235]), .B(n3063), .Z(n3791) );
  XOR U3920 ( .A(key[234]), .B(n3777), .Z(out[106]) );
  XNOR U3921 ( .A(n3792), .B(n3793), .Z(n3777) );
  XOR U3922 ( .A(n3794), .B(n3060), .Z(out[105]) );
  XNOR U3923 ( .A(n3783), .B(n3795), .Z(n3782) );
  XNOR U3924 ( .A(n3796), .B(n3797), .Z(n3795) );
  NANDN U3925 ( .A(n3798), .B(n3770), .Z(n3797) );
  XNOR U3926 ( .A(n3765), .B(n3799), .Z(n3783) );
  XNOR U3927 ( .A(n3800), .B(n3801), .Z(n3799) );
  NANDN U3928 ( .A(n3802), .B(n3803), .Z(n3801) );
  XOR U3929 ( .A(n3793), .B(n3790), .Z(n3066) );
  XNOR U3930 ( .A(n3765), .B(n3804), .Z(n3790) );
  XNOR U3931 ( .A(n3796), .B(n3805), .Z(n3804) );
  NANDN U3932 ( .A(n3806), .B(n3807), .Z(n3805) );
  OR U3933 ( .A(n3808), .B(n3809), .Z(n3796) );
  XOR U3934 ( .A(n3810), .B(n3800), .Z(n3765) );
  NANDN U3935 ( .A(n3811), .B(n3812), .Z(n3800) );
  ANDN U3936 ( .B(n3813), .A(n3814), .Z(n3810) );
  XNOR U3937 ( .A(key[233]), .B(n3792), .Z(n3794) );
  IV U3938 ( .A(n3063), .Z(n3792) );
  XOR U3939 ( .A(n3815), .B(n3816), .Z(n3063) );
  XNOR U3940 ( .A(n3817), .B(n3818), .Z(n3816) );
  NANDN U3941 ( .A(n3819), .B(n3775), .Z(n3818) );
  XNOR U3942 ( .A(n3763), .B(n3820), .Z(out[104]) );
  XOR U3943 ( .A(key[232]), .B(n3793), .Z(n3820) );
  XNOR U3944 ( .A(n3815), .B(n3821), .Z(n3793) );
  XOR U3945 ( .A(n3822), .B(n3767), .Z(n3821) );
  OR U3946 ( .A(n3823), .B(n3808), .Z(n3767) );
  XNOR U3947 ( .A(n3770), .B(n3807), .Z(n3808) );
  ANDN U3948 ( .B(n3824), .A(n3825), .Z(n3822) );
  IV U3949 ( .A(n3779), .Z(n3763) );
  XOR U3950 ( .A(n3771), .B(n3826), .Z(n3779) );
  XOR U3951 ( .A(n3827), .B(n3817), .Z(n3826) );
  XNOR U3952 ( .A(n3789), .B(n3775), .Z(n3786) );
  NOR U3953 ( .A(n3829), .B(n3789), .Z(n3827) );
  XNOR U3954 ( .A(n3815), .B(n3830), .Z(n3771) );
  XNOR U3955 ( .A(n3831), .B(n3832), .Z(n3830) );
  NANDN U3956 ( .A(n3802), .B(n3833), .Z(n3832) );
  XOR U3957 ( .A(n3834), .B(n3831), .Z(n3815) );
  OR U3958 ( .A(n3811), .B(n3835), .Z(n3831) );
  XOR U3959 ( .A(n3836), .B(n3802), .Z(n3811) );
  XNOR U3960 ( .A(n3807), .B(n3775), .Z(n3802) );
  XOR U3961 ( .A(n3837), .B(n3838), .Z(n3775) );
  NANDN U3962 ( .A(n3839), .B(n3840), .Z(n3838) );
  IV U3963 ( .A(n3825), .Z(n3807) );
  XNOR U3964 ( .A(n3841), .B(n3842), .Z(n3825) );
  NANDN U3965 ( .A(n3839), .B(n3843), .Z(n3842) );
  ANDN U3966 ( .B(n3836), .A(n3844), .Z(n3834) );
  IV U3967 ( .A(n3814), .Z(n3836) );
  XOR U3968 ( .A(n3789), .B(n3770), .Z(n3814) );
  XNOR U3969 ( .A(n3845), .B(n3841), .Z(n3770) );
  NANDN U3970 ( .A(n3846), .B(n3847), .Z(n3841) );
  XOR U3971 ( .A(n3843), .B(n3848), .Z(n3847) );
  ANDN U3972 ( .B(n3848), .A(n3849), .Z(n3845) );
  XOR U3973 ( .A(n3850), .B(n3837), .Z(n3789) );
  NANDN U3974 ( .A(n3846), .B(n3851), .Z(n3837) );
  XOR U3975 ( .A(n3852), .B(n3840), .Z(n3851) );
  XNOR U3976 ( .A(n3853), .B(n3854), .Z(n3839) );
  XOR U3977 ( .A(n3855), .B(n3856), .Z(n3854) );
  XNOR U3978 ( .A(n3857), .B(n3858), .Z(n3853) );
  XNOR U3979 ( .A(n3859), .B(n3860), .Z(n3858) );
  ANDN U3980 ( .B(n3852), .A(n3856), .Z(n3859) );
  ANDN U3981 ( .B(n3852), .A(n3849), .Z(n3850) );
  XNOR U3982 ( .A(n3855), .B(n3861), .Z(n3849) );
  XOR U3983 ( .A(n3862), .B(n3860), .Z(n3861) );
  NAND U3984 ( .A(n3863), .B(n3864), .Z(n3860) );
  XNOR U3985 ( .A(n3857), .B(n3840), .Z(n3864) );
  IV U3986 ( .A(n3852), .Z(n3857) );
  XNOR U3987 ( .A(n3843), .B(n3856), .Z(n3863) );
  IV U3988 ( .A(n3848), .Z(n3856) );
  XOR U3989 ( .A(n3865), .B(n3866), .Z(n3848) );
  XNOR U3990 ( .A(n3867), .B(n3868), .Z(n3866) );
  XNOR U3991 ( .A(n3869), .B(n3870), .Z(n3865) );
  ANDN U3992 ( .B(n3871), .A(n3829), .Z(n3869) );
  AND U3993 ( .A(n3840), .B(n3843), .Z(n3862) );
  XNOR U3994 ( .A(n3840), .B(n3843), .Z(n3855) );
  XNOR U3995 ( .A(n3872), .B(n3873), .Z(n3843) );
  XNOR U3996 ( .A(n3874), .B(n3868), .Z(n3873) );
  XOR U3997 ( .A(n3875), .B(n3876), .Z(n3872) );
  XNOR U3998 ( .A(n3877), .B(n3870), .Z(n3876) );
  OR U3999 ( .A(n3787), .B(n3828), .Z(n3870) );
  XNOR U4000 ( .A(n3878), .B(n3879), .Z(n3828) );
  XNOR U4001 ( .A(n3788), .B(n3776), .Z(n3787) );
  ANDN U4002 ( .B(n3880), .A(n3819), .Z(n3877) );
  XNOR U4003 ( .A(n3881), .B(n3882), .Z(n3840) );
  XNOR U4004 ( .A(n3868), .B(n3883), .Z(n3882) );
  XOR U4005 ( .A(n3798), .B(n3875), .Z(n3883) );
  XNOR U4006 ( .A(n3878), .B(n3788), .Z(n3868) );
  XNOR U4007 ( .A(n3884), .B(n3885), .Z(n3881) );
  XNOR U4008 ( .A(n3886), .B(n3887), .Z(n3885) );
  ANDN U4009 ( .B(n3824), .A(n3806), .Z(n3886) );
  XNOR U4010 ( .A(n3888), .B(n3889), .Z(n3852) );
  XNOR U4011 ( .A(n3874), .B(n3890), .Z(n3889) );
  XNOR U4012 ( .A(n3806), .B(n3867), .Z(n3890) );
  XOR U4013 ( .A(n3875), .B(n3891), .Z(n3867) );
  XNOR U4014 ( .A(n3892), .B(n3893), .Z(n3891) );
  NAND U4015 ( .A(n3833), .B(n3803), .Z(n3893) );
  XNOR U4016 ( .A(n3894), .B(n3892), .Z(n3875) );
  NANDN U4017 ( .A(n3835), .B(n3812), .Z(n3892) );
  XOR U4018 ( .A(n3813), .B(n3803), .Z(n3812) );
  XNOR U4019 ( .A(n3895), .B(n3776), .Z(n3803) );
  XOR U4020 ( .A(n3844), .B(n3833), .Z(n3835) );
  XOR U4021 ( .A(n3824), .B(n3879), .Z(n3833) );
  ANDN U4022 ( .B(n3813), .A(n3844), .Z(n3894) );
  XNOR U4023 ( .A(n3884), .B(n3878), .Z(n3844) );
  IV U4024 ( .A(n3829), .Z(n3878) );
  XNOR U4025 ( .A(n3896), .B(n3897), .Z(n3829) );
  XOR U4026 ( .A(n3898), .B(n3899), .Z(n3897) );
  XOR U4027 ( .A(n3900), .B(n3871), .Z(n3813) );
  XOR U4028 ( .A(n3879), .B(n3880), .Z(n3874) );
  IV U4029 ( .A(n3776), .Z(n3880) );
  XOR U4030 ( .A(n3901), .B(n3902), .Z(n3776) );
  XNOR U4031 ( .A(n3903), .B(n3899), .Z(n3902) );
  IV U4032 ( .A(n3819), .Z(n3879) );
  XOR U4033 ( .A(n3899), .B(n3904), .Z(n3819) );
  XNOR U4034 ( .A(n3824), .B(n3905), .Z(n3888) );
  XNOR U4035 ( .A(n3906), .B(n3887), .Z(n3905) );
  OR U4036 ( .A(n3809), .B(n3823), .Z(n3887) );
  XNOR U4037 ( .A(n3884), .B(n3824), .Z(n3823) );
  XOR U4038 ( .A(n3798), .B(n3895), .Z(n3809) );
  IV U4039 ( .A(n3806), .Z(n3895) );
  XOR U4040 ( .A(n3871), .B(n3907), .Z(n3806) );
  XOR U4041 ( .A(n3903), .B(n3896), .Z(n3907) );
  XNOR U4042 ( .A(key[170]), .B(\w0[1][42] ), .Z(n3896) );
  XOR U4043 ( .A(n3908), .B(n3909), .Z(\w0[1][42] ) );
  XOR U4044 ( .A(n1029), .B(n377), .Z(n3909) );
  XNOR U4045 ( .A(n1036), .B(n412), .Z(n3908) );
  IV U4046 ( .A(n3788), .Z(n3871) );
  XOR U4047 ( .A(n3901), .B(n3910), .Z(n3788) );
  XNOR U4048 ( .A(n3899), .B(n3911), .Z(n3910) );
  ANDN U4049 ( .B(n3900), .A(n3769), .Z(n3906) );
  IV U4050 ( .A(n3798), .Z(n3900) );
  XOR U4051 ( .A(n3901), .B(n3912), .Z(n3798) );
  XOR U4052 ( .A(n3899), .B(n3913), .Z(n3912) );
  XOR U4053 ( .A(n3769), .B(n3914), .Z(n3899) );
  XOR U4054 ( .A(key[174]), .B(\w0[1][46] ), .Z(n3914) );
  XNOR U4055 ( .A(n3915), .B(n3916), .Z(\w0[1][46] ) );
  XNOR U4056 ( .A(n1011), .B(n386), .Z(n3916) );
  XOR U4057 ( .A(n399), .B(n3917), .Z(n386) );
  XNOR U4058 ( .A(n3918), .B(n3919), .Z(n399) );
  IV U4059 ( .A(n3884), .Z(n3769) );
  IV U4060 ( .A(n3904), .Z(n3901) );
  XOR U4061 ( .A(key[173]), .B(\w0[1][45] ), .Z(n3904) );
  XOR U4062 ( .A(n3920), .B(n3921), .Z(\w0[1][45] ) );
  XOR U4063 ( .A(n1024), .B(n390), .Z(n3921) );
  XOR U4064 ( .A(n1009), .B(n3922), .Z(n390) );
  XNOR U4065 ( .A(n3923), .B(n1005), .Z(n3920) );
  IV U4066 ( .A(n3924), .Z(n1005) );
  XOR U4067 ( .A(n3925), .B(n3926), .Z(n3824) );
  XOR U4068 ( .A(n3913), .B(n3911), .Z(n3926) );
  XOR U4069 ( .A(key[175]), .B(\w0[1][47] ), .Z(n3911) );
  XNOR U4070 ( .A(n396), .B(n3927), .Z(\w0[1][47] ) );
  XOR U4071 ( .A(n1006), .B(n417), .Z(n3927) );
  XOR U4072 ( .A(n3928), .B(n3929), .Z(n417) );
  XOR U4073 ( .A(n1017), .B(n3930), .Z(n396) );
  XNOR U4074 ( .A(key[172]), .B(\w0[1][44] ), .Z(n3913) );
  XOR U4075 ( .A(n3931), .B(n3932), .Z(\w0[1][44] ) );
  XOR U4076 ( .A(n403), .B(n3933), .Z(n3932) );
  XOR U4077 ( .A(n1021), .B(n3934), .Z(n403) );
  XOR U4078 ( .A(n1031), .B(n402), .Z(n3931) );
  XNOR U4079 ( .A(n393), .B(n3929), .Z(n402) );
  XNOR U4080 ( .A(n3884), .B(n3898), .Z(n3925) );
  XOR U4081 ( .A(n3903), .B(n3935), .Z(n3898) );
  XOR U4082 ( .A(key[171]), .B(\w0[1][43] ), .Z(n3935) );
  XOR U4083 ( .A(n3936), .B(n3937), .Z(\w0[1][43] ) );
  XOR U4084 ( .A(n410), .B(n3938), .Z(n3937) );
  XOR U4085 ( .A(n405), .B(n3929), .Z(n410) );
  IV U4086 ( .A(n3919), .Z(n3929) );
  XOR U4087 ( .A(n997), .B(n409), .Z(n3936) );
  IV U4088 ( .A(n3939), .Z(n409) );
  XOR U4089 ( .A(key[169]), .B(\w0[1][41] ), .Z(n3903) );
  XOR U4090 ( .A(n3940), .B(n3941), .Z(\w0[1][41] ) );
  XNOR U4091 ( .A(n1040), .B(n413), .Z(n3941) );
  XOR U4092 ( .A(n3942), .B(n379), .Z(n3940) );
  XOR U4093 ( .A(key[168]), .B(\w0[1][40] ), .Z(n3884) );
  XOR U4094 ( .A(n3943), .B(n3944), .Z(\w0[1][40] ) );
  XNOR U4095 ( .A(n416), .B(n3928), .Z(n3944) );
  XOR U4096 ( .A(n1015), .B(n1034), .Z(n3943) );
  XOR U4097 ( .A(n3945), .B(n3946), .Z(out[103]) );
  XNOR U4098 ( .A(n16), .B(n3947), .Z(n3946) );
  IV U4099 ( .A(n3948), .Z(n16) );
  XNOR U4100 ( .A(n8), .B(n3949), .Z(n3945) );
  XNOR U4101 ( .A(key[231]), .B(n12), .Z(n3949) );
  XNOR U4102 ( .A(n3950), .B(n3951), .Z(n8) );
  XNOR U4103 ( .A(n3952), .B(n3953), .Z(n3951) );
  NANDN U4104 ( .A(n3954), .B(n3955), .Z(n3953) );
  XOR U4105 ( .A(n3948), .B(n3956), .Z(out[102]) );
  XNOR U4106 ( .A(key[230]), .B(n10), .Z(n3956) );
  XNOR U4107 ( .A(n3958), .B(n3959), .Z(n3957) );
  OR U4108 ( .A(n3960), .B(n3961), .Z(n3959) );
  XNOR U4109 ( .A(n3962), .B(n3963), .Z(n3950) );
  XNOR U4110 ( .A(n3964), .B(n3965), .Z(n3963) );
  NAND U4111 ( .A(n3966), .B(n3967), .Z(n3965) );
  XNOR U4112 ( .A(n9), .B(n19), .Z(n3948) );
  XNOR U4113 ( .A(n3962), .B(n3968), .Z(n9) );
  XNOR U4114 ( .A(n3952), .B(n3969), .Z(n3968) );
  NANDN U4115 ( .A(n3970), .B(n3971), .Z(n3969) );
  OR U4116 ( .A(n3972), .B(n3973), .Z(n3952) );
  XOR U4117 ( .A(n3974), .B(n3975), .Z(out[101]) );
  XNOR U4118 ( .A(n3947), .B(n3976), .Z(n3975) );
  XOR U4119 ( .A(n3962), .B(n17), .Z(n3976) );
  XOR U4120 ( .A(n3977), .B(n3964), .Z(n3962) );
  NANDN U4121 ( .A(n3978), .B(n3979), .Z(n3964) );
  ANDN U4122 ( .B(n3980), .A(n3981), .Z(n3977) );
  XNOR U4123 ( .A(n3982), .B(n3983), .Z(n3947) );
  XNOR U4124 ( .A(n3984), .B(n3985), .Z(n3983) );
  NANDN U4125 ( .A(n3986), .B(n3955), .Z(n3985) );
  XOR U4126 ( .A(n3987), .B(n3988), .Z(n3974) );
  XNOR U4127 ( .A(key[229]), .B(n3958), .Z(n3988) );
  NANDN U4128 ( .A(n3989), .B(n3990), .Z(n3958) );
  ANDN U4129 ( .B(n3991), .A(n3992), .Z(n3987) );
  XOR U4130 ( .A(n17), .B(n3993), .Z(out[100]) );
  XNOR U4131 ( .A(key[228]), .B(n13), .Z(n3993) );
  XOR U4132 ( .A(n3994), .B(n3995), .Z(n19) );
  XOR U4133 ( .A(n3996), .B(n3984), .Z(n3995) );
  OR U4134 ( .A(n3972), .B(n3997), .Z(n3984) );
  XNOR U4135 ( .A(n3955), .B(n3971), .Z(n3972) );
  ANDN U4136 ( .B(n3998), .A(n3999), .Z(n3996) );
  XNOR U4137 ( .A(n3994), .B(n4000), .Z(n12) );
  XNOR U4138 ( .A(n4001), .B(n4002), .Z(n4000) );
  NAND U4139 ( .A(n3991), .B(n4003), .Z(n4002) );
  XOR U4140 ( .A(n3982), .B(n4004), .Z(n17) );
  XOR U4141 ( .A(n4005), .B(n4001), .Z(n4004) );
  NANDN U4142 ( .A(n4006), .B(n3990), .Z(n4001) );
  XNOR U4143 ( .A(n3960), .B(n3991), .Z(n3990) );
  NOR U4144 ( .A(n4007), .B(n3960), .Z(n4005) );
  XNOR U4145 ( .A(n3994), .B(n4008), .Z(n3982) );
  XNOR U4146 ( .A(n4009), .B(n4010), .Z(n4008) );
  NAND U4147 ( .A(n3967), .B(n4011), .Z(n4010) );
  XOR U4148 ( .A(n4012), .B(n4009), .Z(n3994) );
  OR U4149 ( .A(n3978), .B(n4013), .Z(n4009) );
  XOR U4150 ( .A(n3981), .B(n3967), .Z(n3978) );
  XOR U4151 ( .A(n3971), .B(n3991), .Z(n3967) );
  XOR U4152 ( .A(n4014), .B(n4015), .Z(n3991) );
  NANDN U4153 ( .A(n4016), .B(n4017), .Z(n4015) );
  IV U4154 ( .A(n3999), .Z(n3971) );
  XNOR U4155 ( .A(n4018), .B(n4019), .Z(n3999) );
  NANDN U4156 ( .A(n4016), .B(n4020), .Z(n4019) );
  NOR U4157 ( .A(n3981), .B(n4021), .Z(n4012) );
  XOR U4158 ( .A(n3960), .B(n3955), .Z(n3981) );
  XNOR U4159 ( .A(n4022), .B(n4018), .Z(n3955) );
  NANDN U4160 ( .A(n4023), .B(n4024), .Z(n4018) );
  XOR U4161 ( .A(n4020), .B(n4025), .Z(n4024) );
  ANDN U4162 ( .B(n4025), .A(n4026), .Z(n4022) );
  XOR U4163 ( .A(n4027), .B(n4014), .Z(n3960) );
  NANDN U4164 ( .A(n4023), .B(n4028), .Z(n4014) );
  XOR U4165 ( .A(n4029), .B(n4017), .Z(n4028) );
  XNOR U4166 ( .A(n4030), .B(n4031), .Z(n4016) );
  XOR U4167 ( .A(n4032), .B(n4033), .Z(n4031) );
  XNOR U4168 ( .A(n4034), .B(n4035), .Z(n4030) );
  XNOR U4169 ( .A(n4036), .B(n4037), .Z(n4035) );
  ANDN U4170 ( .B(n4029), .A(n4033), .Z(n4036) );
  ANDN U4171 ( .B(n4029), .A(n4026), .Z(n4027) );
  XNOR U4172 ( .A(n4032), .B(n4038), .Z(n4026) );
  XOR U4173 ( .A(n4039), .B(n4037), .Z(n4038) );
  NAND U4174 ( .A(n4040), .B(n4041), .Z(n4037) );
  XNOR U4175 ( .A(n4034), .B(n4017), .Z(n4041) );
  IV U4176 ( .A(n4029), .Z(n4034) );
  XNOR U4177 ( .A(n4020), .B(n4033), .Z(n4040) );
  IV U4178 ( .A(n4025), .Z(n4033) );
  XOR U4179 ( .A(n4042), .B(n4043), .Z(n4025) );
  XNOR U4180 ( .A(n4044), .B(n4045), .Z(n4043) );
  XNOR U4181 ( .A(n4046), .B(n4047), .Z(n4042) );
  ANDN U4182 ( .B(n4048), .A(n4007), .Z(n4046) );
  AND U4183 ( .A(n4017), .B(n4020), .Z(n4039) );
  XNOR U4184 ( .A(n4017), .B(n4020), .Z(n4032) );
  XNOR U4185 ( .A(n4049), .B(n4050), .Z(n4020) );
  XOR U4186 ( .A(n4051), .B(n4045), .Z(n4050) );
  XNOR U4187 ( .A(n4052), .B(n4053), .Z(n4049) );
  XNOR U4188 ( .A(n4054), .B(n4047), .Z(n4053) );
  OR U4189 ( .A(n3989), .B(n4006), .Z(n4047) );
  XNOR U4190 ( .A(n4055), .B(n4003), .Z(n4006) );
  XNOR U4191 ( .A(n3992), .B(n3961), .Z(n3989) );
  ANDN U4192 ( .B(n4003), .A(n3992), .Z(n4054) );
  XNOR U4193 ( .A(n4056), .B(n4057), .Z(n4017) );
  XNOR U4194 ( .A(n4045), .B(n4058), .Z(n4057) );
  XOR U4195 ( .A(n3954), .B(n4051), .Z(n4058) );
  XNOR U4196 ( .A(n4055), .B(n3961), .Z(n4045) );
  XNOR U4197 ( .A(n4059), .B(n4060), .Z(n4056) );
  XNOR U4198 ( .A(n4061), .B(n4062), .Z(n4060) );
  ANDN U4199 ( .B(n3998), .A(n3970), .Z(n4061) );
  XNOR U4200 ( .A(n4063), .B(n4064), .Z(n4029) );
  XNOR U4201 ( .A(n4044), .B(n4065), .Z(n4064) );
  XNOR U4202 ( .A(n4052), .B(n3970), .Z(n4065) );
  XOR U4203 ( .A(n4003), .B(n4066), .Z(n4052) );
  XOR U4204 ( .A(n4051), .B(n4067), .Z(n4044) );
  XNOR U4205 ( .A(n4068), .B(n4069), .Z(n4067) );
  NAND U4206 ( .A(n4011), .B(n3966), .Z(n4069) );
  XNOR U4207 ( .A(n4070), .B(n4068), .Z(n4051) );
  NANDN U4208 ( .A(n4013), .B(n3979), .Z(n4068) );
  XOR U4209 ( .A(n3980), .B(n3966), .Z(n3979) );
  XNOR U4210 ( .A(n4066), .B(n3970), .Z(n3966) );
  IV U4211 ( .A(n3992), .Z(n4066) );
  XOR U4212 ( .A(n4071), .B(n4072), .Z(n3992) );
  XOR U4213 ( .A(n4073), .B(n4074), .Z(n4072) );
  XOR U4214 ( .A(n4021), .B(n4011), .Z(n4013) );
  XOR U4215 ( .A(n4003), .B(n3998), .Z(n4011) );
  ANDN U4216 ( .B(n3980), .A(n4021), .Z(n4070) );
  XNOR U4217 ( .A(n4059), .B(n4055), .Z(n4021) );
  IV U4218 ( .A(n4007), .Z(n4055) );
  XOR U4219 ( .A(n4075), .B(n4076), .Z(n4007) );
  XOR U4220 ( .A(n4077), .B(n4073), .Z(n4076) );
  XOR U4221 ( .A(n4078), .B(n4048), .Z(n3980) );
  XNOR U4222 ( .A(n3998), .B(n4079), .Z(n4063) );
  XNOR U4223 ( .A(n4080), .B(n4062), .Z(n4079) );
  OR U4224 ( .A(n3973), .B(n3997), .Z(n4062) );
  XNOR U4225 ( .A(n4059), .B(n3998), .Z(n3997) );
  XNOR U4226 ( .A(n3954), .B(n3970), .Z(n3973) );
  XOR U4227 ( .A(n4048), .B(n4081), .Z(n3970) );
  XNOR U4228 ( .A(n4077), .B(n4074), .Z(n4081) );
  XOR U4229 ( .A(key[130]), .B(\w0[1][2] ), .Z(n4077) );
  XOR U4230 ( .A(n612), .B(n4082), .Z(\w0[1][2] ) );
  XNOR U4231 ( .A(n1824), .B(n1232), .Z(n4082) );
  XNOR U4232 ( .A(n4083), .B(n626), .Z(n1232) );
  IV U4233 ( .A(n1231), .Z(n612) );
  XNOR U4234 ( .A(n1797), .B(n624), .Z(n1231) );
  XOR U4235 ( .A(n4084), .B(n4085), .Z(n624) );
  XNOR U4236 ( .A(n4086), .B(n4087), .Z(n4085) );
  XNOR U4237 ( .A(n4088), .B(n4089), .Z(n4084) );
  IV U4238 ( .A(n3961), .Z(n4048) );
  XNOR U4239 ( .A(n4090), .B(n4003), .Z(n3961) );
  IV U4240 ( .A(n4078), .Z(n3954) );
  ANDN U4241 ( .B(n4078), .A(n3986), .Z(n4080) );
  XOR U4242 ( .A(n4091), .B(n4003), .Z(n4078) );
  XNOR U4243 ( .A(n4073), .B(n4071), .Z(n4003) );
  XNOR U4244 ( .A(key[133]), .B(\w0[1][5] ), .Z(n4071) );
  XNOR U4245 ( .A(n1209), .B(n4092), .Z(\w0[1][5] ) );
  XNOR U4246 ( .A(n1204), .B(n1808), .Z(n4092) );
  XNOR U4247 ( .A(n1208), .B(n593), .Z(n1808) );
  XNOR U4248 ( .A(n4093), .B(n4094), .Z(n593) );
  XNOR U4249 ( .A(n4095), .B(n4096), .Z(n4094) );
  XNOR U4250 ( .A(n4097), .B(n4098), .Z(n4093) );
  XOR U4251 ( .A(n4099), .B(n4100), .Z(n4098) );
  ANDN U4252 ( .B(n4101), .A(n4102), .Z(n4100) );
  IV U4253 ( .A(n1225), .Z(n1208) );
  XOR U4254 ( .A(n4103), .B(n4104), .Z(n1225) );
  XNOR U4255 ( .A(n4105), .B(n4106), .Z(n4104) );
  XNOR U4256 ( .A(n4107), .B(n4108), .Z(n4103) );
  XNOR U4257 ( .A(n4109), .B(n4110), .Z(n4108) );
  ANDN U4258 ( .B(n4111), .A(n4112), .Z(n4110) );
  XOR U4259 ( .A(n1809), .B(n596), .Z(n1204) );
  XOR U4260 ( .A(n4113), .B(n4087), .Z(n596) );
  XNOR U4261 ( .A(n4114), .B(n4115), .Z(n4087) );
  XNOR U4262 ( .A(n4116), .B(n4117), .Z(n4115) );
  ANDN U4263 ( .B(n4118), .A(n4119), .Z(n4116) );
  XNOR U4264 ( .A(n3986), .B(n4120), .Z(n4073) );
  XOR U4265 ( .A(key[134]), .B(\w0[1][6] ), .Z(n4120) );
  XNOR U4266 ( .A(n1809), .B(n4121), .Z(\w0[1][6] ) );
  XOR U4267 ( .A(n601), .B(n1804), .Z(n4121) );
  XOR U4268 ( .A(n4122), .B(n1207), .Z(n1804) );
  XNOR U4269 ( .A(n602), .B(n595), .Z(n1207) );
  XNOR U4270 ( .A(n4123), .B(n4124), .Z(n595) );
  XOR U4271 ( .A(n4125), .B(n4126), .Z(n602) );
  XOR U4272 ( .A(n605), .B(n1218), .Z(n601) );
  XOR U4273 ( .A(n4127), .B(n4128), .Z(n1218) );
  XNOR U4274 ( .A(n4113), .B(n4129), .Z(n4128) );
  XOR U4275 ( .A(n4130), .B(n4089), .Z(n4127) );
  XOR U4276 ( .A(n4131), .B(n4132), .Z(n1809) );
  IV U4277 ( .A(n4059), .Z(n3986) );
  XOR U4278 ( .A(n4133), .B(n4134), .Z(n3998) );
  XNOR U4279 ( .A(n4091), .B(n4090), .Z(n4134) );
  XOR U4280 ( .A(key[135]), .B(\w0[1][7] ), .Z(n4090) );
  XNOR U4281 ( .A(n4122), .B(n4135), .Z(\w0[1][7] ) );
  XNOR U4282 ( .A(n605), .B(n1813), .Z(n4135) );
  XNOR U4283 ( .A(n589), .B(n1215), .Z(n1813) );
  XOR U4284 ( .A(n4136), .B(n4137), .Z(n1215) );
  XNOR U4285 ( .A(n4138), .B(n4105), .Z(n4137) );
  XNOR U4286 ( .A(n4139), .B(n4140), .Z(n4105) );
  XNOR U4287 ( .A(n4141), .B(n4142), .Z(n4140) );
  OR U4288 ( .A(n4143), .B(n4144), .Z(n4142) );
  XNOR U4289 ( .A(n4145), .B(n4123), .Z(n4136) );
  XNOR U4290 ( .A(n4146), .B(n4147), .Z(n589) );
  XNOR U4291 ( .A(n4125), .B(n4096), .Z(n4147) );
  XNOR U4292 ( .A(n4148), .B(n4149), .Z(n4096) );
  XNOR U4293 ( .A(n4150), .B(n4151), .Z(n4149) );
  NANDN U4294 ( .A(n4152), .B(n4153), .Z(n4151) );
  XOR U4295 ( .A(n1235), .B(n1217), .Z(n4122) );
  XOR U4296 ( .A(n4154), .B(n4155), .Z(n1217) );
  XNOR U4297 ( .A(n4131), .B(n4156), .Z(n4155) );
  XOR U4298 ( .A(key[132]), .B(\w0[1][4] ), .Z(n4091) );
  XOR U4299 ( .A(n4157), .B(n4158), .Z(\w0[1][4] ) );
  XOR U4300 ( .A(n4159), .B(n1817), .Z(n4158) );
  XOR U4301 ( .A(n1220), .B(n581), .Z(n1817) );
  XNOR U4302 ( .A(n4095), .B(n626), .Z(n581) );
  XOR U4303 ( .A(n4160), .B(n4161), .Z(n626) );
  XNOR U4304 ( .A(n621), .B(n4106), .Z(n1220) );
  IV U4305 ( .A(n4083), .Z(n621) );
  XOR U4306 ( .A(n4162), .B(n4163), .Z(n4083) );
  XOR U4307 ( .A(n580), .B(n1816), .Z(n4157) );
  XNOR U4308 ( .A(n4164), .B(n1209), .Z(n1816) );
  XOR U4309 ( .A(n4165), .B(n4166), .Z(n1209) );
  XNOR U4310 ( .A(n4167), .B(n4156), .Z(n4166) );
  XNOR U4311 ( .A(n4168), .B(n4169), .Z(n4156) );
  XNOR U4312 ( .A(n4170), .B(n4171), .Z(n4169) );
  NANDN U4313 ( .A(n4172), .B(n4173), .Z(n4171) );
  XNOR U4314 ( .A(n4174), .B(n4175), .Z(n4165) );
  XOR U4315 ( .A(n4176), .B(n4177), .Z(n4175) );
  ANDN U4316 ( .B(n4178), .A(n4179), .Z(n4177) );
  XNOR U4317 ( .A(n605), .B(n1210), .Z(n580) );
  XNOR U4318 ( .A(n4180), .B(n4181), .Z(n1210) );
  XOR U4319 ( .A(n4182), .B(n4129), .Z(n4181) );
  XNOR U4320 ( .A(n4183), .B(n4184), .Z(n4129) );
  XNOR U4321 ( .A(n4185), .B(n4186), .Z(n4184) );
  NANDN U4322 ( .A(n4187), .B(n4188), .Z(n4186) );
  XNOR U4323 ( .A(n4189), .B(n4190), .Z(n4180) );
  XOR U4324 ( .A(n4117), .B(n4191), .Z(n4190) );
  ANDN U4325 ( .B(n4192), .A(n4193), .Z(n4191) );
  NOR U4326 ( .A(n4194), .B(n4195), .Z(n4117) );
  XOR U4327 ( .A(n4059), .B(n4075), .Z(n4133) );
  XNOR U4328 ( .A(n4074), .B(n4196), .Z(n4075) );
  XOR U4329 ( .A(key[131]), .B(\w0[1][3] ), .Z(n4196) );
  XOR U4330 ( .A(n4197), .B(n4198), .Z(\w0[1][3] ) );
  XNOR U4331 ( .A(n1797), .B(n1196), .Z(n4198) );
  XNOR U4332 ( .A(n615), .B(n627), .Z(n1196) );
  XOR U4333 ( .A(n4199), .B(n4200), .Z(n627) );
  XNOR U4334 ( .A(n4201), .B(n4124), .Z(n4200) );
  XNOR U4335 ( .A(n4202), .B(n4203), .Z(n4124) );
  XOR U4336 ( .A(n4204), .B(n4109), .Z(n4203) );
  OR U4337 ( .A(n4205), .B(n4206), .Z(n4109) );
  ANDN U4338 ( .B(n4207), .A(n4208), .Z(n4204) );
  XNOR U4339 ( .A(n4162), .B(n4209), .Z(n4199) );
  IV U4340 ( .A(n4145), .Z(n4162) );
  XOR U4341 ( .A(n4146), .B(n4210), .Z(n615) );
  XOR U4342 ( .A(n4211), .B(n4126), .Z(n4210) );
  XOR U4343 ( .A(n4212), .B(n4213), .Z(n4126) );
  XNOR U4344 ( .A(n4214), .B(n4099), .Z(n4213) );
  NOR U4345 ( .A(n4215), .B(n4216), .Z(n4099) );
  ANDN U4346 ( .B(n4217), .A(n4218), .Z(n4214) );
  XNOR U4347 ( .A(n4219), .B(n4220), .Z(n4146) );
  XOR U4348 ( .A(n4154), .B(n4221), .Z(n1797) );
  XOR U4349 ( .A(n4222), .B(n4132), .Z(n4221) );
  XOR U4350 ( .A(n4223), .B(n4224), .Z(n4132) );
  XNOR U4351 ( .A(n4225), .B(n4176), .Z(n4224) );
  NOR U4352 ( .A(n4226), .B(n4227), .Z(n4176) );
  ANDN U4353 ( .B(n4228), .A(n4229), .Z(n4225) );
  XNOR U4354 ( .A(n4230), .B(n4231), .Z(n4154) );
  XNOR U4355 ( .A(n614), .B(n1821), .Z(n4197) );
  XNOR U4356 ( .A(n4164), .B(n4159), .Z(n1821) );
  IV U4357 ( .A(n1226), .Z(n4159) );
  XNOR U4358 ( .A(n4167), .B(n1824), .Z(n1226) );
  XOR U4359 ( .A(n605), .B(n1224), .Z(n614) );
  XOR U4360 ( .A(n619), .B(n4182), .Z(n1224) );
  XOR U4361 ( .A(n4232), .B(n4182), .Z(n605) );
  XOR U4362 ( .A(n4183), .B(n4233), .Z(n4182) );
  XOR U4363 ( .A(n4234), .B(n4235), .Z(n4233) );
  NOR U4364 ( .A(n4236), .B(n4119), .Z(n4234) );
  XNOR U4365 ( .A(n4237), .B(n4238), .Z(n4183) );
  XNOR U4366 ( .A(n4239), .B(n4240), .Z(n4238) );
  NANDN U4367 ( .A(n4241), .B(n4242), .Z(n4240) );
  XOR U4368 ( .A(key[129]), .B(\w0[1][1] ), .Z(n4074) );
  XNOR U4369 ( .A(n625), .B(n4243), .Z(\w0[1][1] ) );
  XOR U4370 ( .A(n4244), .B(n1236), .Z(n4243) );
  XOR U4371 ( .A(n618), .B(n606), .Z(n1236) );
  XNOR U4372 ( .A(n4201), .B(n4245), .Z(n606) );
  XOR U4373 ( .A(n4145), .B(n4123), .Z(n4245) );
  XOR U4374 ( .A(n4163), .B(n4209), .Z(n4123) );
  XNOR U4375 ( .A(n4107), .B(n4246), .Z(n4209) );
  XNOR U4376 ( .A(n4247), .B(n4248), .Z(n4246) );
  NANDN U4377 ( .A(n4249), .B(n4250), .Z(n4248) );
  XNOR U4378 ( .A(n4251), .B(n4252), .Z(n4145) );
  XNOR U4379 ( .A(n4253), .B(n4254), .Z(n4252) );
  NANDN U4380 ( .A(n4255), .B(n4111), .Z(n4254) );
  IV U4381 ( .A(n4138), .Z(n4201) );
  XOR U4382 ( .A(n4202), .B(n4256), .Z(n4138) );
  XNOR U4383 ( .A(n4247), .B(n4257), .Z(n4256) );
  OR U4384 ( .A(n4143), .B(n4258), .Z(n4257) );
  OR U4385 ( .A(n4259), .B(n4260), .Z(n4247) );
  XOR U4386 ( .A(n4107), .B(n4261), .Z(n4202) );
  XNOR U4387 ( .A(n4262), .B(n4263), .Z(n4261) );
  NANDN U4388 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U4389 ( .A(n4266), .B(n4262), .Z(n4107) );
  NANDN U4390 ( .A(n4267), .B(n4268), .Z(n4262) );
  AND U4391 ( .A(n4269), .B(n4270), .Z(n4266) );
  XNOR U4392 ( .A(n4125), .B(n4271), .Z(n618) );
  XOR U4393 ( .A(n4219), .B(n4220), .Z(n4271) );
  XOR U4394 ( .A(n4212), .B(n4272), .Z(n4220) );
  XNOR U4395 ( .A(n4273), .B(n4274), .Z(n4272) );
  NANDN U4396 ( .A(n4152), .B(n4275), .Z(n4274) );
  XNOR U4397 ( .A(n4097), .B(n4276), .Z(n4212) );
  XNOR U4398 ( .A(n4277), .B(n4278), .Z(n4276) );
  NANDN U4399 ( .A(n4279), .B(n4280), .Z(n4278) );
  IV U4400 ( .A(n4160), .Z(n4219) );
  XOR U4401 ( .A(n4281), .B(n4282), .Z(n4160) );
  XNOR U4402 ( .A(n4283), .B(n4284), .Z(n4282) );
  NANDN U4403 ( .A(n4285), .B(n4286), .Z(n4284) );
  XOR U4404 ( .A(n4161), .B(n4211), .Z(n4125) );
  XNOR U4405 ( .A(n4097), .B(n4287), .Z(n4211) );
  XNOR U4406 ( .A(n4273), .B(n4288), .Z(n4287) );
  OR U4407 ( .A(n4289), .B(n4290), .Z(n4288) );
  OR U4408 ( .A(n4291), .B(n4292), .Z(n4273) );
  XOR U4409 ( .A(n4293), .B(n4277), .Z(n4097) );
  NANDN U4410 ( .A(n4294), .B(n4295), .Z(n4277) );
  AND U4411 ( .A(n4296), .B(n4297), .Z(n4293) );
  XNOR U4412 ( .A(n619), .B(n1824), .Z(n625) );
  XOR U4413 ( .A(n4298), .B(n4299), .Z(n1824) );
  XOR U4414 ( .A(n4130), .B(n4232), .Z(n619) );
  XOR U4415 ( .A(key[128]), .B(\w0[1][0] ), .Z(n4059) );
  XOR U4416 ( .A(n1216), .B(n4300), .Z(\w0[1][0] ) );
  XNOR U4417 ( .A(n620), .B(n608), .Z(n4300) );
  XNOR U4418 ( .A(n1214), .B(n1235), .Z(n608) );
  IV U4419 ( .A(n4164), .Z(n1235) );
  XOR U4420 ( .A(n4299), .B(n4167), .Z(n4164) );
  XNOR U4421 ( .A(n4168), .B(n4301), .Z(n4167) );
  XOR U4422 ( .A(n4302), .B(n4303), .Z(n4301) );
  NOR U4423 ( .A(n4304), .B(n4229), .Z(n4302) );
  XNOR U4424 ( .A(n4305), .B(n4306), .Z(n4168) );
  XNOR U4425 ( .A(n4307), .B(n4308), .Z(n4306) );
  NANDN U4426 ( .A(n4309), .B(n4310), .Z(n4308) );
  IV U4427 ( .A(n1805), .Z(n1214) );
  XOR U4428 ( .A(n4161), .B(n4095), .Z(n1805) );
  XNOR U4429 ( .A(n4148), .B(n4311), .Z(n4095) );
  XOR U4430 ( .A(n4312), .B(n4283), .Z(n4311) );
  OR U4431 ( .A(n4313), .B(n4215), .Z(n4283) );
  XOR U4432 ( .A(n4218), .B(n4286), .Z(n4215) );
  NOR U4433 ( .A(n4314), .B(n4218), .Z(n4312) );
  XNOR U4434 ( .A(n4281), .B(n4315), .Z(n4148) );
  XNOR U4435 ( .A(n4316), .B(n4317), .Z(n4315) );
  NANDN U4436 ( .A(n4279), .B(n4318), .Z(n4317) );
  XOR U4437 ( .A(n4281), .B(n4319), .Z(n4161) );
  XOR U4438 ( .A(n4320), .B(n4150), .Z(n4319) );
  OR U4439 ( .A(n4321), .B(n4291), .Z(n4150) );
  XNOR U4440 ( .A(n4152), .B(n4289), .Z(n4291) );
  NOR U4441 ( .A(n4322), .B(n4289), .Z(n4320) );
  XOR U4442 ( .A(n4323), .B(n4316), .Z(n4281) );
  OR U4443 ( .A(n4294), .B(n4324), .Z(n4316) );
  XOR U4444 ( .A(n4289), .B(n4286), .Z(n4279) );
  IV U4445 ( .A(n4102), .Z(n4286) );
  XNOR U4446 ( .A(n4325), .B(n4326), .Z(n4102) );
  NANDN U4447 ( .A(n4327), .B(n4328), .Z(n4326) );
  XNOR U4448 ( .A(n4329), .B(n4330), .Z(n4289) );
  NANDN U4449 ( .A(n4327), .B(n4331), .Z(n4330) );
  ANDN U4450 ( .B(n4296), .A(n4332), .Z(n4323) );
  XOR U4451 ( .A(n4152), .B(n4218), .Z(n4296) );
  XOR U4452 ( .A(n4333), .B(n4325), .Z(n4218) );
  NANDN U4453 ( .A(n4334), .B(n4335), .Z(n4325) );
  XOR U4454 ( .A(n4328), .B(n4336), .Z(n4335) );
  ANDN U4455 ( .B(n4336), .A(n4337), .Z(n4333) );
  NANDN U4456 ( .A(n4334), .B(n4339), .Z(n4329) );
  XOR U4457 ( .A(n4340), .B(n4341), .Z(n4327) );
  XOR U4458 ( .A(n4342), .B(n4343), .Z(n4341) );
  XNOR U4459 ( .A(n4344), .B(n4345), .Z(n4340) );
  XNOR U4460 ( .A(n4346), .B(n4347), .Z(n4345) );
  ANDN U4461 ( .B(n4343), .A(n4342), .Z(n4346) );
  ANDN U4462 ( .B(n4343), .A(n4337), .Z(n4338) );
  XNOR U4463 ( .A(n4344), .B(n4348), .Z(n4337) );
  XOR U4464 ( .A(n4349), .B(n4347), .Z(n4348) );
  NAND U4465 ( .A(n4339), .B(n4350), .Z(n4347) );
  XNOR U4466 ( .A(n4328), .B(n4342), .Z(n4350) );
  IV U4467 ( .A(n4336), .Z(n4342) );
  XNOR U4468 ( .A(n4351), .B(n4352), .Z(n4336) );
  XNOR U4469 ( .A(n4353), .B(n4354), .Z(n4352) );
  XOR U4470 ( .A(n4290), .B(n4355), .Z(n4354) );
  XNOR U4471 ( .A(n4322), .B(n4356), .Z(n4351) );
  XNOR U4472 ( .A(n4357), .B(n4358), .Z(n4356) );
  AND U4473 ( .A(n4275), .B(n4153), .Z(n4357) );
  XOR U4474 ( .A(n4331), .B(n4343), .Z(n4339) );
  AND U4475 ( .A(n4328), .B(n4331), .Z(n4349) );
  XNOR U4476 ( .A(n4328), .B(n4331), .Z(n4344) );
  XNOR U4477 ( .A(n4359), .B(n4360), .Z(n4331) );
  XNOR U4478 ( .A(n4361), .B(n4355), .Z(n4360) );
  XOR U4479 ( .A(n4362), .B(n4363), .Z(n4359) );
  XNOR U4480 ( .A(n4364), .B(n4365), .Z(n4363) );
  ANDN U4481 ( .B(n4101), .A(n4285), .Z(n4364) );
  XNOR U4482 ( .A(n4366), .B(n4367), .Z(n4328) );
  XNOR U4483 ( .A(n4275), .B(n4362), .Z(n4368) );
  XOR U4484 ( .A(n4153), .B(n4369), .Z(n4366) );
  XNOR U4485 ( .A(n4370), .B(n4358), .Z(n4369) );
  OR U4486 ( .A(n4292), .B(n4321), .Z(n4358) );
  XOR U4487 ( .A(n4153), .B(n4322), .Z(n4321) );
  XNOR U4488 ( .A(n4275), .B(n4371), .Z(n4292) );
  ANDN U4489 ( .B(n4372), .A(n4290), .Z(n4370) );
  XNOR U4490 ( .A(n4373), .B(n4374), .Z(n4343) );
  XOR U4491 ( .A(n4361), .B(n4353), .Z(n4374) );
  XOR U4492 ( .A(n4362), .B(n4375), .Z(n4353) );
  XNOR U4493 ( .A(n4376), .B(n4377), .Z(n4375) );
  NAND U4494 ( .A(n4318), .B(n4280), .Z(n4377) );
  XNOR U4495 ( .A(n4378), .B(n4376), .Z(n4362) );
  NANDN U4496 ( .A(n4324), .B(n4295), .Z(n4376) );
  XOR U4497 ( .A(n4297), .B(n4280), .Z(n4295) );
  XOR U4498 ( .A(n4371), .B(n4101), .Z(n4280) );
  IV U4499 ( .A(n4290), .Z(n4371) );
  XOR U4500 ( .A(n4217), .B(n4379), .Z(n4290) );
  XNOR U4501 ( .A(n4380), .B(n4381), .Z(n4379) );
  XOR U4502 ( .A(n4332), .B(n4318), .Z(n4324) );
  XNOR U4503 ( .A(n4372), .B(n4285), .Z(n4318) );
  IV U4504 ( .A(n4322), .Z(n4372) );
  XOR U4505 ( .A(n4382), .B(n4383), .Z(n4322) );
  XOR U4506 ( .A(n4384), .B(n4385), .Z(n4383) );
  XNOR U4507 ( .A(n4153), .B(n4386), .Z(n4382) );
  ANDN U4508 ( .B(n4297), .A(n4332), .Z(n4378) );
  XNOR U4509 ( .A(n4153), .B(n4387), .Z(n4332) );
  XOR U4510 ( .A(n4275), .B(n4217), .Z(n4297) );
  XOR U4511 ( .A(n4388), .B(n4389), .Z(n4275) );
  XOR U4512 ( .A(n4390), .B(n4385), .Z(n4389) );
  XOR U4513 ( .A(state[116]), .B(key[116]), .Z(n4385) );
  XOR U4514 ( .A(n4387), .B(n4217), .Z(n4361) );
  IV U4515 ( .A(n4314), .Z(n4387) );
  XNOR U4516 ( .A(n4391), .B(n4365), .Z(n4373) );
  OR U4517 ( .A(n4216), .B(n4313), .Z(n4365) );
  XNOR U4518 ( .A(n4314), .B(n4285), .Z(n4313) );
  XOR U4519 ( .A(n4392), .B(n4388), .Z(n4285) );
  XNOR U4520 ( .A(n4217), .B(n4101), .Z(n4216) );
  XOR U4521 ( .A(n4388), .B(n4393), .Z(n4101) );
  XOR U4522 ( .A(n4380), .B(n4392), .Z(n4393) );
  ANDN U4523 ( .B(n4217), .A(n4314), .Z(n4391) );
  XNOR U4524 ( .A(n4381), .B(n4394), .Z(n4314) );
  XOR U4525 ( .A(n4386), .B(n4392), .Z(n4394) );
  IV U4526 ( .A(n4390), .Z(n4392) );
  XNOR U4527 ( .A(n4380), .B(n4395), .Z(n4386) );
  XNOR U4528 ( .A(state[115]), .B(key[115]), .Z(n4395) );
  XNOR U4529 ( .A(state[113]), .B(key[113]), .Z(n4380) );
  XNOR U4530 ( .A(state[114]), .B(key[114]), .Z(n4381) );
  XOR U4531 ( .A(n4388), .B(n4396), .Z(n4217) );
  XNOR U4532 ( .A(n4390), .B(n4384), .Z(n4396) );
  XNOR U4533 ( .A(state[119]), .B(key[119]), .Z(n4384) );
  XOR U4534 ( .A(n4153), .B(n4397), .Z(n4390) );
  XNOR U4535 ( .A(state[118]), .B(key[118]), .Z(n4397) );
  XOR U4536 ( .A(state[112]), .B(key[112]), .Z(n4153) );
  XNOR U4537 ( .A(state[117]), .B(key[117]), .Z(n4388) );
  XNOR U4538 ( .A(n4244), .B(n607), .Z(n620) );
  XOR U4539 ( .A(n4113), .B(n4398), .Z(n607) );
  XOR U4540 ( .A(n4088), .B(n4089), .Z(n4398) );
  XOR U4541 ( .A(n4114), .B(n4399), .Z(n4089) );
  XNOR U4542 ( .A(n4400), .B(n4401), .Z(n4399) );
  NANDN U4543 ( .A(n4187), .B(n4402), .Z(n4401) );
  XNOR U4544 ( .A(n4189), .B(n4403), .Z(n4114) );
  XNOR U4545 ( .A(n4404), .B(n4405), .Z(n4403) );
  NANDN U4546 ( .A(n4241), .B(n4406), .Z(n4405) );
  IV U4547 ( .A(n4130), .Z(n4088) );
  XOR U4548 ( .A(n4237), .B(n4407), .Z(n4130) );
  XNOR U4549 ( .A(n4235), .B(n4408), .Z(n4407) );
  NANDN U4550 ( .A(n4409), .B(n4410), .Z(n4408) );
  OR U4551 ( .A(n4411), .B(n4194), .Z(n4235) );
  XOR U4552 ( .A(n4119), .B(n4410), .Z(n4194) );
  XOR U4553 ( .A(n4086), .B(n4232), .Z(n4113) );
  XOR U4554 ( .A(n4237), .B(n4412), .Z(n4232) );
  XOR U4555 ( .A(n4413), .B(n4185), .Z(n4412) );
  OR U4556 ( .A(n4414), .B(n4415), .Z(n4185) );
  ANDN U4557 ( .B(n4416), .A(n4417), .Z(n4413) );
  XOR U4558 ( .A(n4418), .B(n4239), .Z(n4237) );
  OR U4559 ( .A(n4419), .B(n4420), .Z(n4239) );
  ANDN U4560 ( .B(n4421), .A(n4422), .Z(n4418) );
  XNOR U4561 ( .A(n4189), .B(n4423), .Z(n4086) );
  XNOR U4562 ( .A(n4400), .B(n4424), .Z(n4423) );
  NANDN U4563 ( .A(n4425), .B(n4416), .Z(n4424) );
  OR U4564 ( .A(n4414), .B(n4426), .Z(n4400) );
  XOR U4565 ( .A(n4187), .B(n4416), .Z(n4414) );
  XOR U4566 ( .A(n4427), .B(n4404), .Z(n4189) );
  NANDN U4567 ( .A(n4419), .B(n4428), .Z(n4404) );
  XOR U4568 ( .A(n4421), .B(n4241), .Z(n4419) );
  XNOR U4569 ( .A(n4416), .B(n4410), .Z(n4241) );
  IV U4570 ( .A(n4193), .Z(n4410) );
  XNOR U4571 ( .A(n4429), .B(n4430), .Z(n4193) );
  NANDN U4572 ( .A(n4431), .B(n4432), .Z(n4430) );
  XOR U4573 ( .A(n4433), .B(n4434), .Z(n4416) );
  NANDN U4574 ( .A(n4431), .B(n4435), .Z(n4434) );
  XOR U4575 ( .A(n4187), .B(n4119), .Z(n4421) );
  XOR U4576 ( .A(n4437), .B(n4429), .Z(n4119) );
  NANDN U4577 ( .A(n4438), .B(n4439), .Z(n4429) );
  XOR U4578 ( .A(n4432), .B(n4440), .Z(n4439) );
  ANDN U4579 ( .B(n4440), .A(n4441), .Z(n4437) );
  NANDN U4580 ( .A(n4438), .B(n4443), .Z(n4433) );
  XOR U4581 ( .A(n4444), .B(n4445), .Z(n4431) );
  XOR U4582 ( .A(n4446), .B(n4447), .Z(n4445) );
  XNOR U4583 ( .A(n4448), .B(n4449), .Z(n4444) );
  XNOR U4584 ( .A(n4450), .B(n4451), .Z(n4449) );
  ANDN U4585 ( .B(n4447), .A(n4446), .Z(n4450) );
  ANDN U4586 ( .B(n4447), .A(n4441), .Z(n4442) );
  XNOR U4587 ( .A(n4448), .B(n4452), .Z(n4441) );
  XOR U4588 ( .A(n4453), .B(n4451), .Z(n4452) );
  NAND U4589 ( .A(n4443), .B(n4454), .Z(n4451) );
  XNOR U4590 ( .A(n4432), .B(n4446), .Z(n4454) );
  IV U4591 ( .A(n4440), .Z(n4446) );
  XNOR U4592 ( .A(n4455), .B(n4456), .Z(n4440) );
  XNOR U4593 ( .A(n4457), .B(n4458), .Z(n4456) );
  XOR U4594 ( .A(n4425), .B(n4459), .Z(n4458) );
  XNOR U4595 ( .A(n4417), .B(n4460), .Z(n4455) );
  XNOR U4596 ( .A(n4461), .B(n4462), .Z(n4460) );
  AND U4597 ( .A(n4402), .B(n4188), .Z(n4461) );
  XOR U4598 ( .A(n4435), .B(n4447), .Z(n4443) );
  AND U4599 ( .A(n4432), .B(n4435), .Z(n4453) );
  XNOR U4600 ( .A(n4432), .B(n4435), .Z(n4448) );
  XNOR U4601 ( .A(n4463), .B(n4464), .Z(n4435) );
  XNOR U4602 ( .A(n4465), .B(n4459), .Z(n4464) );
  XOR U4603 ( .A(n4466), .B(n4467), .Z(n4463) );
  XNOR U4604 ( .A(n4468), .B(n4469), .Z(n4467) );
  ANDN U4605 ( .B(n4192), .A(n4409), .Z(n4468) );
  XNOR U4606 ( .A(n4470), .B(n4471), .Z(n4432) );
  XNOR U4607 ( .A(n4402), .B(n4466), .Z(n4472) );
  XOR U4608 ( .A(n4188), .B(n4473), .Z(n4470) );
  XNOR U4609 ( .A(n4474), .B(n4462), .Z(n4473) );
  OR U4610 ( .A(n4426), .B(n4415), .Z(n4462) );
  XOR U4611 ( .A(n4188), .B(n4417), .Z(n4415) );
  XNOR U4612 ( .A(n4402), .B(n4475), .Z(n4426) );
  ANDN U4613 ( .B(n4476), .A(n4425), .Z(n4474) );
  XNOR U4614 ( .A(n4477), .B(n4478), .Z(n4447) );
  XOR U4615 ( .A(n4465), .B(n4457), .Z(n4478) );
  XOR U4616 ( .A(n4466), .B(n4479), .Z(n4457) );
  XNOR U4617 ( .A(n4480), .B(n4481), .Z(n4479) );
  NAND U4618 ( .A(n4242), .B(n4406), .Z(n4481) );
  XNOR U4619 ( .A(n4482), .B(n4480), .Z(n4466) );
  NANDN U4620 ( .A(n4420), .B(n4428), .Z(n4480) );
  XOR U4621 ( .A(n4436), .B(n4406), .Z(n4428) );
  XOR U4622 ( .A(n4475), .B(n4192), .Z(n4406) );
  IV U4623 ( .A(n4425), .Z(n4475) );
  XOR U4624 ( .A(n4118), .B(n4483), .Z(n4425) );
  XNOR U4625 ( .A(n4484), .B(n4485), .Z(n4483) );
  XOR U4626 ( .A(n4422), .B(n4242), .Z(n4420) );
  XNOR U4627 ( .A(n4476), .B(n4409), .Z(n4242) );
  IV U4628 ( .A(n4417), .Z(n4476) );
  XOR U4629 ( .A(n4486), .B(n4487), .Z(n4417) );
  XOR U4630 ( .A(n4488), .B(n4489), .Z(n4487) );
  XNOR U4631 ( .A(n4188), .B(n4490), .Z(n4486) );
  ANDN U4632 ( .B(n4436), .A(n4422), .Z(n4482) );
  XNOR U4633 ( .A(n4188), .B(n4491), .Z(n4422) );
  XOR U4634 ( .A(n4491), .B(n4118), .Z(n4465) );
  IV U4635 ( .A(n4236), .Z(n4491) );
  XNOR U4636 ( .A(n4492), .B(n4469), .Z(n4477) );
  OR U4637 ( .A(n4195), .B(n4411), .Z(n4469) );
  XNOR U4638 ( .A(n4236), .B(n4409), .Z(n4411) );
  XOR U4639 ( .A(n4493), .B(n4494), .Z(n4409) );
  XNOR U4640 ( .A(n4118), .B(n4192), .Z(n4195) );
  XOR U4641 ( .A(n4494), .B(n4495), .Z(n4192) );
  XOR U4642 ( .A(n4484), .B(n4493), .Z(n4495) );
  ANDN U4643 ( .B(n4118), .A(n4236), .Z(n4492) );
  XNOR U4644 ( .A(n4485), .B(n4496), .Z(n4236) );
  XOR U4645 ( .A(n4490), .B(n4493), .Z(n4496) );
  IV U4646 ( .A(n4497), .Z(n4493) );
  XNOR U4647 ( .A(n4484), .B(n4498), .Z(n4490) );
  XNOR U4648 ( .A(state[35]), .B(key[35]), .Z(n4498) );
  XNOR U4649 ( .A(state[33]), .B(key[33]), .Z(n4484) );
  XNOR U4650 ( .A(state[34]), .B(key[34]), .Z(n4485) );
  XOR U4651 ( .A(n4402), .B(n4118), .Z(n4436) );
  XOR U4652 ( .A(n4494), .B(n4499), .Z(n4118) );
  XNOR U4653 ( .A(n4497), .B(n4488), .Z(n4499) );
  XNOR U4654 ( .A(state[39]), .B(key[39]), .Z(n4488) );
  XOR U4655 ( .A(n4494), .B(n4500), .Z(n4402) );
  XOR U4656 ( .A(n4497), .B(n4489), .Z(n4500) );
  XOR U4657 ( .A(state[36]), .B(key[36]), .Z(n4489) );
  XOR U4658 ( .A(n4188), .B(n4501), .Z(n4497) );
  XNOR U4659 ( .A(state[38]), .B(key[38]), .Z(n4501) );
  XOR U4660 ( .A(state[32]), .B(key[32]), .Z(n4188) );
  XNOR U4661 ( .A(state[37]), .B(key[37]), .Z(n4494) );
  IV U4662 ( .A(n1827), .Z(n4244) );
  XNOR U4663 ( .A(n4131), .B(n4502), .Z(n1827) );
  XOR U4664 ( .A(n4230), .B(n4231), .Z(n4502) );
  XOR U4665 ( .A(n4223), .B(n4503), .Z(n4231) );
  XNOR U4666 ( .A(n4504), .B(n4505), .Z(n4503) );
  NANDN U4667 ( .A(n4172), .B(n4506), .Z(n4505) );
  XNOR U4668 ( .A(n4174), .B(n4507), .Z(n4223) );
  XNOR U4669 ( .A(n4508), .B(n4509), .Z(n4507) );
  NANDN U4670 ( .A(n4309), .B(n4510), .Z(n4509) );
  IV U4671 ( .A(n4298), .Z(n4230) );
  XOR U4672 ( .A(n4305), .B(n4511), .Z(n4298) );
  XNOR U4673 ( .A(n4303), .B(n4512), .Z(n4511) );
  NANDN U4674 ( .A(n4513), .B(n4514), .Z(n4512) );
  OR U4675 ( .A(n4515), .B(n4226), .Z(n4303) );
  XOR U4676 ( .A(n4229), .B(n4514), .Z(n4226) );
  XOR U4677 ( .A(n4299), .B(n4222), .Z(n4131) );
  XNOR U4678 ( .A(n4174), .B(n4516), .Z(n4222) );
  XNOR U4679 ( .A(n4504), .B(n4517), .Z(n4516) );
  OR U4680 ( .A(n4518), .B(n4519), .Z(n4517) );
  OR U4681 ( .A(n4520), .B(n4521), .Z(n4504) );
  XOR U4682 ( .A(n4522), .B(n4508), .Z(n4174) );
  NANDN U4683 ( .A(n4523), .B(n4524), .Z(n4508) );
  AND U4684 ( .A(n4525), .B(n4526), .Z(n4522) );
  XOR U4685 ( .A(n4305), .B(n4527), .Z(n4299) );
  XOR U4686 ( .A(n4528), .B(n4170), .Z(n4527) );
  OR U4687 ( .A(n4529), .B(n4520), .Z(n4170) );
  XNOR U4688 ( .A(n4172), .B(n4518), .Z(n4520) );
  NOR U4689 ( .A(n4530), .B(n4518), .Z(n4528) );
  XOR U4690 ( .A(n4531), .B(n4307), .Z(n4305) );
  OR U4691 ( .A(n4523), .B(n4532), .Z(n4307) );
  XOR U4692 ( .A(n4518), .B(n4514), .Z(n4309) );
  IV U4693 ( .A(n4179), .Z(n4514) );
  XNOR U4694 ( .A(n4533), .B(n4534), .Z(n4179) );
  NANDN U4695 ( .A(n4535), .B(n4536), .Z(n4534) );
  XNOR U4696 ( .A(n4537), .B(n4538), .Z(n4518) );
  NANDN U4697 ( .A(n4535), .B(n4539), .Z(n4538) );
  ANDN U4698 ( .B(n4525), .A(n4540), .Z(n4531) );
  XOR U4699 ( .A(n4172), .B(n4229), .Z(n4525) );
  XOR U4700 ( .A(n4541), .B(n4533), .Z(n4229) );
  NANDN U4701 ( .A(n4542), .B(n4543), .Z(n4533) );
  XOR U4702 ( .A(n4536), .B(n4544), .Z(n4543) );
  ANDN U4703 ( .B(n4544), .A(n4545), .Z(n4541) );
  NANDN U4704 ( .A(n4542), .B(n4547), .Z(n4537) );
  XOR U4705 ( .A(n4548), .B(n4549), .Z(n4535) );
  XOR U4706 ( .A(n4550), .B(n4551), .Z(n4549) );
  XNOR U4707 ( .A(n4552), .B(n4553), .Z(n4548) );
  XNOR U4708 ( .A(n4554), .B(n4555), .Z(n4553) );
  ANDN U4709 ( .B(n4551), .A(n4550), .Z(n4554) );
  ANDN U4710 ( .B(n4551), .A(n4545), .Z(n4546) );
  XNOR U4711 ( .A(n4552), .B(n4556), .Z(n4545) );
  XOR U4712 ( .A(n4557), .B(n4555), .Z(n4556) );
  NAND U4713 ( .A(n4547), .B(n4558), .Z(n4555) );
  XNOR U4714 ( .A(n4536), .B(n4550), .Z(n4558) );
  IV U4715 ( .A(n4544), .Z(n4550) );
  XNOR U4716 ( .A(n4559), .B(n4560), .Z(n4544) );
  XNOR U4717 ( .A(n4561), .B(n4562), .Z(n4560) );
  XOR U4718 ( .A(n4519), .B(n4563), .Z(n4562) );
  XNOR U4719 ( .A(n4530), .B(n4564), .Z(n4559) );
  XNOR U4720 ( .A(n4565), .B(n4566), .Z(n4564) );
  AND U4721 ( .A(n4506), .B(n4173), .Z(n4565) );
  XOR U4722 ( .A(n4539), .B(n4551), .Z(n4547) );
  AND U4723 ( .A(n4536), .B(n4539), .Z(n4557) );
  XNOR U4724 ( .A(n4536), .B(n4539), .Z(n4552) );
  XNOR U4725 ( .A(n4567), .B(n4568), .Z(n4539) );
  XNOR U4726 ( .A(n4569), .B(n4563), .Z(n4568) );
  XOR U4727 ( .A(n4570), .B(n4571), .Z(n4567) );
  XNOR U4728 ( .A(n4572), .B(n4573), .Z(n4571) );
  ANDN U4729 ( .B(n4178), .A(n4513), .Z(n4572) );
  XNOR U4730 ( .A(n4574), .B(n4575), .Z(n4536) );
  XNOR U4731 ( .A(n4506), .B(n4570), .Z(n4576) );
  XOR U4732 ( .A(n4173), .B(n4577), .Z(n4574) );
  XNOR U4733 ( .A(n4578), .B(n4566), .Z(n4577) );
  OR U4734 ( .A(n4521), .B(n4529), .Z(n4566) );
  XOR U4735 ( .A(n4173), .B(n4530), .Z(n4529) );
  XNOR U4736 ( .A(n4506), .B(n4579), .Z(n4521) );
  ANDN U4737 ( .B(n4580), .A(n4519), .Z(n4578) );
  XNOR U4738 ( .A(n4581), .B(n4582), .Z(n4551) );
  XOR U4739 ( .A(n4569), .B(n4561), .Z(n4582) );
  XOR U4740 ( .A(n4570), .B(n4583), .Z(n4561) );
  XNOR U4741 ( .A(n4584), .B(n4585), .Z(n4583) );
  NAND U4742 ( .A(n4310), .B(n4510), .Z(n4585) );
  XNOR U4743 ( .A(n4586), .B(n4584), .Z(n4570) );
  NANDN U4744 ( .A(n4532), .B(n4524), .Z(n4584) );
  XOR U4745 ( .A(n4526), .B(n4510), .Z(n4524) );
  XOR U4746 ( .A(n4579), .B(n4178), .Z(n4510) );
  IV U4747 ( .A(n4519), .Z(n4579) );
  XOR U4748 ( .A(n4228), .B(n4587), .Z(n4519) );
  XNOR U4749 ( .A(n4588), .B(n4589), .Z(n4587) );
  XOR U4750 ( .A(n4540), .B(n4310), .Z(n4532) );
  XNOR U4751 ( .A(n4580), .B(n4513), .Z(n4310) );
  IV U4752 ( .A(n4530), .Z(n4580) );
  XOR U4753 ( .A(n4590), .B(n4591), .Z(n4530) );
  XOR U4754 ( .A(n4592), .B(n4593), .Z(n4591) );
  XNOR U4755 ( .A(n4173), .B(n4594), .Z(n4590) );
  ANDN U4756 ( .B(n4526), .A(n4540), .Z(n4586) );
  XNOR U4757 ( .A(n4173), .B(n4595), .Z(n4540) );
  XOR U4758 ( .A(n4506), .B(n4228), .Z(n4526) );
  XOR U4759 ( .A(n4596), .B(n4597), .Z(n4506) );
  XOR U4760 ( .A(n4598), .B(n4593), .Z(n4597) );
  XOR U4761 ( .A(state[28]), .B(key[28]), .Z(n4593) );
  XOR U4762 ( .A(n4595), .B(n4228), .Z(n4569) );
  IV U4763 ( .A(n4304), .Z(n4595) );
  XNOR U4764 ( .A(n4599), .B(n4573), .Z(n4581) );
  OR U4765 ( .A(n4227), .B(n4515), .Z(n4573) );
  XNOR U4766 ( .A(n4304), .B(n4513), .Z(n4515) );
  XOR U4767 ( .A(n4600), .B(n4596), .Z(n4513) );
  XNOR U4768 ( .A(n4228), .B(n4178), .Z(n4227) );
  XOR U4769 ( .A(n4596), .B(n4601), .Z(n4178) );
  XOR U4770 ( .A(n4588), .B(n4600), .Z(n4601) );
  ANDN U4771 ( .B(n4228), .A(n4304), .Z(n4599) );
  XNOR U4772 ( .A(n4589), .B(n4602), .Z(n4304) );
  XOR U4773 ( .A(n4594), .B(n4600), .Z(n4602) );
  IV U4774 ( .A(n4598), .Z(n4600) );
  XNOR U4775 ( .A(n4588), .B(n4603), .Z(n4594) );
  XNOR U4776 ( .A(state[27]), .B(key[27]), .Z(n4603) );
  XNOR U4777 ( .A(state[25]), .B(key[25]), .Z(n4588) );
  XNOR U4778 ( .A(state[26]), .B(key[26]), .Z(n4589) );
  XOR U4779 ( .A(n4596), .B(n4604), .Z(n4228) );
  XNOR U4780 ( .A(n4598), .B(n4592), .Z(n4604) );
  XNOR U4781 ( .A(state[31]), .B(key[31]), .Z(n4592) );
  XOR U4782 ( .A(n4173), .B(n4605), .Z(n4598) );
  XNOR U4783 ( .A(state[30]), .B(key[30]), .Z(n4605) );
  XOR U4784 ( .A(state[24]), .B(key[24]), .Z(n4173) );
  XNOR U4785 ( .A(state[29]), .B(key[29]), .Z(n4596) );
  XOR U4786 ( .A(n4163), .B(n4106), .Z(n1216) );
  XNOR U4787 ( .A(n4139), .B(n4606), .Z(n4106) );
  XOR U4788 ( .A(n4607), .B(n4253), .Z(n4606) );
  OR U4789 ( .A(n4608), .B(n4205), .Z(n4253) );
  XOR U4790 ( .A(n4208), .B(n4111), .Z(n4205) );
  NOR U4791 ( .A(n4609), .B(n4208), .Z(n4607) );
  XNOR U4792 ( .A(n4251), .B(n4610), .Z(n4139) );
  XNOR U4793 ( .A(n4611), .B(n4612), .Z(n4610) );
  NANDN U4794 ( .A(n4613), .B(n4265), .Z(n4612) );
  XNOR U4795 ( .A(n4251), .B(n4614), .Z(n4163) );
  XOR U4796 ( .A(n4615), .B(n4141), .Z(n4614) );
  OR U4797 ( .A(n4616), .B(n4259), .Z(n4141) );
  XOR U4798 ( .A(n4143), .B(n4617), .Z(n4259) );
  ANDN U4799 ( .B(n4617), .A(n4618), .Z(n4615) );
  IV U4800 ( .A(n4249), .Z(n4617) );
  XOR U4801 ( .A(n4619), .B(n4611), .Z(n4251) );
  OR U4802 ( .A(n4267), .B(n4620), .Z(n4611) );
  XNOR U4803 ( .A(n4269), .B(n4265), .Z(n4267) );
  XNOR U4804 ( .A(n4111), .B(n4249), .Z(n4265) );
  XNOR U4805 ( .A(n4621), .B(n4622), .Z(n4249) );
  NAND U4806 ( .A(n4623), .B(n4624), .Z(n4622) );
  XOR U4807 ( .A(n4625), .B(n4626), .Z(n4111) );
  NAND U4808 ( .A(n4627), .B(n4623), .Z(n4626) );
  ANDN U4809 ( .B(n4269), .A(n4628), .Z(n4619) );
  XOR U4810 ( .A(n4208), .B(n4143), .Z(n4269) );
  XOR U4811 ( .A(n4629), .B(n4621), .Z(n4143) );
  NANDN U4812 ( .A(n4630), .B(n4631), .Z(n4621) );
  NANDN U4813 ( .A(n4630), .B(n4635), .Z(n4625) );
  XOR U4814 ( .A(n4632), .B(n4623), .Z(n4630) );
  XNOR U4815 ( .A(n4636), .B(n4637), .Z(n4623) );
  XOR U4816 ( .A(n4638), .B(n4633), .Z(n4637) );
  XNOR U4817 ( .A(n4639), .B(n4640), .Z(n4636) );
  XNOR U4818 ( .A(n4641), .B(n4642), .Z(n4640) );
  ANDN U4819 ( .B(n4638), .A(n4633), .Z(n4641) );
  ANDN U4820 ( .B(n4638), .A(n4632), .Z(n4634) );
  XNOR U4821 ( .A(n4639), .B(n4643), .Z(n4632) );
  XOR U4822 ( .A(n4644), .B(n4642), .Z(n4643) );
  NAND U4823 ( .A(n4631), .B(n4635), .Z(n4642) );
  XNOR U4824 ( .A(n4624), .B(n4633), .Z(n4631) );
  XOR U4825 ( .A(n4645), .B(n4646), .Z(n4633) );
  XOR U4826 ( .A(n4647), .B(n4648), .Z(n4646) );
  XNOR U4827 ( .A(n4649), .B(n4650), .Z(n4645) );
  ANDN U4828 ( .B(n4207), .A(n4609), .Z(n4649) );
  AND U4829 ( .A(n4627), .B(n4624), .Z(n4644) );
  XNOR U4830 ( .A(n4627), .B(n4624), .Z(n4639) );
  XNOR U4831 ( .A(n4651), .B(n4652), .Z(n4624) );
  XOR U4832 ( .A(n4653), .B(n4654), .Z(n4652) );
  XOR U4833 ( .A(n4647), .B(n4655), .Z(n4651) );
  XNOR U4834 ( .A(n4656), .B(n4650), .Z(n4655) );
  OR U4835 ( .A(n4206), .B(n4608), .Z(n4650) );
  XOR U4836 ( .A(n4609), .B(n4657), .Z(n4608) );
  XNOR U4837 ( .A(n4207), .B(n4658), .Z(n4206) );
  ANDN U4838 ( .B(n4658), .A(n4255), .Z(n4656) );
  IV U4839 ( .A(n4112), .Z(n4658) );
  XNOR U4840 ( .A(n4659), .B(n4660), .Z(n4627) );
  XNOR U4841 ( .A(n4661), .B(n4662), .Z(n4660) );
  XOR U4842 ( .A(n4258), .B(n4647), .Z(n4662) );
  XNOR U4843 ( .A(n4609), .B(n4207), .Z(n4647) );
  XNOR U4844 ( .A(n4144), .B(n4663), .Z(n4659) );
  XNOR U4845 ( .A(n4664), .B(n4665), .Z(n4663) );
  ANDN U4846 ( .B(n4250), .A(n4618), .Z(n4664) );
  XNOR U4847 ( .A(n4666), .B(n4667), .Z(n4638) );
  XNOR U4848 ( .A(n4648), .B(n4668), .Z(n4667) );
  XOR U4849 ( .A(n4250), .B(n4654), .Z(n4668) );
  XOR U4850 ( .A(n4657), .B(n4112), .Z(n4654) );
  XNOR U4851 ( .A(n4661), .B(n4669), .Z(n4648) );
  XNOR U4852 ( .A(n4670), .B(n4671), .Z(n4669) );
  OR U4853 ( .A(n4613), .B(n4264), .Z(n4671) );
  IV U4854 ( .A(n4653), .Z(n4661) );
  XNOR U4855 ( .A(n4672), .B(n4670), .Z(n4653) );
  NANDN U4856 ( .A(n4620), .B(n4268), .Z(n4670) );
  XOR U4857 ( .A(n4250), .B(n4112), .Z(n4264) );
  XOR U4858 ( .A(n4673), .B(n4674), .Z(n4112) );
  XOR U4859 ( .A(n4675), .B(n4676), .Z(n4674) );
  XOR U4860 ( .A(n4657), .B(n4618), .Z(n4613) );
  IV U4861 ( .A(n4255), .Z(n4657) );
  ANDN U4862 ( .B(n4270), .A(n4628), .Z(n4672) );
  XOR U4863 ( .A(n4677), .B(n4609), .Z(n4628) );
  XOR U4864 ( .A(n4678), .B(n4679), .Z(n4609) );
  XOR U4865 ( .A(n4680), .B(n4675), .Z(n4679) );
  XOR U4866 ( .A(n4681), .B(n4207), .Z(n4270) );
  XNOR U4867 ( .A(n4618), .B(n4682), .Z(n4666) );
  XNOR U4868 ( .A(n4683), .B(n4665), .Z(n4682) );
  OR U4869 ( .A(n4260), .B(n4616), .Z(n4665) );
  XNOR U4870 ( .A(n4144), .B(n4618), .Z(n4616) );
  XOR U4871 ( .A(n4258), .B(n4250), .Z(n4260) );
  XNOR U4872 ( .A(n4207), .B(n4684), .Z(n4250) );
  XNOR U4873 ( .A(n4680), .B(n4676), .Z(n4684) );
  XNOR U4874 ( .A(state[74]), .B(key[74]), .Z(n4680) );
  XOR U4875 ( .A(n4685), .B(n4686), .Z(n4207) );
  IV U4876 ( .A(n4681), .Z(n4258) );
  ANDN U4877 ( .B(n4681), .A(n4144), .Z(n4683) );
  XOR U4878 ( .A(n4687), .B(n4686), .Z(n4681) );
  XNOR U4879 ( .A(n4675), .B(n4673), .Z(n4686) );
  XOR U4880 ( .A(state[77]), .B(key[77]), .Z(n4673) );
  XNOR U4881 ( .A(n4677), .B(n4688), .Z(n4675) );
  XNOR U4882 ( .A(state[78]), .B(key[78]), .Z(n4688) );
  XOR U4883 ( .A(n4689), .B(n4690), .Z(n4618) );
  XNOR U4884 ( .A(n4687), .B(n4685), .Z(n4690) );
  XNOR U4885 ( .A(state[79]), .B(key[79]), .Z(n4685) );
  XNOR U4886 ( .A(state[76]), .B(key[76]), .Z(n4687) );
  XNOR U4887 ( .A(n4144), .B(n4678), .Z(n4689) );
  XOR U4888 ( .A(n4676), .B(n4691), .Z(n4678) );
  XNOR U4889 ( .A(state[75]), .B(key[75]), .Z(n4691) );
  XNOR U4890 ( .A(state[73]), .B(key[73]), .Z(n4676) );
  IV U4891 ( .A(n4677), .Z(n4144) );
  XOR U4892 ( .A(state[72]), .B(key[72]), .Z(n4677) );
  XNOR U4893 ( .A(n854), .B(n4692), .Z(out[0]) );
  XOR U4894 ( .A(key[128]), .B(n1651), .Z(n4692) );
  XNOR U4895 ( .A(n1876), .B(n4693), .Z(n1651) );
  XOR U4896 ( .A(n4694), .B(n858), .Z(n4693) );
  OR U4897 ( .A(n4695), .B(n1869), .Z(n858) );
  XNOR U4898 ( .A(n861), .B(n1868), .Z(n1869) );
  ANDN U4899 ( .B(n4696), .A(n4697), .Z(n4694) );
  IV U4900 ( .A(n1084), .Z(n854) );
  XOR U4901 ( .A(n862), .B(n4698), .Z(n1084) );
  XOR U4902 ( .A(n4699), .B(n1878), .Z(n4698) );
  XNOR U4903 ( .A(n1445), .B(n866), .Z(n1442) );
  NOR U4904 ( .A(n4701), .B(n1445), .Z(n4699) );
  XNOR U4905 ( .A(n1876), .B(n4702), .Z(n862) );
  XNOR U4906 ( .A(n4703), .B(n4704), .Z(n4702) );
  NANDN U4907 ( .A(n1863), .B(n4705), .Z(n4704) );
  XOR U4908 ( .A(n4706), .B(n4703), .Z(n1876) );
  OR U4909 ( .A(n1872), .B(n4707), .Z(n4703) );
  XOR U4910 ( .A(n4708), .B(n1863), .Z(n1872) );
  XNOR U4911 ( .A(n1868), .B(n866), .Z(n1863) );
  XOR U4912 ( .A(n4709), .B(n4710), .Z(n866) );
  NANDN U4913 ( .A(n4711), .B(n4712), .Z(n4710) );
  IV U4914 ( .A(n4697), .Z(n1868) );
  XNOR U4915 ( .A(n4713), .B(n4714), .Z(n4697) );
  NANDN U4916 ( .A(n4711), .B(n4715), .Z(n4714) );
  ANDN U4917 ( .B(n4708), .A(n4716), .Z(n4706) );
  IV U4918 ( .A(n1875), .Z(n4708) );
  XOR U4919 ( .A(n1445), .B(n861), .Z(n1875) );
  XNOR U4920 ( .A(n4717), .B(n4713), .Z(n861) );
  NANDN U4921 ( .A(n4718), .B(n4719), .Z(n4713) );
  XOR U4922 ( .A(n4715), .B(n4720), .Z(n4719) );
  ANDN U4923 ( .B(n4720), .A(n4721), .Z(n4717) );
  XOR U4924 ( .A(n4722), .B(n4709), .Z(n1445) );
  NANDN U4925 ( .A(n4718), .B(n4723), .Z(n4709) );
  XOR U4926 ( .A(n4724), .B(n4712), .Z(n4723) );
  XNOR U4927 ( .A(n4725), .B(n4726), .Z(n4711) );
  XOR U4928 ( .A(n4727), .B(n4728), .Z(n4726) );
  XNOR U4929 ( .A(n4729), .B(n4730), .Z(n4725) );
  XNOR U4930 ( .A(n4731), .B(n4732), .Z(n4730) );
  ANDN U4931 ( .B(n4724), .A(n4728), .Z(n4731) );
  ANDN U4932 ( .B(n4724), .A(n4721), .Z(n4722) );
  XNOR U4933 ( .A(n4727), .B(n4733), .Z(n4721) );
  XOR U4934 ( .A(n4734), .B(n4732), .Z(n4733) );
  NAND U4935 ( .A(n4735), .B(n4736), .Z(n4732) );
  XNOR U4936 ( .A(n4729), .B(n4712), .Z(n4736) );
  IV U4937 ( .A(n4724), .Z(n4729) );
  XNOR U4938 ( .A(n4715), .B(n4728), .Z(n4735) );
  IV U4939 ( .A(n4720), .Z(n4728) );
  XOR U4940 ( .A(n4737), .B(n4738), .Z(n4720) );
  XNOR U4941 ( .A(n4739), .B(n4740), .Z(n4738) );
  XNOR U4942 ( .A(n4741), .B(n4742), .Z(n4737) );
  ANDN U4943 ( .B(n4743), .A(n4701), .Z(n4741) );
  AND U4944 ( .A(n4712), .B(n4715), .Z(n4734) );
  XNOR U4945 ( .A(n4712), .B(n4715), .Z(n4727) );
  XNOR U4946 ( .A(n4744), .B(n4745), .Z(n4715) );
  XNOR U4947 ( .A(n4746), .B(n4740), .Z(n4745) );
  XOR U4948 ( .A(n4747), .B(n4748), .Z(n4744) );
  XNOR U4949 ( .A(n4749), .B(n4742), .Z(n4748) );
  OR U4950 ( .A(n1443), .B(n4700), .Z(n4742) );
  XNOR U4951 ( .A(n4750), .B(n1880), .Z(n4700) );
  XNOR U4952 ( .A(n1444), .B(n867), .Z(n1443) );
  ANDN U4953 ( .B(n1880), .A(n867), .Z(n4749) );
  XNOR U4954 ( .A(n4751), .B(n4752), .Z(n4712) );
  XNOR U4955 ( .A(n4740), .B(n4753), .Z(n4752) );
  XOR U4956 ( .A(n1859), .B(n4747), .Z(n4753) );
  XNOR U4957 ( .A(n4750), .B(n1444), .Z(n4740) );
  XNOR U4958 ( .A(n4754), .B(n4755), .Z(n4751) );
  XNOR U4959 ( .A(n4756), .B(n4757), .Z(n4755) );
  ANDN U4960 ( .B(n4696), .A(n1867), .Z(n4756) );
  XNOR U4961 ( .A(n4758), .B(n4759), .Z(n4724) );
  XNOR U4962 ( .A(n4746), .B(n4760), .Z(n4759) );
  XNOR U4963 ( .A(n1867), .B(n4739), .Z(n4760) );
  XOR U4964 ( .A(n4747), .B(n4761), .Z(n4739) );
  XNOR U4965 ( .A(n4762), .B(n4763), .Z(n4761) );
  NAND U4966 ( .A(n4705), .B(n1864), .Z(n4763) );
  XNOR U4967 ( .A(n4764), .B(n4762), .Z(n4747) );
  NANDN U4968 ( .A(n4707), .B(n1873), .Z(n4762) );
  XOR U4969 ( .A(n1874), .B(n1864), .Z(n1873) );
  XNOR U4970 ( .A(n4765), .B(n867), .Z(n1864) );
  XOR U4971 ( .A(n4716), .B(n4705), .Z(n4707) );
  XOR U4972 ( .A(n4696), .B(n1880), .Z(n4705) );
  ANDN U4973 ( .B(n1874), .A(n4716), .Z(n4764) );
  XNOR U4974 ( .A(n4754), .B(n4750), .Z(n4716) );
  IV U4975 ( .A(n4701), .Z(n4750) );
  XNOR U4976 ( .A(n4766), .B(n4767), .Z(n4701) );
  XOR U4977 ( .A(n4768), .B(n4769), .Z(n4767) );
  XOR U4978 ( .A(n4770), .B(n4743), .Z(n1874) );
  XNOR U4979 ( .A(n4771), .B(n4772), .Z(n867) );
  XNOR U4980 ( .A(n4773), .B(n4769), .Z(n4772) );
  XNOR U4981 ( .A(n4769), .B(n4771), .Z(n1880) );
  XNOR U4982 ( .A(n4696), .B(n4774), .Z(n4758) );
  XNOR U4983 ( .A(n4775), .B(n4757), .Z(n4774) );
  OR U4984 ( .A(n1870), .B(n4695), .Z(n4757) );
  XNOR U4985 ( .A(n4754), .B(n4696), .Z(n4695) );
  XOR U4986 ( .A(n1859), .B(n4765), .Z(n1870) );
  IV U4987 ( .A(n1867), .Z(n4765) );
  XOR U4988 ( .A(n4743), .B(n4776), .Z(n1867) );
  XOR U4989 ( .A(n4773), .B(n4766), .Z(n4776) );
  XNOR U4990 ( .A(key[162]), .B(\w0[1][34] ), .Z(n4766) );
  XOR U4991 ( .A(n3939), .B(n4777), .Z(\w0[1][34] ) );
  XNOR U4992 ( .A(n1035), .B(n995), .Z(n4777) );
  XOR U4993 ( .A(n1036), .B(n379), .Z(n995) );
  XOR U4994 ( .A(n1029), .B(n994), .Z(n3939) );
  XNOR U4995 ( .A(n4778), .B(n4779), .Z(n1029) );
  XNOR U4996 ( .A(n4780), .B(n4781), .Z(n4779) );
  XNOR U4997 ( .A(n4782), .B(n4783), .Z(n4778) );
  IV U4998 ( .A(n1444), .Z(n4743) );
  XNOR U4999 ( .A(n4771), .B(n4784), .Z(n1444) );
  XNOR U5000 ( .A(n4769), .B(n4785), .Z(n4784) );
  ANDN U5001 ( .B(n4770), .A(n860), .Z(n4775) );
  IV U5002 ( .A(n1859), .Z(n4770) );
  XNOR U5003 ( .A(n4771), .B(n4786), .Z(n1859) );
  XNOR U5004 ( .A(n4769), .B(n4787), .Z(n4786) );
  XOR U5005 ( .A(n860), .B(n4788), .Z(n4769) );
  XOR U5006 ( .A(key[166]), .B(\w0[1][38] ), .Z(n4788) );
  XNOR U5007 ( .A(n3915), .B(n4789), .Z(\w0[1][38] ) );
  XOR U5008 ( .A(n1004), .B(n1010), .Z(n4789) );
  XNOR U5009 ( .A(n392), .B(n4790), .Z(n1004) );
  XOR U5010 ( .A(n1011), .B(n3923), .Z(n392) );
  IV U5011 ( .A(n388), .Z(n3923) );
  XOR U5012 ( .A(n4791), .B(n4792), .Z(n388) );
  XOR U5013 ( .A(n4793), .B(n4794), .Z(n1011) );
  XNOR U5014 ( .A(n1017), .B(n4795), .Z(n3915) );
  XOR U5015 ( .A(n4796), .B(n4797), .Z(n1017) );
  XNOR U5016 ( .A(n4798), .B(n4780), .Z(n4797) );
  IV U5017 ( .A(n4754), .Z(n860) );
  XOR U5018 ( .A(key[165]), .B(\w0[1][37] ), .Z(n4771) );
  XOR U5019 ( .A(n3917), .B(n4800), .Z(\w0[1][37] ) );
  XOR U5020 ( .A(n1012), .B(n3922), .Z(n4800) );
  XNOR U5021 ( .A(n1024), .B(n393), .Z(n1012) );
  XNOR U5022 ( .A(n4801), .B(n4802), .Z(n393) );
  XNOR U5023 ( .A(n4803), .B(n4804), .Z(n4802) );
  XOR U5024 ( .A(n4805), .B(n4806), .Z(n4801) );
  XOR U5025 ( .A(n4807), .B(n4808), .Z(n4806) );
  ANDN U5026 ( .B(n4809), .A(n4810), .Z(n4808) );
  XNOR U5027 ( .A(n4811), .B(n4812), .Z(n1024) );
  XOR U5028 ( .A(n4813), .B(n4814), .Z(n4812) );
  XNOR U5029 ( .A(n4815), .B(n4816), .Z(n4811) );
  XNOR U5030 ( .A(n4817), .B(n4818), .Z(n4816) );
  ANDN U5031 ( .B(n4819), .A(n4820), .Z(n4818) );
  XOR U5032 ( .A(n3924), .B(n1010), .Z(n3917) );
  XOR U5033 ( .A(n4821), .B(n4822), .Z(n1010) );
  XOR U5034 ( .A(n4798), .B(n4781), .Z(n3924) );
  XOR U5035 ( .A(n4823), .B(n4824), .Z(n4781) );
  XNOR U5036 ( .A(n4825), .B(n4826), .Z(n4824) );
  NOR U5037 ( .A(n4827), .B(n4828), .Z(n4825) );
  XOR U5038 ( .A(n4829), .B(n4830), .Z(n4696) );
  XNOR U5039 ( .A(n4787), .B(n4785), .Z(n4830) );
  XOR U5040 ( .A(key[167]), .B(\w0[1][39] ), .Z(n4785) );
  XNOR U5041 ( .A(n4795), .B(n4831), .Z(\w0[1][39] ) );
  XNOR U5042 ( .A(n1018), .B(n4790), .Z(n4831) );
  XNOR U5043 ( .A(n419), .B(n3930), .Z(n4790) );
  XNOR U5044 ( .A(n4832), .B(n4833), .Z(n3930) );
  XNOR U5045 ( .A(n4835), .B(n4836), .Z(n4832) );
  IV U5046 ( .A(n4837), .Z(n419) );
  XNOR U5047 ( .A(n1006), .B(n3918), .Z(n1018) );
  XOR U5048 ( .A(n4838), .B(n4839), .Z(n3918) );
  XOR U5049 ( .A(n4840), .B(n4791), .Z(n4839) );
  XNOR U5050 ( .A(n4843), .B(n4844), .Z(n4842) );
  OR U5051 ( .A(n4845), .B(n4846), .Z(n4844) );
  XOR U5052 ( .A(n4848), .B(n4849), .Z(n1006) );
  XOR U5053 ( .A(n4850), .B(n4793), .Z(n4849) );
  XNOR U5054 ( .A(n4852), .B(n4853), .Z(n4815) );
  XNOR U5055 ( .A(n4854), .B(n4855), .Z(n4853) );
  OR U5056 ( .A(n4856), .B(n4857), .Z(n4855) );
  XOR U5057 ( .A(key[164]), .B(\w0[1][36] ), .Z(n4787) );
  XOR U5058 ( .A(n4858), .B(n4859), .Z(\w0[1][36] ) );
  XNOR U5059 ( .A(n3934), .B(n3933), .Z(n4859) );
  XNOR U5060 ( .A(n1009), .B(n3928), .Z(n3933) );
  XOR U5061 ( .A(n4860), .B(n4861), .Z(n1009) );
  XNOR U5062 ( .A(n4862), .B(n4863), .Z(n4861) );
  XOR U5063 ( .A(n4799), .B(n4864), .Z(n4860) );
  XOR U5064 ( .A(n4826), .B(n4865), .Z(n4864) );
  ANDN U5065 ( .B(n4866), .A(n4867), .Z(n4865) );
  NOR U5066 ( .A(n4868), .B(n4869), .Z(n4826) );
  XNOR U5067 ( .A(n4871), .B(n4872), .Z(n4870) );
  OR U5068 ( .A(n4873), .B(n4874), .Z(n4872) );
  XOR U5069 ( .A(n1023), .B(n1022), .Z(n4858) );
  XOR U5070 ( .A(n4804), .B(n379), .Z(n405) );
  XOR U5071 ( .A(n4841), .B(n4876), .Z(n379) );
  XNOR U5072 ( .A(n4814), .B(n1036), .Z(n1031) );
  XNOR U5073 ( .A(n4851), .B(n4877), .Z(n1036) );
  XOR U5074 ( .A(n4837), .B(n3922), .Z(n1023) );
  XNOR U5075 ( .A(n4878), .B(n4879), .Z(n3922) );
  XNOR U5076 ( .A(n4835), .B(n4880), .Z(n4879) );
  XNOR U5077 ( .A(n4881), .B(n4882), .Z(n4835) );
  XNOR U5078 ( .A(n4883), .B(n4884), .Z(n4882) );
  OR U5079 ( .A(n4885), .B(n4886), .Z(n4884) );
  XNOR U5080 ( .A(n4887), .B(n4888), .Z(n4878) );
  XNOR U5081 ( .A(n4889), .B(n4890), .Z(n4888) );
  ANDN U5082 ( .B(n4891), .A(n4892), .Z(n4890) );
  XNOR U5083 ( .A(n4754), .B(n4768), .Z(n4829) );
  XOR U5084 ( .A(n4773), .B(n4893), .Z(n4768) );
  XOR U5085 ( .A(key[163]), .B(\w0[1][35] ), .Z(n4893) );
  XOR U5086 ( .A(n4894), .B(n4895), .Z(\w0[1][35] ) );
  XNOR U5087 ( .A(n994), .B(n3938), .Z(n4895) );
  XNOR U5088 ( .A(n1021), .B(n3928), .Z(n3938) );
  IV U5089 ( .A(n4795), .Z(n3928) );
  XOR U5090 ( .A(n4896), .B(n4863), .Z(n4795) );
  XOR U5091 ( .A(n4863), .B(n3942), .Z(n1021) );
  IV U5092 ( .A(n996), .Z(n3942) );
  XNOR U5093 ( .A(n4875), .B(n4897), .Z(n4863) );
  XOR U5094 ( .A(n4898), .B(n4899), .Z(n4897) );
  NOR U5095 ( .A(n4900), .B(n4828), .Z(n4898) );
  XNOR U5096 ( .A(n4901), .B(n4902), .Z(n4875) );
  XNOR U5097 ( .A(n4903), .B(n4904), .Z(n4902) );
  NANDN U5098 ( .A(n4905), .B(n4906), .Z(n4904) );
  XNOR U5099 ( .A(n4907), .B(n4908), .Z(n994) );
  XNOR U5100 ( .A(n4834), .B(n4822), .Z(n4908) );
  XOR U5101 ( .A(n4909), .B(n4910), .Z(n4822) );
  XOR U5102 ( .A(n4911), .B(n4889), .Z(n4910) );
  NANDN U5103 ( .A(n4912), .B(n4913), .Z(n4889) );
  NOR U5104 ( .A(n4914), .B(n4915), .Z(n4911) );
  XNOR U5105 ( .A(n4836), .B(n4916), .Z(n4907) );
  XOR U5106 ( .A(n1030), .B(n1028), .Z(n4894) );
  IV U5107 ( .A(n380), .Z(n1028) );
  XOR U5108 ( .A(n997), .B(n412), .Z(n380) );
  XOR U5109 ( .A(n4917), .B(n4918), .Z(n412) );
  XOR U5110 ( .A(n4919), .B(n4792), .Z(n4918) );
  XNOR U5111 ( .A(n4920), .B(n4921), .Z(n4792) );
  XNOR U5112 ( .A(n4922), .B(n4807), .Z(n4921) );
  NOR U5113 ( .A(n4923), .B(n4924), .Z(n4807) );
  NOR U5114 ( .A(n4925), .B(n4926), .Z(n4922) );
  XOR U5115 ( .A(n4841), .B(n4840), .Z(n4917) );
  XOR U5116 ( .A(n4927), .B(n4928), .Z(n997) );
  XOR U5117 ( .A(n4929), .B(n4794), .Z(n4928) );
  XNOR U5118 ( .A(n4930), .B(n4931), .Z(n4794) );
  XOR U5119 ( .A(n4932), .B(n4817), .Z(n4931) );
  NANDN U5120 ( .A(n4933), .B(n4934), .Z(n4817) );
  NOR U5121 ( .A(n4935), .B(n4936), .Z(n4932) );
  XOR U5122 ( .A(n4851), .B(n4850), .Z(n4927) );
  XOR U5123 ( .A(n4837), .B(n3934), .Z(n1030) );
  XNOR U5124 ( .A(n4887), .B(n1035), .Z(n3934) );
  XOR U5125 ( .A(key[161]), .B(\w0[1][33] ), .Z(n4773) );
  XNOR U5126 ( .A(n377), .B(n4937), .Z(\w0[1][33] ) );
  XOR U5127 ( .A(n420), .B(n1039), .Z(n4937) );
  XNOR U5128 ( .A(n1040), .B(n416), .Z(n420) );
  XOR U5129 ( .A(n4791), .B(n4938), .Z(n416) );
  XNOR U5130 ( .A(n4841), .B(n4840), .Z(n4938) );
  XNOR U5131 ( .A(n4920), .B(n4939), .Z(n4840) );
  XNOR U5132 ( .A(n4940), .B(n4941), .Z(n4939) );
  OR U5133 ( .A(n4845), .B(n4942), .Z(n4941) );
  XOR U5134 ( .A(n4803), .B(n4943), .Z(n4920) );
  XNOR U5135 ( .A(n4944), .B(n4945), .Z(n4943) );
  OR U5136 ( .A(n4946), .B(n4947), .Z(n4945) );
  XOR U5137 ( .A(n4948), .B(n4949), .Z(n4841) );
  XNOR U5138 ( .A(n4950), .B(n4951), .Z(n4949) );
  OR U5139 ( .A(n4952), .B(n4810), .Z(n4951) );
  XOR U5140 ( .A(n4876), .B(n4919), .Z(n4791) );
  XNOR U5141 ( .A(n4803), .B(n4953), .Z(n4919) );
  XNOR U5142 ( .A(n4940), .B(n4954), .Z(n4953) );
  NANDN U5143 ( .A(n4955), .B(n4956), .Z(n4954) );
  OR U5144 ( .A(n4957), .B(n4958), .Z(n4940) );
  XOR U5145 ( .A(n4959), .B(n4944), .Z(n4803) );
  NANDN U5146 ( .A(n4960), .B(n4961), .Z(n4944) );
  AND U5147 ( .A(n4962), .B(n4963), .Z(n4959) );
  XNOR U5148 ( .A(n4793), .B(n4964), .Z(n1040) );
  XNOR U5149 ( .A(n4851), .B(n4850), .Z(n4964) );
  XNOR U5150 ( .A(n4930), .B(n4965), .Z(n4850) );
  XNOR U5151 ( .A(n4966), .B(n4967), .Z(n4965) );
  OR U5152 ( .A(n4856), .B(n4968), .Z(n4967) );
  XOR U5153 ( .A(n4813), .B(n4969), .Z(n4930) );
  XNOR U5154 ( .A(n4970), .B(n4971), .Z(n4969) );
  OR U5155 ( .A(n4972), .B(n4973), .Z(n4971) );
  XOR U5156 ( .A(n4974), .B(n4975), .Z(n4851) );
  XOR U5157 ( .A(n4976), .B(n4977), .Z(n4975) );
  OR U5158 ( .A(n4978), .B(n4820), .Z(n4977) );
  XOR U5159 ( .A(n4979), .B(n4929), .Z(n4793) );
  XNOR U5160 ( .A(n4813), .B(n4980), .Z(n4929) );
  XNOR U5161 ( .A(n4966), .B(n4981), .Z(n4980) );
  NANDN U5162 ( .A(n4982), .B(n4983), .Z(n4981) );
  OR U5163 ( .A(n4984), .B(n4985), .Z(n4966) );
  XOR U5164 ( .A(n4986), .B(n4970), .Z(n4813) );
  NANDN U5165 ( .A(n4987), .B(n4988), .Z(n4970) );
  AND U5166 ( .A(n4989), .B(n4990), .Z(n4986) );
  XOR U5167 ( .A(n996), .B(n1035), .Z(n377) );
  XNOR U5168 ( .A(n4991), .B(n4836), .Z(n1035) );
  XNOR U5169 ( .A(n4782), .B(n4896), .Z(n996) );
  XOR U5170 ( .A(key[160]), .B(\w0[1][32] ), .Z(n4754) );
  XNOR U5171 ( .A(n413), .B(n4992), .Z(\w0[1][32] ) );
  XNOR U5172 ( .A(n1015), .B(n3919), .Z(n4992) );
  XOR U5173 ( .A(n4876), .B(n4804), .Z(n3919) );
  XNOR U5174 ( .A(n4847), .B(n4993), .Z(n4804) );
  XOR U5175 ( .A(n4994), .B(n4950), .Z(n4993) );
  OR U5176 ( .A(n4995), .B(n4923), .Z(n4950) );
  XNOR U5177 ( .A(n4926), .B(n4810), .Z(n4923) );
  NOR U5178 ( .A(n4996), .B(n4926), .Z(n4994) );
  XNOR U5179 ( .A(n4948), .B(n4997), .Z(n4847) );
  XNOR U5180 ( .A(n4998), .B(n4999), .Z(n4997) );
  NANDN U5181 ( .A(n4946), .B(n5000), .Z(n4999) );
  XOR U5182 ( .A(n4948), .B(n5001), .Z(n4876) );
  XOR U5183 ( .A(n5002), .B(n4843), .Z(n5001) );
  OR U5184 ( .A(n5003), .B(n4957), .Z(n4843) );
  XOR U5185 ( .A(n4845), .B(n5004), .Z(n4957) );
  ANDN U5186 ( .B(n5005), .A(n4955), .Z(n5002) );
  XOR U5187 ( .A(n5006), .B(n4998), .Z(n4948) );
  OR U5188 ( .A(n4960), .B(n5007), .Z(n4998) );
  XOR U5189 ( .A(n4962), .B(n4946), .Z(n4960) );
  XOR U5190 ( .A(n5004), .B(n4810), .Z(n4946) );
  XNOR U5191 ( .A(n5008), .B(n5009), .Z(n4810) );
  NANDN U5192 ( .A(n5010), .B(n5011), .Z(n5009) );
  IV U5193 ( .A(n4955), .Z(n5004) );
  XNOR U5194 ( .A(n5012), .B(n5013), .Z(n4955) );
  NANDN U5195 ( .A(n5010), .B(n5014), .Z(n5013) );
  ANDN U5196 ( .B(n4962), .A(n5015), .Z(n5006) );
  XOR U5197 ( .A(n4926), .B(n4845), .Z(n4962) );
  XOR U5198 ( .A(n5016), .B(n5012), .Z(n4845) );
  NANDN U5199 ( .A(n5017), .B(n5018), .Z(n5012) );
  NANDN U5200 ( .A(n5017), .B(n5022), .Z(n5008) );
  XOR U5201 ( .A(n5023), .B(n5024), .Z(n5010) );
  XOR U5202 ( .A(n5025), .B(n5020), .Z(n5024) );
  XNOR U5203 ( .A(n5026), .B(n5027), .Z(n5023) );
  XNOR U5204 ( .A(n5028), .B(n5029), .Z(n5027) );
  ANDN U5205 ( .B(n5025), .A(n5020), .Z(n5028) );
  ANDN U5206 ( .B(n5025), .A(n5019), .Z(n5021) );
  XNOR U5207 ( .A(n5026), .B(n5030), .Z(n5019) );
  XOR U5208 ( .A(n5031), .B(n5029), .Z(n5030) );
  NAND U5209 ( .A(n5018), .B(n5022), .Z(n5029) );
  XNOR U5210 ( .A(n5014), .B(n5020), .Z(n5018) );
  XOR U5211 ( .A(n5032), .B(n5033), .Z(n5020) );
  XOR U5212 ( .A(n5034), .B(n5035), .Z(n5033) );
  XNOR U5213 ( .A(n5036), .B(n5037), .Z(n5032) );
  ANDN U5214 ( .B(n5038), .A(n4925), .Z(n5036) );
  AND U5215 ( .A(n5011), .B(n5014), .Z(n5031) );
  XNOR U5216 ( .A(n5011), .B(n5014), .Z(n5026) );
  XNOR U5217 ( .A(n5039), .B(n5040), .Z(n5014) );
  XNOR U5218 ( .A(n5041), .B(n5042), .Z(n5040) );
  XOR U5219 ( .A(n5034), .B(n5043), .Z(n5039) );
  XNOR U5220 ( .A(n5044), .B(n5037), .Z(n5043) );
  OR U5221 ( .A(n4924), .B(n4995), .Z(n5037) );
  XNOR U5222 ( .A(n4996), .B(n4952), .Z(n4995) );
  XNOR U5223 ( .A(n4925), .B(n5045), .Z(n4924) );
  NOR U5224 ( .A(n5045), .B(n4952), .Z(n5044) );
  XNOR U5225 ( .A(n5046), .B(n5047), .Z(n5011) );
  XNOR U5226 ( .A(n5048), .B(n5049), .Z(n5047) );
  XOR U5227 ( .A(n4942), .B(n5034), .Z(n5049) );
  XOR U5228 ( .A(n5038), .B(n5050), .Z(n5034) );
  XNOR U5229 ( .A(n4846), .B(n5051), .Z(n5046) );
  XNOR U5230 ( .A(n5052), .B(n5053), .Z(n5051) );
  ANDN U5231 ( .B(n4956), .A(n5054), .Z(n5052) );
  XNOR U5232 ( .A(n5055), .B(n5056), .Z(n5025) );
  XNOR U5233 ( .A(n5035), .B(n5057), .Z(n5056) );
  XNOR U5234 ( .A(n4956), .B(n5042), .Z(n5057) );
  XOR U5235 ( .A(n4952), .B(n5045), .Z(n5042) );
  XNOR U5236 ( .A(n5048), .B(n5058), .Z(n5035) );
  XNOR U5237 ( .A(n5059), .B(n5060), .Z(n5058) );
  NANDN U5238 ( .A(n4947), .B(n5000), .Z(n5060) );
  IV U5239 ( .A(n5041), .Z(n5048) );
  XNOR U5240 ( .A(n5061), .B(n5059), .Z(n5041) );
  NANDN U5241 ( .A(n5007), .B(n4961), .Z(n5059) );
  XOR U5242 ( .A(n4956), .B(n5045), .Z(n4947) );
  IV U5243 ( .A(n4809), .Z(n5045) );
  XOR U5244 ( .A(n5062), .B(n5063), .Z(n4809) );
  XNOR U5245 ( .A(n5064), .B(n5065), .Z(n5063) );
  XOR U5246 ( .A(n5015), .B(n5000), .Z(n5007) );
  XNOR U5247 ( .A(n5005), .B(n4952), .Z(n5000) );
  XNOR U5248 ( .A(n5065), .B(n5062), .Z(n4952) );
  ANDN U5249 ( .B(n4963), .A(n5015), .Z(n5061) );
  XNOR U5250 ( .A(n5066), .B(n5038), .Z(n5015) );
  IV U5251 ( .A(n4996), .Z(n5038) );
  XNOR U5252 ( .A(n5067), .B(n5068), .Z(n4996) );
  XNOR U5253 ( .A(n5069), .B(n5065), .Z(n5068) );
  XOR U5254 ( .A(n5070), .B(n5050), .Z(n4963) );
  XNOR U5255 ( .A(n5054), .B(n5071), .Z(n5055) );
  XNOR U5256 ( .A(n5072), .B(n5053), .Z(n5071) );
  OR U5257 ( .A(n4958), .B(n5003), .Z(n5053) );
  XOR U5258 ( .A(n4846), .B(n5005), .Z(n5003) );
  IV U5259 ( .A(n5054), .Z(n5005) );
  XOR U5260 ( .A(n4942), .B(n4956), .Z(n4958) );
  XNOR U5261 ( .A(n5050), .B(n5073), .Z(n4956) );
  XNOR U5262 ( .A(n5064), .B(n5067), .Z(n5073) );
  XNOR U5263 ( .A(state[106]), .B(key[106]), .Z(n5067) );
  IV U5264 ( .A(n4925), .Z(n5050) );
  XOR U5265 ( .A(n5074), .B(n5075), .Z(n4925) );
  XOR U5266 ( .A(n5065), .B(n5076), .Z(n5075) );
  IV U5267 ( .A(n5070), .Z(n4942) );
  ANDN U5268 ( .B(n5070), .A(n4846), .Z(n5072) );
  XOR U5269 ( .A(n5062), .B(n5077), .Z(n5070) );
  XNOR U5270 ( .A(n5065), .B(n5078), .Z(n5077) );
  XOR U5271 ( .A(n5066), .B(n5079), .Z(n5065) );
  XNOR U5272 ( .A(state[110]), .B(key[110]), .Z(n5079) );
  IV U5273 ( .A(n5074), .Z(n5062) );
  XOR U5274 ( .A(state[109]), .B(key[109]), .Z(n5074) );
  XOR U5275 ( .A(n5080), .B(n5081), .Z(n5054) );
  XOR U5276 ( .A(n5078), .B(n5076), .Z(n5081) );
  XOR U5277 ( .A(state[111]), .B(key[111]), .Z(n5076) );
  XNOR U5278 ( .A(state[108]), .B(key[108]), .Z(n5078) );
  XOR U5279 ( .A(n4846), .B(n5069), .Z(n5080) );
  XNOR U5280 ( .A(n5064), .B(n5082), .Z(n5069) );
  XNOR U5281 ( .A(state[107]), .B(key[107]), .Z(n5082) );
  XNOR U5282 ( .A(state[105]), .B(key[105]), .Z(n5064) );
  IV U5283 ( .A(n5066), .Z(n4846) );
  XOR U5284 ( .A(state[104]), .B(key[104]), .Z(n5066) );
  XOR U5285 ( .A(n4837), .B(n398), .Z(n1015) );
  XOR U5286 ( .A(n4979), .B(n4814), .Z(n398) );
  XOR U5287 ( .A(n4852), .B(n5083), .Z(n4814) );
  XNOR U5288 ( .A(n5084), .B(n4976), .Z(n5083) );
  ANDN U5289 ( .B(n4934), .A(n5085), .Z(n4976) );
  XOR U5290 ( .A(n4936), .B(n4820), .Z(n4934) );
  NOR U5291 ( .A(n5086), .B(n4936), .Z(n5084) );
  XNOR U5292 ( .A(n4974), .B(n5087), .Z(n4852) );
  XNOR U5293 ( .A(n5088), .B(n5089), .Z(n5087) );
  NANDN U5294 ( .A(n4972), .B(n5090), .Z(n5089) );
  IV U5295 ( .A(n4877), .Z(n4979) );
  XNOR U5296 ( .A(n4974), .B(n5091), .Z(n4877) );
  XOR U5297 ( .A(n5092), .B(n4854), .Z(n5091) );
  OR U5298 ( .A(n5093), .B(n4984), .Z(n4854) );
  XOR U5299 ( .A(n4856), .B(n5094), .Z(n4984) );
  ANDN U5300 ( .B(n5095), .A(n4982), .Z(n5092) );
  XOR U5301 ( .A(n5096), .B(n5088), .Z(n4974) );
  OR U5302 ( .A(n4987), .B(n5097), .Z(n5088) );
  XOR U5303 ( .A(n4989), .B(n4972), .Z(n4987) );
  XOR U5304 ( .A(n5094), .B(n4820), .Z(n4972) );
  XNOR U5305 ( .A(n5098), .B(n5099), .Z(n4820) );
  NANDN U5306 ( .A(n5100), .B(n5101), .Z(n5099) );
  IV U5307 ( .A(n4982), .Z(n5094) );
  XNOR U5308 ( .A(n5102), .B(n5103), .Z(n4982) );
  NANDN U5309 ( .A(n5100), .B(n5104), .Z(n5103) );
  ANDN U5310 ( .B(n4989), .A(n5105), .Z(n5096) );
  XOR U5311 ( .A(n4936), .B(n4856), .Z(n4989) );
  XOR U5312 ( .A(n5106), .B(n5102), .Z(n4856) );
  NANDN U5313 ( .A(n5107), .B(n5108), .Z(n5102) );
  NANDN U5314 ( .A(n5107), .B(n5112), .Z(n5098) );
  XOR U5315 ( .A(n5113), .B(n5114), .Z(n5100) );
  XOR U5316 ( .A(n5115), .B(n5110), .Z(n5114) );
  XNOR U5317 ( .A(n5116), .B(n5117), .Z(n5113) );
  XNOR U5318 ( .A(n5118), .B(n5119), .Z(n5117) );
  ANDN U5319 ( .B(n5115), .A(n5110), .Z(n5118) );
  ANDN U5320 ( .B(n5115), .A(n5109), .Z(n5111) );
  XNOR U5321 ( .A(n5116), .B(n5120), .Z(n5109) );
  XOR U5322 ( .A(n5121), .B(n5119), .Z(n5120) );
  NAND U5323 ( .A(n5108), .B(n5112), .Z(n5119) );
  XNOR U5324 ( .A(n5104), .B(n5110), .Z(n5108) );
  XOR U5325 ( .A(n5122), .B(n5123), .Z(n5110) );
  XOR U5326 ( .A(n5124), .B(n5125), .Z(n5123) );
  XNOR U5327 ( .A(n5126), .B(n5127), .Z(n5122) );
  ANDN U5328 ( .B(n5128), .A(n4935), .Z(n5126) );
  AND U5329 ( .A(n5101), .B(n5104), .Z(n5121) );
  XNOR U5330 ( .A(n5101), .B(n5104), .Z(n5116) );
  XNOR U5331 ( .A(n5129), .B(n5130), .Z(n5104) );
  XNOR U5332 ( .A(n5131), .B(n5132), .Z(n5130) );
  XOR U5333 ( .A(n5124), .B(n5133), .Z(n5129) );
  XNOR U5334 ( .A(n5134), .B(n5127), .Z(n5133) );
  OR U5335 ( .A(n4933), .B(n5085), .Z(n5127) );
  XNOR U5336 ( .A(n5086), .B(n4978), .Z(n5085) );
  XNOR U5337 ( .A(n4935), .B(n5135), .Z(n4933) );
  NOR U5338 ( .A(n5135), .B(n4978), .Z(n5134) );
  XNOR U5339 ( .A(n5136), .B(n5137), .Z(n5101) );
  XNOR U5340 ( .A(n5138), .B(n5139), .Z(n5137) );
  XOR U5341 ( .A(n4968), .B(n5124), .Z(n5139) );
  XOR U5342 ( .A(n5128), .B(n5140), .Z(n5124) );
  XNOR U5343 ( .A(n4857), .B(n5141), .Z(n5136) );
  XNOR U5344 ( .A(n5142), .B(n5143), .Z(n5141) );
  ANDN U5345 ( .B(n4983), .A(n5144), .Z(n5142) );
  XNOR U5346 ( .A(n5145), .B(n5146), .Z(n5115) );
  XNOR U5347 ( .A(n5125), .B(n5147), .Z(n5146) );
  XNOR U5348 ( .A(n4983), .B(n5132), .Z(n5147) );
  XOR U5349 ( .A(n4978), .B(n5135), .Z(n5132) );
  XNOR U5350 ( .A(n5138), .B(n5148), .Z(n5125) );
  XNOR U5351 ( .A(n5149), .B(n5150), .Z(n5148) );
  NANDN U5352 ( .A(n4973), .B(n5090), .Z(n5150) );
  IV U5353 ( .A(n5131), .Z(n5138) );
  XNOR U5354 ( .A(n5151), .B(n5149), .Z(n5131) );
  NANDN U5355 ( .A(n5097), .B(n4988), .Z(n5149) );
  XOR U5356 ( .A(n4983), .B(n5135), .Z(n4973) );
  IV U5357 ( .A(n4819), .Z(n5135) );
  XOR U5358 ( .A(n5152), .B(n5153), .Z(n4819) );
  XNOR U5359 ( .A(n5154), .B(n5155), .Z(n5153) );
  XOR U5360 ( .A(n5105), .B(n5090), .Z(n5097) );
  XNOR U5361 ( .A(n5095), .B(n4978), .Z(n5090) );
  XNOR U5362 ( .A(n5155), .B(n5152), .Z(n4978) );
  ANDN U5363 ( .B(n4990), .A(n5105), .Z(n5151) );
  XNOR U5364 ( .A(n5156), .B(n5128), .Z(n5105) );
  IV U5365 ( .A(n5086), .Z(n5128) );
  XNOR U5366 ( .A(n5157), .B(n5158), .Z(n5086) );
  XNOR U5367 ( .A(n5159), .B(n5155), .Z(n5158) );
  XOR U5368 ( .A(n5160), .B(n5140), .Z(n4990) );
  XNOR U5369 ( .A(n5144), .B(n5161), .Z(n5145) );
  XNOR U5370 ( .A(n5162), .B(n5143), .Z(n5161) );
  OR U5371 ( .A(n4985), .B(n5093), .Z(n5143) );
  XOR U5372 ( .A(n4857), .B(n5095), .Z(n5093) );
  IV U5373 ( .A(n5144), .Z(n5095) );
  XOR U5374 ( .A(n4968), .B(n4983), .Z(n4985) );
  XNOR U5375 ( .A(n5140), .B(n5163), .Z(n4983) );
  XNOR U5376 ( .A(n5154), .B(n5157), .Z(n5163) );
  XNOR U5377 ( .A(state[18]), .B(key[18]), .Z(n5157) );
  IV U5378 ( .A(n4935), .Z(n5140) );
  XOR U5379 ( .A(n5164), .B(n5165), .Z(n4935) );
  XOR U5380 ( .A(n5155), .B(n5166), .Z(n5165) );
  IV U5381 ( .A(n5160), .Z(n4968) );
  ANDN U5382 ( .B(n5160), .A(n4857), .Z(n5162) );
  XOR U5383 ( .A(n5152), .B(n5167), .Z(n5160) );
  XNOR U5384 ( .A(n5155), .B(n5168), .Z(n5167) );
  XOR U5385 ( .A(n5156), .B(n5169), .Z(n5155) );
  XNOR U5386 ( .A(state[22]), .B(key[22]), .Z(n5169) );
  IV U5387 ( .A(n5164), .Z(n5152) );
  XOR U5388 ( .A(state[21]), .B(key[21]), .Z(n5164) );
  XOR U5389 ( .A(n5170), .B(n5171), .Z(n5144) );
  XOR U5390 ( .A(n5168), .B(n5166), .Z(n5171) );
  XOR U5391 ( .A(state[23]), .B(key[23]), .Z(n5166) );
  XNOR U5392 ( .A(state[20]), .B(key[20]), .Z(n5168) );
  XOR U5393 ( .A(n4857), .B(n5159), .Z(n5170) );
  XNOR U5394 ( .A(n5154), .B(n5172), .Z(n5159) );
  XNOR U5395 ( .A(state[19]), .B(key[19]), .Z(n5172) );
  XNOR U5396 ( .A(state[17]), .B(key[17]), .Z(n5154) );
  IV U5397 ( .A(n5156), .Z(n4857) );
  XOR U5398 ( .A(state[16]), .B(key[16]), .Z(n5156) );
  XNOR U5399 ( .A(n4881), .B(n5173), .Z(n4887) );
  XNOR U5400 ( .A(n5174), .B(n5175), .Z(n5173) );
  NOR U5401 ( .A(n5176), .B(n4915), .Z(n5174) );
  XNOR U5402 ( .A(n5177), .B(n5178), .Z(n4881) );
  XNOR U5403 ( .A(n5179), .B(n5180), .Z(n5178) );
  NANDN U5404 ( .A(n5181), .B(n5182), .Z(n5180) );
  XNOR U5405 ( .A(n1034), .B(n1039), .Z(n413) );
  XOR U5406 ( .A(n4834), .B(n5183), .Z(n1039) );
  XNOR U5407 ( .A(n4836), .B(n4821), .Z(n5183) );
  XOR U5408 ( .A(n4991), .B(n4916), .Z(n4821) );
  XNOR U5409 ( .A(n4880), .B(n5184), .Z(n4916) );
  XNOR U5410 ( .A(n5185), .B(n5186), .Z(n5184) );
  NANDN U5411 ( .A(n5187), .B(n5188), .Z(n5186) );
  XNOR U5412 ( .A(n5177), .B(n5189), .Z(n4991) );
  XOR U5413 ( .A(n5190), .B(n4883), .Z(n5189) );
  OR U5414 ( .A(n5191), .B(n5192), .Z(n4883) );
  ANDN U5415 ( .B(n5193), .A(n5187), .Z(n5190) );
  XOR U5416 ( .A(n5177), .B(n5194), .Z(n4836) );
  XOR U5417 ( .A(n5175), .B(n5195), .Z(n5194) );
  OR U5418 ( .A(n5196), .B(n4892), .Z(n5195) );
  ANDN U5419 ( .B(n4913), .A(n5197), .Z(n5175) );
  XOR U5420 ( .A(n4915), .B(n4892), .Z(n4913) );
  XOR U5421 ( .A(n5198), .B(n5179), .Z(n5177) );
  OR U5422 ( .A(n5199), .B(n5200), .Z(n5179) );
  ANDN U5423 ( .B(n5201), .A(n5202), .Z(n5198) );
  XOR U5424 ( .A(n4909), .B(n5203), .Z(n4834) );
  XNOR U5425 ( .A(n5185), .B(n5204), .Z(n5203) );
  OR U5426 ( .A(n4885), .B(n5205), .Z(n5204) );
  OR U5427 ( .A(n5192), .B(n5206), .Z(n5185) );
  XOR U5428 ( .A(n4885), .B(n5207), .Z(n5192) );
  XNOR U5429 ( .A(n4880), .B(n5208), .Z(n4909) );
  XNOR U5430 ( .A(n5209), .B(n5210), .Z(n5208) );
  OR U5431 ( .A(n5181), .B(n5211), .Z(n5210) );
  XOR U5432 ( .A(n5212), .B(n5209), .Z(n4880) );
  NANDN U5433 ( .A(n5199), .B(n5213), .Z(n5209) );
  XOR U5434 ( .A(n5201), .B(n5181), .Z(n5199) );
  XOR U5435 ( .A(n5207), .B(n4892), .Z(n5181) );
  XNOR U5436 ( .A(n5214), .B(n5215), .Z(n4892) );
  NANDN U5437 ( .A(n5216), .B(n5217), .Z(n5215) );
  IV U5438 ( .A(n5187), .Z(n5207) );
  XNOR U5439 ( .A(n5218), .B(n5219), .Z(n5187) );
  NANDN U5440 ( .A(n5216), .B(n5220), .Z(n5219) );
  AND U5441 ( .A(n5201), .B(n5221), .Z(n5212) );
  XOR U5442 ( .A(n4915), .B(n4885), .Z(n5201) );
  XOR U5443 ( .A(n5222), .B(n5218), .Z(n4885) );
  NANDN U5444 ( .A(n5223), .B(n5224), .Z(n5218) );
  NANDN U5445 ( .A(n5223), .B(n5228), .Z(n5214) );
  XOR U5446 ( .A(n5229), .B(n5230), .Z(n5216) );
  XOR U5447 ( .A(n5231), .B(n5226), .Z(n5230) );
  XNOR U5448 ( .A(n5232), .B(n5233), .Z(n5229) );
  XNOR U5449 ( .A(n5234), .B(n5235), .Z(n5233) );
  ANDN U5450 ( .B(n5231), .A(n5226), .Z(n5234) );
  ANDN U5451 ( .B(n5231), .A(n5225), .Z(n5227) );
  XNOR U5452 ( .A(n5232), .B(n5236), .Z(n5225) );
  XOR U5453 ( .A(n5237), .B(n5235), .Z(n5236) );
  NAND U5454 ( .A(n5224), .B(n5228), .Z(n5235) );
  XNOR U5455 ( .A(n5220), .B(n5226), .Z(n5224) );
  XOR U5456 ( .A(n5238), .B(n5239), .Z(n5226) );
  XOR U5457 ( .A(n5240), .B(n5241), .Z(n5239) );
  XNOR U5458 ( .A(n5242), .B(n5243), .Z(n5238) );
  ANDN U5459 ( .B(n5244), .A(n4914), .Z(n5242) );
  AND U5460 ( .A(n5217), .B(n5220), .Z(n5237) );
  XNOR U5461 ( .A(n5217), .B(n5220), .Z(n5232) );
  XNOR U5462 ( .A(n5245), .B(n5246), .Z(n5220) );
  XNOR U5463 ( .A(n5247), .B(n5248), .Z(n5246) );
  XOR U5464 ( .A(n5240), .B(n5249), .Z(n5245) );
  XNOR U5465 ( .A(n5250), .B(n5243), .Z(n5249) );
  OR U5466 ( .A(n4912), .B(n5197), .Z(n5243) );
  XNOR U5467 ( .A(n5176), .B(n5196), .Z(n5197) );
  XNOR U5468 ( .A(n4914), .B(n5251), .Z(n4912) );
  NOR U5469 ( .A(n5251), .B(n5196), .Z(n5250) );
  XNOR U5470 ( .A(n5252), .B(n5253), .Z(n5217) );
  XNOR U5471 ( .A(n5254), .B(n5255), .Z(n5253) );
  XOR U5472 ( .A(n5205), .B(n5240), .Z(n5255) );
  XOR U5473 ( .A(n5244), .B(n5256), .Z(n5240) );
  XNOR U5474 ( .A(n4886), .B(n5257), .Z(n5252) );
  XNOR U5475 ( .A(n5258), .B(n5259), .Z(n5257) );
  ANDN U5476 ( .B(n5188), .A(n5260), .Z(n5258) );
  XNOR U5477 ( .A(n5261), .B(n5262), .Z(n5231) );
  XNOR U5478 ( .A(n5241), .B(n5263), .Z(n5262) );
  XNOR U5479 ( .A(n5188), .B(n5248), .Z(n5263) );
  XOR U5480 ( .A(n5196), .B(n5251), .Z(n5248) );
  XNOR U5481 ( .A(n5254), .B(n5264), .Z(n5241) );
  XNOR U5482 ( .A(n5265), .B(n5266), .Z(n5264) );
  NANDN U5483 ( .A(n5211), .B(n5182), .Z(n5266) );
  IV U5484 ( .A(n5247), .Z(n5254) );
  XNOR U5485 ( .A(n5267), .B(n5265), .Z(n5247) );
  NANDN U5486 ( .A(n5200), .B(n5213), .Z(n5265) );
  XOR U5487 ( .A(n5188), .B(n5251), .Z(n5211) );
  IV U5488 ( .A(n4891), .Z(n5251) );
  XOR U5489 ( .A(n5268), .B(n5269), .Z(n4891) );
  XNOR U5490 ( .A(n5270), .B(n5271), .Z(n5269) );
  XOR U5491 ( .A(n5202), .B(n5182), .Z(n5200) );
  XNOR U5492 ( .A(n5193), .B(n5196), .Z(n5182) );
  XNOR U5493 ( .A(n5271), .B(n5268), .Z(n5196) );
  ANDN U5494 ( .B(n5221), .A(n5202), .Z(n5267) );
  XNOR U5495 ( .A(n5272), .B(n5244), .Z(n5202) );
  IV U5496 ( .A(n5176), .Z(n5244) );
  XNOR U5497 ( .A(n5273), .B(n5274), .Z(n5176) );
  XNOR U5498 ( .A(n5275), .B(n5271), .Z(n5274) );
  XOR U5499 ( .A(n5276), .B(n5256), .Z(n5221) );
  XNOR U5500 ( .A(n5260), .B(n5277), .Z(n5261) );
  XNOR U5501 ( .A(n5278), .B(n5259), .Z(n5277) );
  OR U5502 ( .A(n5206), .B(n5191), .Z(n5259) );
  XOR U5503 ( .A(n4886), .B(n5193), .Z(n5191) );
  IV U5504 ( .A(n5260), .Z(n5193) );
  XOR U5505 ( .A(n5205), .B(n5188), .Z(n5206) );
  XNOR U5506 ( .A(n5256), .B(n5279), .Z(n5188) );
  XNOR U5507 ( .A(n5270), .B(n5273), .Z(n5279) );
  XNOR U5508 ( .A(state[58]), .B(key[58]), .Z(n5273) );
  IV U5509 ( .A(n4914), .Z(n5256) );
  XOR U5510 ( .A(n5280), .B(n5281), .Z(n4914) );
  XOR U5511 ( .A(n5271), .B(n5282), .Z(n5281) );
  IV U5512 ( .A(n5276), .Z(n5205) );
  ANDN U5513 ( .B(n5276), .A(n4886), .Z(n5278) );
  XOR U5514 ( .A(n5268), .B(n5283), .Z(n5276) );
  XNOR U5515 ( .A(n5271), .B(n5284), .Z(n5283) );
  XOR U5516 ( .A(n5272), .B(n5285), .Z(n5271) );
  XNOR U5517 ( .A(state[62]), .B(key[62]), .Z(n5285) );
  IV U5518 ( .A(n5280), .Z(n5268) );
  XOR U5519 ( .A(state[61]), .B(key[61]), .Z(n5280) );
  XOR U5520 ( .A(n5286), .B(n5287), .Z(n5260) );
  XOR U5521 ( .A(n5284), .B(n5282), .Z(n5287) );
  XOR U5522 ( .A(state[63]), .B(key[63]), .Z(n5282) );
  XNOR U5523 ( .A(state[60]), .B(key[60]), .Z(n5284) );
  XOR U5524 ( .A(n4886), .B(n5275), .Z(n5286) );
  XNOR U5525 ( .A(n5270), .B(n5288), .Z(n5275) );
  XNOR U5526 ( .A(state[59]), .B(key[59]), .Z(n5288) );
  XNOR U5527 ( .A(state[57]), .B(key[57]), .Z(n5270) );
  IV U5528 ( .A(n5272), .Z(n4886) );
  XOR U5529 ( .A(state[56]), .B(key[56]), .Z(n5272) );
  XOR U5530 ( .A(n4780), .B(n5289), .Z(n1034) );
  XNOR U5531 ( .A(n4782), .B(n4798), .Z(n5289) );
  XOR U5532 ( .A(n4901), .B(n5290), .Z(n4896) );
  XOR U5533 ( .A(n5291), .B(n4871), .Z(n5290) );
  OR U5534 ( .A(n5292), .B(n5293), .Z(n4871) );
  ANDN U5535 ( .B(n5294), .A(n5295), .Z(n5291) );
  XNOR U5536 ( .A(n4862), .B(n5296), .Z(n4783) );
  XNOR U5537 ( .A(n5297), .B(n5298), .Z(n5296) );
  NANDN U5538 ( .A(n5295), .B(n5299), .Z(n5298) );
  XOR U5539 ( .A(n4901), .B(n5300), .Z(n4782) );
  XNOR U5540 ( .A(n4899), .B(n5301), .Z(n5300) );
  OR U5541 ( .A(n5302), .B(n4867), .Z(n5301) );
  OR U5542 ( .A(n5303), .B(n4868), .Z(n4899) );
  XNOR U5543 ( .A(n4828), .B(n4867), .Z(n4868) );
  XOR U5544 ( .A(n5304), .B(n4903), .Z(n4901) );
  OR U5545 ( .A(n5305), .B(n5306), .Z(n4903) );
  ANDN U5546 ( .B(n5307), .A(n5308), .Z(n5304) );
  XOR U5547 ( .A(n4823), .B(n5309), .Z(n4780) );
  XNOR U5548 ( .A(n5297), .B(n5310), .Z(n5309) );
  OR U5549 ( .A(n4873), .B(n5311), .Z(n5310) );
  OR U5550 ( .A(n5293), .B(n5312), .Z(n5297) );
  XOR U5551 ( .A(n4873), .B(n5313), .Z(n5293) );
  XNOR U5552 ( .A(n4862), .B(n5314), .Z(n4823) );
  XNOR U5553 ( .A(n5315), .B(n5316), .Z(n5314) );
  OR U5554 ( .A(n4905), .B(n5317), .Z(n5316) );
  XOR U5555 ( .A(n5318), .B(n5315), .Z(n4862) );
  NANDN U5556 ( .A(n5305), .B(n5319), .Z(n5315) );
  XOR U5557 ( .A(n5307), .B(n4905), .Z(n5305) );
  XOR U5558 ( .A(n5313), .B(n4867), .Z(n4905) );
  XNOR U5559 ( .A(n5320), .B(n5321), .Z(n4867) );
  NANDN U5560 ( .A(n5322), .B(n5323), .Z(n5321) );
  IV U5561 ( .A(n5295), .Z(n5313) );
  XNOR U5562 ( .A(n5324), .B(n5325), .Z(n5295) );
  NANDN U5563 ( .A(n5322), .B(n5326), .Z(n5325) );
  AND U5564 ( .A(n5307), .B(n5327), .Z(n5318) );
  XOR U5565 ( .A(n4828), .B(n4873), .Z(n5307) );
  XOR U5566 ( .A(n5328), .B(n5324), .Z(n4873) );
  NANDN U5567 ( .A(n5329), .B(n5330), .Z(n5324) );
  NANDN U5568 ( .A(n5329), .B(n5334), .Z(n5320) );
  XOR U5569 ( .A(n5335), .B(n5336), .Z(n5322) );
  XOR U5570 ( .A(n5337), .B(n5332), .Z(n5336) );
  XNOR U5571 ( .A(n5338), .B(n5339), .Z(n5335) );
  XNOR U5572 ( .A(n5340), .B(n5341), .Z(n5339) );
  ANDN U5573 ( .B(n5337), .A(n5332), .Z(n5340) );
  ANDN U5574 ( .B(n5337), .A(n5331), .Z(n5333) );
  XNOR U5575 ( .A(n5338), .B(n5342), .Z(n5331) );
  XOR U5576 ( .A(n5343), .B(n5341), .Z(n5342) );
  NAND U5577 ( .A(n5330), .B(n5334), .Z(n5341) );
  XNOR U5578 ( .A(n5326), .B(n5332), .Z(n5330) );
  XOR U5579 ( .A(n5344), .B(n5345), .Z(n5332) );
  XOR U5580 ( .A(n5346), .B(n5347), .Z(n5345) );
  XNOR U5581 ( .A(n5348), .B(n5349), .Z(n5344) );
  ANDN U5582 ( .B(n5350), .A(n4827), .Z(n5348) );
  AND U5583 ( .A(n5323), .B(n5326), .Z(n5343) );
  XNOR U5584 ( .A(n5323), .B(n5326), .Z(n5338) );
  XNOR U5585 ( .A(n5351), .B(n5352), .Z(n5326) );
  XNOR U5586 ( .A(n5353), .B(n5354), .Z(n5352) );
  XOR U5587 ( .A(n5346), .B(n5355), .Z(n5351) );
  XNOR U5588 ( .A(n5356), .B(n5349), .Z(n5355) );
  OR U5589 ( .A(n4869), .B(n5303), .Z(n5349) );
  XNOR U5590 ( .A(n4900), .B(n5302), .Z(n5303) );
  XNOR U5591 ( .A(n4827), .B(n5357), .Z(n4869) );
  NOR U5592 ( .A(n5357), .B(n5302), .Z(n5356) );
  XNOR U5593 ( .A(n5358), .B(n5359), .Z(n5323) );
  XNOR U5594 ( .A(n5360), .B(n5361), .Z(n5359) );
  XOR U5595 ( .A(n5311), .B(n5346), .Z(n5361) );
  XOR U5596 ( .A(n5350), .B(n5362), .Z(n5346) );
  XNOR U5597 ( .A(n4874), .B(n5363), .Z(n5358) );
  XNOR U5598 ( .A(n5364), .B(n5365), .Z(n5363) );
  ANDN U5599 ( .B(n5299), .A(n5366), .Z(n5364) );
  XNOR U5600 ( .A(n5367), .B(n5368), .Z(n5337) );
  XNOR U5601 ( .A(n5347), .B(n5369), .Z(n5368) );
  XNOR U5602 ( .A(n5299), .B(n5354), .Z(n5369) );
  XOR U5603 ( .A(n5302), .B(n5357), .Z(n5354) );
  XNOR U5604 ( .A(n5360), .B(n5370), .Z(n5347) );
  XNOR U5605 ( .A(n5371), .B(n5372), .Z(n5370) );
  NANDN U5606 ( .A(n5317), .B(n4906), .Z(n5372) );
  IV U5607 ( .A(n5353), .Z(n5360) );
  XNOR U5608 ( .A(n5373), .B(n5371), .Z(n5353) );
  NANDN U5609 ( .A(n5306), .B(n5319), .Z(n5371) );
  XOR U5610 ( .A(n5299), .B(n5357), .Z(n5317) );
  IV U5611 ( .A(n4866), .Z(n5357) );
  XOR U5612 ( .A(n5374), .B(n5375), .Z(n4866) );
  XNOR U5613 ( .A(n5376), .B(n5377), .Z(n5375) );
  XOR U5614 ( .A(n5308), .B(n4906), .Z(n5306) );
  XNOR U5615 ( .A(n5294), .B(n5302), .Z(n4906) );
  XNOR U5616 ( .A(n5377), .B(n5374), .Z(n5302) );
  ANDN U5617 ( .B(n5327), .A(n5308), .Z(n5373) );
  XNOR U5618 ( .A(n5378), .B(n5350), .Z(n5308) );
  IV U5619 ( .A(n4900), .Z(n5350) );
  XNOR U5620 ( .A(n5379), .B(n5380), .Z(n4900) );
  XNOR U5621 ( .A(n5381), .B(n5377), .Z(n5380) );
  XOR U5622 ( .A(n5382), .B(n5362), .Z(n5327) );
  XNOR U5623 ( .A(n5366), .B(n5383), .Z(n5367) );
  XNOR U5624 ( .A(n5384), .B(n5365), .Z(n5383) );
  OR U5625 ( .A(n5312), .B(n5292), .Z(n5365) );
  XOR U5626 ( .A(n4874), .B(n5294), .Z(n5292) );
  IV U5627 ( .A(n5366), .Z(n5294) );
  XOR U5628 ( .A(n5311), .B(n5299), .Z(n5312) );
  XNOR U5629 ( .A(n5362), .B(n5385), .Z(n5299) );
  XNOR U5630 ( .A(n5376), .B(n5379), .Z(n5385) );
  XNOR U5631 ( .A(state[66]), .B(key[66]), .Z(n5379) );
  IV U5632 ( .A(n4827), .Z(n5362) );
  XOR U5633 ( .A(n5386), .B(n5387), .Z(n4827) );
  XOR U5634 ( .A(n5377), .B(n5388), .Z(n5387) );
  IV U5635 ( .A(n5382), .Z(n5311) );
  ANDN U5636 ( .B(n5382), .A(n4874), .Z(n5384) );
  XOR U5637 ( .A(n5374), .B(n5389), .Z(n5382) );
  XNOR U5638 ( .A(n5377), .B(n5390), .Z(n5389) );
  XOR U5639 ( .A(n5378), .B(n5391), .Z(n5377) );
  XNOR U5640 ( .A(state[70]), .B(key[70]), .Z(n5391) );
  IV U5641 ( .A(n5386), .Z(n5374) );
  XOR U5642 ( .A(state[69]), .B(key[69]), .Z(n5386) );
  XOR U5643 ( .A(n5392), .B(n5393), .Z(n5366) );
  XOR U5644 ( .A(n5390), .B(n5388), .Z(n5393) );
  XOR U5645 ( .A(state[71]), .B(key[71]), .Z(n5388) );
  XNOR U5646 ( .A(state[68]), .B(key[68]), .Z(n5390) );
  XOR U5647 ( .A(n4874), .B(n5381), .Z(n5392) );
  XNOR U5648 ( .A(n5376), .B(n5394), .Z(n5381) );
  XNOR U5649 ( .A(state[67]), .B(key[67]), .Z(n5394) );
  XNOR U5650 ( .A(state[65]), .B(key[65]), .Z(n5376) );
  IV U5651 ( .A(n5378), .Z(n4874) );
  XOR U5652 ( .A(state[64]), .B(key[64]), .Z(n5378) );
endmodule

