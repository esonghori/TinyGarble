
module compare_N16384_CC64 ( clk, rst, x, y, g, e );
  input [255:0] x;
  input [255:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  IV U10 ( .A(ebreg), .Z(e) );
  XNOR U11 ( .A(y[189]), .B(x[189]), .Z(n9) );
  NANDN U12 ( .A(x[188]), .B(y[188]), .Z(n8) );
  NAND U13 ( .A(n9), .B(n8), .Z(n1085) );
  XNOR U14 ( .A(y[185]), .B(x[185]), .Z(n11) );
  NANDN U15 ( .A(x[184]), .B(y[184]), .Z(n10) );
  NAND U16 ( .A(n11), .B(n10), .Z(n1073) );
  XNOR U17 ( .A(y[187]), .B(x[187]), .Z(n13) );
  NANDN U18 ( .A(x[186]), .B(y[186]), .Z(n12) );
  NAND U19 ( .A(n13), .B(n12), .Z(n1079) );
  NOR U20 ( .A(n1073), .B(n1079), .Z(n16) );
  XNOR U21 ( .A(y[191]), .B(x[191]), .Z(n15) );
  NANDN U22 ( .A(x[190]), .B(y[190]), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n1091) );
  ANDN U24 ( .B(n16), .A(n1091), .Z(n17) );
  NANDN U25 ( .A(n1085), .B(n17), .Z(n53) );
  XNOR U26 ( .A(y[173]), .B(x[173]), .Z(n19) );
  NANDN U27 ( .A(x[172]), .B(y[172]), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n1037) );
  XNOR U29 ( .A(y[169]), .B(x[169]), .Z(n21) );
  NANDN U30 ( .A(x[168]), .B(y[168]), .Z(n20) );
  NAND U31 ( .A(n21), .B(n20), .Z(n1025) );
  XNOR U32 ( .A(y[171]), .B(x[171]), .Z(n23) );
  NANDN U33 ( .A(x[170]), .B(y[170]), .Z(n22) );
  NAND U34 ( .A(n23), .B(n22), .Z(n1031) );
  NOR U35 ( .A(n1025), .B(n1031), .Z(n26) );
  XNOR U36 ( .A(y[175]), .B(x[175]), .Z(n25) );
  NANDN U37 ( .A(x[174]), .B(y[174]), .Z(n24) );
  NAND U38 ( .A(n25), .B(n24), .Z(n1043) );
  ANDN U39 ( .B(n26), .A(n1043), .Z(n27) );
  NANDN U40 ( .A(n1037), .B(n27), .Z(n39) );
  XNOR U41 ( .A(y[165]), .B(x[165]), .Z(n29) );
  NANDN U42 ( .A(x[164]), .B(y[164]), .Z(n28) );
  NAND U43 ( .A(n29), .B(n28), .Z(n1013) );
  XNOR U44 ( .A(y[161]), .B(x[161]), .Z(n31) );
  NANDN U45 ( .A(x[160]), .B(y[160]), .Z(n30) );
  NAND U46 ( .A(n31), .B(n30), .Z(n1001) );
  XNOR U47 ( .A(y[163]), .B(x[163]), .Z(n33) );
  NANDN U48 ( .A(x[162]), .B(y[162]), .Z(n32) );
  NAND U49 ( .A(n33), .B(n32), .Z(n1007) );
  NOR U50 ( .A(n1001), .B(n1007), .Z(n36) );
  XNOR U51 ( .A(y[167]), .B(x[167]), .Z(n35) );
  NANDN U52 ( .A(x[166]), .B(y[166]), .Z(n34) );
  NAND U53 ( .A(n35), .B(n34), .Z(n1019) );
  ANDN U54 ( .B(n36), .A(n1019), .Z(n37) );
  NANDN U55 ( .A(n1013), .B(n37), .Z(n38) );
  NOR U56 ( .A(n39), .B(n38), .Z(n51) );
  XNOR U57 ( .A(y[181]), .B(x[181]), .Z(n41) );
  NANDN U58 ( .A(x[180]), .B(y[180]), .Z(n40) );
  NAND U59 ( .A(n41), .B(n40), .Z(n1061) );
  XNOR U60 ( .A(y[177]), .B(x[177]), .Z(n43) );
  NANDN U61 ( .A(x[176]), .B(y[176]), .Z(n42) );
  NAND U62 ( .A(n43), .B(n42), .Z(n1049) );
  XNOR U63 ( .A(y[179]), .B(x[179]), .Z(n45) );
  NANDN U64 ( .A(x[178]), .B(y[178]), .Z(n44) );
  NAND U65 ( .A(n45), .B(n44), .Z(n1055) );
  NOR U66 ( .A(n1049), .B(n1055), .Z(n48) );
  XNOR U67 ( .A(y[183]), .B(x[183]), .Z(n47) );
  NANDN U68 ( .A(x[182]), .B(y[182]), .Z(n46) );
  NAND U69 ( .A(n47), .B(n46), .Z(n1067) );
  ANDN U70 ( .B(n48), .A(n1067), .Z(n49) );
  NANDN U71 ( .A(n1061), .B(n49), .Z(n50) );
  ANDN U72 ( .B(n51), .A(n50), .Z(n52) );
  NANDN U73 ( .A(n53), .B(n52), .Z(n101) );
  XNOR U74 ( .A(y[157]), .B(x[157]), .Z(n55) );
  NANDN U75 ( .A(x[156]), .B(y[156]), .Z(n54) );
  NAND U76 ( .A(n55), .B(n54), .Z(n989) );
  XNOR U77 ( .A(y[153]), .B(x[153]), .Z(n57) );
  NANDN U78 ( .A(x[152]), .B(y[152]), .Z(n56) );
  NAND U79 ( .A(n57), .B(n56), .Z(n977) );
  XNOR U80 ( .A(y[155]), .B(x[155]), .Z(n59) );
  NANDN U81 ( .A(x[154]), .B(y[154]), .Z(n58) );
  NAND U82 ( .A(n59), .B(n58), .Z(n983) );
  NOR U83 ( .A(n977), .B(n983), .Z(n62) );
  XNOR U84 ( .A(y[159]), .B(x[159]), .Z(n61) );
  NANDN U85 ( .A(x[158]), .B(y[158]), .Z(n60) );
  NAND U86 ( .A(n61), .B(n60), .Z(n995) );
  ANDN U87 ( .B(n62), .A(n995), .Z(n63) );
  NANDN U88 ( .A(n989), .B(n63), .Z(n99) );
  XNOR U89 ( .A(y[141]), .B(x[141]), .Z(n65) );
  NANDN U90 ( .A(x[140]), .B(y[140]), .Z(n64) );
  NAND U91 ( .A(n65), .B(n64), .Z(n941) );
  XNOR U92 ( .A(y[137]), .B(x[137]), .Z(n67) );
  NANDN U93 ( .A(x[136]), .B(y[136]), .Z(n66) );
  NAND U94 ( .A(n67), .B(n66), .Z(n929) );
  XNOR U95 ( .A(y[139]), .B(x[139]), .Z(n69) );
  NANDN U96 ( .A(x[138]), .B(y[138]), .Z(n68) );
  NAND U97 ( .A(n69), .B(n68), .Z(n935) );
  NOR U98 ( .A(n929), .B(n935), .Z(n72) );
  XNOR U99 ( .A(y[143]), .B(x[143]), .Z(n71) );
  NANDN U100 ( .A(x[142]), .B(y[142]), .Z(n70) );
  NAND U101 ( .A(n71), .B(n70), .Z(n947) );
  ANDN U102 ( .B(n72), .A(n947), .Z(n73) );
  NANDN U103 ( .A(n941), .B(n73), .Z(n85) );
  XNOR U104 ( .A(y[133]), .B(x[133]), .Z(n75) );
  NANDN U105 ( .A(x[132]), .B(y[132]), .Z(n74) );
  NAND U106 ( .A(n75), .B(n74), .Z(n917) );
  XNOR U107 ( .A(y[129]), .B(x[129]), .Z(n77) );
  NANDN U108 ( .A(x[128]), .B(y[128]), .Z(n76) );
  NAND U109 ( .A(n77), .B(n76), .Z(n905) );
  XNOR U110 ( .A(y[131]), .B(x[131]), .Z(n79) );
  NANDN U111 ( .A(x[130]), .B(y[130]), .Z(n78) );
  NAND U112 ( .A(n79), .B(n78), .Z(n911) );
  NOR U113 ( .A(n905), .B(n911), .Z(n82) );
  XNOR U114 ( .A(y[135]), .B(x[135]), .Z(n81) );
  NANDN U115 ( .A(x[134]), .B(y[134]), .Z(n80) );
  NAND U116 ( .A(n81), .B(n80), .Z(n923) );
  ANDN U117 ( .B(n82), .A(n923), .Z(n83) );
  NANDN U118 ( .A(n917), .B(n83), .Z(n84) );
  NOR U119 ( .A(n85), .B(n84), .Z(n97) );
  XNOR U120 ( .A(y[149]), .B(x[149]), .Z(n87) );
  NANDN U121 ( .A(x[148]), .B(y[148]), .Z(n86) );
  NAND U122 ( .A(n87), .B(n86), .Z(n965) );
  XNOR U123 ( .A(y[145]), .B(x[145]), .Z(n89) );
  NANDN U124 ( .A(x[144]), .B(y[144]), .Z(n88) );
  NAND U125 ( .A(n89), .B(n88), .Z(n953) );
  XNOR U126 ( .A(y[147]), .B(x[147]), .Z(n91) );
  NANDN U127 ( .A(x[146]), .B(y[146]), .Z(n90) );
  NAND U128 ( .A(n91), .B(n90), .Z(n959) );
  NOR U129 ( .A(n953), .B(n959), .Z(n94) );
  XNOR U130 ( .A(y[151]), .B(x[151]), .Z(n93) );
  NANDN U131 ( .A(x[150]), .B(y[150]), .Z(n92) );
  NAND U132 ( .A(n93), .B(n92), .Z(n971) );
  ANDN U133 ( .B(n94), .A(n971), .Z(n95) );
  NANDN U134 ( .A(n965), .B(n95), .Z(n96) );
  ANDN U135 ( .B(n97), .A(n96), .Z(n98) );
  NANDN U136 ( .A(n99), .B(n98), .Z(n100) );
  NOR U137 ( .A(n101), .B(n100), .Z(n325) );
  ANDN U138 ( .B(x[252]), .A(y[252]), .Z(n1273) );
  ANDN U139 ( .B(x[248]), .A(y[248]), .Z(n1261) );
  ANDN U140 ( .B(x[250]), .A(y[250]), .Z(n1267) );
  NOR U141 ( .A(n1261), .B(n1267), .Z(n102) );
  ANDN U142 ( .B(x[254]), .A(y[254]), .Z(n1279) );
  ANDN U143 ( .B(n102), .A(n1279), .Z(n103) );
  NANDN U144 ( .A(n1273), .B(n103), .Z(n115) );
  ANDN U145 ( .B(x[236]), .A(y[236]), .Z(n1225) );
  ANDN U146 ( .B(x[232]), .A(y[232]), .Z(n1213) );
  ANDN U147 ( .B(x[234]), .A(y[234]), .Z(n1219) );
  NOR U148 ( .A(n1213), .B(n1219), .Z(n104) );
  ANDN U149 ( .B(x[238]), .A(y[238]), .Z(n1231) );
  ANDN U150 ( .B(n104), .A(n1231), .Z(n105) );
  NANDN U151 ( .A(n1225), .B(n105), .Z(n109) );
  ANDN U152 ( .B(x[228]), .A(y[228]), .Z(n1201) );
  ANDN U153 ( .B(x[224]), .A(y[224]), .Z(n1189) );
  ANDN U154 ( .B(x[226]), .A(y[226]), .Z(n1195) );
  NOR U155 ( .A(n1189), .B(n1195), .Z(n106) );
  ANDN U156 ( .B(x[230]), .A(y[230]), .Z(n1207) );
  ANDN U157 ( .B(n106), .A(n1207), .Z(n107) );
  NANDN U158 ( .A(n1201), .B(n107), .Z(n108) );
  NOR U159 ( .A(n109), .B(n108), .Z(n113) );
  ANDN U160 ( .B(x[244]), .A(y[244]), .Z(n1249) );
  ANDN U161 ( .B(x[240]), .A(y[240]), .Z(n1237) );
  ANDN U162 ( .B(x[242]), .A(y[242]), .Z(n1243) );
  NOR U163 ( .A(n1237), .B(n1243), .Z(n110) );
  ANDN U164 ( .B(x[246]), .A(y[246]), .Z(n1255) );
  ANDN U165 ( .B(n110), .A(n1255), .Z(n111) );
  NANDN U166 ( .A(n1249), .B(n111), .Z(n112) );
  ANDN U167 ( .B(n113), .A(n112), .Z(n114) );
  NANDN U168 ( .A(n115), .B(n114), .Z(n163) );
  ANDN U169 ( .B(x[188]), .A(y[188]), .Z(n1081) );
  ANDN U170 ( .B(x[184]), .A(y[184]), .Z(n1069) );
  ANDN U171 ( .B(x[186]), .A(y[186]), .Z(n1075) );
  NOR U172 ( .A(n1069), .B(n1075), .Z(n116) );
  ANDN U173 ( .B(x[190]), .A(y[190]), .Z(n1087) );
  ANDN U174 ( .B(n116), .A(n1087), .Z(n117) );
  NANDN U175 ( .A(n1081), .B(n117), .Z(n129) );
  ANDN U176 ( .B(x[172]), .A(y[172]), .Z(n1033) );
  ANDN U177 ( .B(x[168]), .A(y[168]), .Z(n1021) );
  ANDN U178 ( .B(x[170]), .A(y[170]), .Z(n1027) );
  NOR U179 ( .A(n1021), .B(n1027), .Z(n118) );
  ANDN U180 ( .B(x[174]), .A(y[174]), .Z(n1039) );
  ANDN U181 ( .B(n118), .A(n1039), .Z(n119) );
  NANDN U182 ( .A(n1033), .B(n119), .Z(n123) );
  ANDN U183 ( .B(x[164]), .A(y[164]), .Z(n1009) );
  ANDN U184 ( .B(x[160]), .A(y[160]), .Z(n997) );
  ANDN U185 ( .B(x[162]), .A(y[162]), .Z(n1003) );
  NOR U186 ( .A(n997), .B(n1003), .Z(n120) );
  ANDN U187 ( .B(x[166]), .A(y[166]), .Z(n1015) );
  ANDN U188 ( .B(n120), .A(n1015), .Z(n121) );
  NANDN U189 ( .A(n1009), .B(n121), .Z(n122) );
  NOR U190 ( .A(n123), .B(n122), .Z(n127) );
  ANDN U191 ( .B(x[180]), .A(y[180]), .Z(n1057) );
  ANDN U192 ( .B(x[176]), .A(y[176]), .Z(n1045) );
  ANDN U193 ( .B(x[178]), .A(y[178]), .Z(n1051) );
  NOR U194 ( .A(n1045), .B(n1051), .Z(n124) );
  ANDN U195 ( .B(x[182]), .A(y[182]), .Z(n1063) );
  ANDN U196 ( .B(n124), .A(n1063), .Z(n125) );
  NANDN U197 ( .A(n1057), .B(n125), .Z(n126) );
  ANDN U198 ( .B(n127), .A(n126), .Z(n128) );
  NANDN U199 ( .A(n129), .B(n128), .Z(n145) );
  ANDN U200 ( .B(x[156]), .A(y[156]), .Z(n985) );
  ANDN U201 ( .B(x[152]), .A(y[152]), .Z(n973) );
  ANDN U202 ( .B(x[154]), .A(y[154]), .Z(n979) );
  NOR U203 ( .A(n973), .B(n979), .Z(n130) );
  ANDN U204 ( .B(x[158]), .A(y[158]), .Z(n991) );
  ANDN U205 ( .B(n130), .A(n991), .Z(n131) );
  NANDN U206 ( .A(n985), .B(n131), .Z(n143) );
  ANDN U207 ( .B(x[140]), .A(y[140]), .Z(n937) );
  ANDN U208 ( .B(x[136]), .A(y[136]), .Z(n925) );
  ANDN U209 ( .B(x[138]), .A(y[138]), .Z(n931) );
  NOR U210 ( .A(n925), .B(n931), .Z(n132) );
  ANDN U211 ( .B(x[142]), .A(y[142]), .Z(n943) );
  ANDN U212 ( .B(n132), .A(n943), .Z(n133) );
  NANDN U213 ( .A(n937), .B(n133), .Z(n137) );
  ANDN U214 ( .B(x[132]), .A(y[132]), .Z(n913) );
  ANDN U215 ( .B(x[128]), .A(y[128]), .Z(n903) );
  ANDN U216 ( .B(x[130]), .A(y[130]), .Z(n907) );
  NOR U217 ( .A(n903), .B(n907), .Z(n134) );
  ANDN U218 ( .B(x[134]), .A(y[134]), .Z(n919) );
  ANDN U219 ( .B(n134), .A(n919), .Z(n135) );
  NANDN U220 ( .A(n913), .B(n135), .Z(n136) );
  NOR U221 ( .A(n137), .B(n136), .Z(n141) );
  ANDN U222 ( .B(x[148]), .A(y[148]), .Z(n961) );
  ANDN U223 ( .B(x[144]), .A(y[144]), .Z(n949) );
  ANDN U224 ( .B(x[146]), .A(y[146]), .Z(n955) );
  NOR U225 ( .A(n949), .B(n955), .Z(n138) );
  ANDN U226 ( .B(x[150]), .A(y[150]), .Z(n967) );
  ANDN U227 ( .B(n138), .A(n967), .Z(n139) );
  NANDN U228 ( .A(n961), .B(n139), .Z(n140) );
  ANDN U229 ( .B(n141), .A(n140), .Z(n142) );
  NANDN U230 ( .A(n143), .B(n142), .Z(n144) );
  NOR U231 ( .A(n145), .B(n144), .Z(n161) );
  ANDN U232 ( .B(x[220]), .A(y[220]), .Z(n1177) );
  ANDN U233 ( .B(x[216]), .A(y[216]), .Z(n1165) );
  ANDN U234 ( .B(x[218]), .A(y[218]), .Z(n1171) );
  NOR U235 ( .A(n1165), .B(n1171), .Z(n146) );
  ANDN U236 ( .B(x[222]), .A(y[222]), .Z(n1183) );
  ANDN U237 ( .B(n146), .A(n1183), .Z(n147) );
  NANDN U238 ( .A(n1177), .B(n147), .Z(n159) );
  ANDN U239 ( .B(x[204]), .A(y[204]), .Z(n1129) );
  ANDN U240 ( .B(x[200]), .A(y[200]), .Z(n1117) );
  ANDN U241 ( .B(x[202]), .A(y[202]), .Z(n1123) );
  NOR U242 ( .A(n1117), .B(n1123), .Z(n148) );
  ANDN U243 ( .B(x[206]), .A(y[206]), .Z(n1135) );
  ANDN U244 ( .B(n148), .A(n1135), .Z(n149) );
  NANDN U245 ( .A(n1129), .B(n149), .Z(n153) );
  ANDN U246 ( .B(x[196]), .A(y[196]), .Z(n1105) );
  ANDN U247 ( .B(x[192]), .A(y[192]), .Z(n1093) );
  ANDN U248 ( .B(x[194]), .A(y[194]), .Z(n1099) );
  NOR U249 ( .A(n1093), .B(n1099), .Z(n150) );
  ANDN U250 ( .B(x[198]), .A(y[198]), .Z(n1111) );
  ANDN U251 ( .B(n150), .A(n1111), .Z(n151) );
  NANDN U252 ( .A(n1105), .B(n151), .Z(n152) );
  NOR U253 ( .A(n153), .B(n152), .Z(n157) );
  ANDN U254 ( .B(x[212]), .A(y[212]), .Z(n1153) );
  ANDN U255 ( .B(x[208]), .A(y[208]), .Z(n1141) );
  ANDN U256 ( .B(x[210]), .A(y[210]), .Z(n1147) );
  NOR U257 ( .A(n1141), .B(n1147), .Z(n154) );
  ANDN U258 ( .B(x[214]), .A(y[214]), .Z(n1159) );
  ANDN U259 ( .B(n154), .A(n1159), .Z(n155) );
  NANDN U260 ( .A(n1153), .B(n155), .Z(n156) );
  ANDN U261 ( .B(n157), .A(n156), .Z(n158) );
  NANDN U262 ( .A(n159), .B(n158), .Z(n160) );
  ANDN U263 ( .B(n161), .A(n160), .Z(n162) );
  NANDN U264 ( .A(n163), .B(n162), .Z(n323) );
  XNOR U265 ( .A(y[253]), .B(x[253]), .Z(n165) );
  NANDN U266 ( .A(x[252]), .B(y[252]), .Z(n164) );
  NAND U267 ( .A(n165), .B(n164), .Z(n1277) );
  XNOR U268 ( .A(y[249]), .B(x[249]), .Z(n167) );
  NANDN U269 ( .A(x[248]), .B(y[248]), .Z(n166) );
  NAND U270 ( .A(n167), .B(n166), .Z(n1265) );
  XNOR U271 ( .A(y[251]), .B(x[251]), .Z(n169) );
  NANDN U272 ( .A(x[250]), .B(y[250]), .Z(n168) );
  NAND U273 ( .A(n169), .B(n168), .Z(n1271) );
  NOR U274 ( .A(n1265), .B(n1271), .Z(n172) );
  XNOR U275 ( .A(y[255]), .B(x[255]), .Z(n171) );
  NANDN U276 ( .A(x[254]), .B(y[254]), .Z(n170) );
  NAND U277 ( .A(n171), .B(n170), .Z(n1283) );
  ANDN U278 ( .B(n172), .A(n1283), .Z(n173) );
  NANDN U279 ( .A(n1277), .B(n173), .Z(n209) );
  XNOR U280 ( .A(y[237]), .B(x[237]), .Z(n175) );
  NANDN U281 ( .A(x[236]), .B(y[236]), .Z(n174) );
  NAND U282 ( .A(n175), .B(n174), .Z(n1229) );
  XNOR U283 ( .A(y[233]), .B(x[233]), .Z(n177) );
  NANDN U284 ( .A(x[232]), .B(y[232]), .Z(n176) );
  NAND U285 ( .A(n177), .B(n176), .Z(n1217) );
  XNOR U286 ( .A(y[235]), .B(x[235]), .Z(n179) );
  NANDN U287 ( .A(x[234]), .B(y[234]), .Z(n178) );
  NAND U288 ( .A(n179), .B(n178), .Z(n1223) );
  NOR U289 ( .A(n1217), .B(n1223), .Z(n182) );
  XNOR U290 ( .A(y[239]), .B(x[239]), .Z(n181) );
  NANDN U291 ( .A(x[238]), .B(y[238]), .Z(n180) );
  NAND U292 ( .A(n181), .B(n180), .Z(n1235) );
  ANDN U293 ( .B(n182), .A(n1235), .Z(n183) );
  NANDN U294 ( .A(n1229), .B(n183), .Z(n195) );
  XNOR U295 ( .A(y[229]), .B(x[229]), .Z(n185) );
  NANDN U296 ( .A(x[228]), .B(y[228]), .Z(n184) );
  NAND U297 ( .A(n185), .B(n184), .Z(n1205) );
  XNOR U298 ( .A(y[225]), .B(x[225]), .Z(n187) );
  NANDN U299 ( .A(x[224]), .B(y[224]), .Z(n186) );
  NAND U300 ( .A(n187), .B(n186), .Z(n1193) );
  XNOR U301 ( .A(y[227]), .B(x[227]), .Z(n189) );
  NANDN U302 ( .A(x[226]), .B(y[226]), .Z(n188) );
  NAND U303 ( .A(n189), .B(n188), .Z(n1199) );
  NOR U304 ( .A(n1193), .B(n1199), .Z(n192) );
  XNOR U305 ( .A(y[231]), .B(x[231]), .Z(n191) );
  NANDN U306 ( .A(x[230]), .B(y[230]), .Z(n190) );
  NAND U307 ( .A(n191), .B(n190), .Z(n1211) );
  ANDN U308 ( .B(n192), .A(n1211), .Z(n193) );
  NANDN U309 ( .A(n1205), .B(n193), .Z(n194) );
  NOR U310 ( .A(n195), .B(n194), .Z(n207) );
  XNOR U311 ( .A(y[245]), .B(x[245]), .Z(n197) );
  NANDN U312 ( .A(x[244]), .B(y[244]), .Z(n196) );
  NAND U313 ( .A(n197), .B(n196), .Z(n1253) );
  XNOR U314 ( .A(y[241]), .B(x[241]), .Z(n199) );
  NANDN U315 ( .A(x[240]), .B(y[240]), .Z(n198) );
  NAND U316 ( .A(n199), .B(n198), .Z(n1241) );
  XNOR U317 ( .A(y[243]), .B(x[243]), .Z(n201) );
  NANDN U318 ( .A(x[242]), .B(y[242]), .Z(n200) );
  NAND U319 ( .A(n201), .B(n200), .Z(n1247) );
  NOR U320 ( .A(n1241), .B(n1247), .Z(n204) );
  XNOR U321 ( .A(y[247]), .B(x[247]), .Z(n203) );
  NANDN U322 ( .A(x[246]), .B(y[246]), .Z(n202) );
  NAND U323 ( .A(n203), .B(n202), .Z(n1259) );
  ANDN U324 ( .B(n204), .A(n1259), .Z(n205) );
  NANDN U325 ( .A(n1253), .B(n205), .Z(n206) );
  ANDN U326 ( .B(n207), .A(n206), .Z(n208) );
  NANDN U327 ( .A(n209), .B(n208), .Z(n257) );
  XNOR U328 ( .A(y[221]), .B(x[221]), .Z(n211) );
  NANDN U329 ( .A(x[220]), .B(y[220]), .Z(n210) );
  NAND U330 ( .A(n211), .B(n210), .Z(n1181) );
  XNOR U331 ( .A(y[217]), .B(x[217]), .Z(n213) );
  NANDN U332 ( .A(x[216]), .B(y[216]), .Z(n212) );
  NAND U333 ( .A(n213), .B(n212), .Z(n1169) );
  XNOR U334 ( .A(y[219]), .B(x[219]), .Z(n215) );
  NANDN U335 ( .A(x[218]), .B(y[218]), .Z(n214) );
  NAND U336 ( .A(n215), .B(n214), .Z(n1175) );
  NOR U337 ( .A(n1169), .B(n1175), .Z(n218) );
  XNOR U338 ( .A(y[223]), .B(x[223]), .Z(n217) );
  NANDN U339 ( .A(x[222]), .B(y[222]), .Z(n216) );
  NAND U340 ( .A(n217), .B(n216), .Z(n1187) );
  ANDN U341 ( .B(n218), .A(n1187), .Z(n219) );
  NANDN U342 ( .A(n1181), .B(n219), .Z(n255) );
  XNOR U343 ( .A(y[205]), .B(x[205]), .Z(n221) );
  NANDN U344 ( .A(x[204]), .B(y[204]), .Z(n220) );
  NAND U345 ( .A(n221), .B(n220), .Z(n1133) );
  XNOR U346 ( .A(y[201]), .B(x[201]), .Z(n223) );
  NANDN U347 ( .A(x[200]), .B(y[200]), .Z(n222) );
  NAND U348 ( .A(n223), .B(n222), .Z(n1121) );
  XNOR U349 ( .A(y[203]), .B(x[203]), .Z(n225) );
  NANDN U350 ( .A(x[202]), .B(y[202]), .Z(n224) );
  NAND U351 ( .A(n225), .B(n224), .Z(n1127) );
  NOR U352 ( .A(n1121), .B(n1127), .Z(n228) );
  XNOR U353 ( .A(y[207]), .B(x[207]), .Z(n227) );
  NANDN U354 ( .A(x[206]), .B(y[206]), .Z(n226) );
  NAND U355 ( .A(n227), .B(n226), .Z(n1139) );
  ANDN U356 ( .B(n228), .A(n1139), .Z(n229) );
  NANDN U357 ( .A(n1133), .B(n229), .Z(n241) );
  XNOR U358 ( .A(y[197]), .B(x[197]), .Z(n231) );
  NANDN U359 ( .A(x[196]), .B(y[196]), .Z(n230) );
  NAND U360 ( .A(n231), .B(n230), .Z(n1109) );
  XNOR U361 ( .A(y[193]), .B(x[193]), .Z(n233) );
  NANDN U362 ( .A(x[192]), .B(y[192]), .Z(n232) );
  NAND U363 ( .A(n233), .B(n232), .Z(n1097) );
  XNOR U364 ( .A(y[195]), .B(x[195]), .Z(n235) );
  NANDN U365 ( .A(x[194]), .B(y[194]), .Z(n234) );
  NAND U366 ( .A(n235), .B(n234), .Z(n1103) );
  NOR U367 ( .A(n1097), .B(n1103), .Z(n238) );
  XNOR U368 ( .A(y[199]), .B(x[199]), .Z(n237) );
  NANDN U369 ( .A(x[198]), .B(y[198]), .Z(n236) );
  NAND U370 ( .A(n237), .B(n236), .Z(n1115) );
  ANDN U371 ( .B(n238), .A(n1115), .Z(n239) );
  NANDN U372 ( .A(n1109), .B(n239), .Z(n240) );
  NOR U373 ( .A(n241), .B(n240), .Z(n253) );
  XNOR U374 ( .A(y[213]), .B(x[213]), .Z(n243) );
  NANDN U375 ( .A(x[212]), .B(y[212]), .Z(n242) );
  NAND U376 ( .A(n243), .B(n242), .Z(n1157) );
  XNOR U377 ( .A(y[209]), .B(x[209]), .Z(n245) );
  NANDN U378 ( .A(x[208]), .B(y[208]), .Z(n244) );
  NAND U379 ( .A(n245), .B(n244), .Z(n1145) );
  XNOR U380 ( .A(y[211]), .B(x[211]), .Z(n247) );
  NANDN U381 ( .A(x[210]), .B(y[210]), .Z(n246) );
  NAND U382 ( .A(n247), .B(n246), .Z(n1151) );
  NOR U383 ( .A(n1145), .B(n1151), .Z(n250) );
  XNOR U384 ( .A(y[215]), .B(x[215]), .Z(n249) );
  NANDN U385 ( .A(x[214]), .B(y[214]), .Z(n248) );
  NAND U386 ( .A(n249), .B(n248), .Z(n1163) );
  ANDN U387 ( .B(n250), .A(n1163), .Z(n251) );
  NANDN U388 ( .A(n1157), .B(n251), .Z(n252) );
  ANDN U389 ( .B(n253), .A(n252), .Z(n254) );
  NANDN U390 ( .A(n255), .B(n254), .Z(n256) );
  NOR U391 ( .A(n257), .B(n256), .Z(n321) );
  ANDN U392 ( .B(x[124]), .A(y[124]), .Z(n891) );
  ANDN U393 ( .B(x[120]), .A(y[120]), .Z(n879) );
  ANDN U394 ( .B(x[122]), .A(y[122]), .Z(n885) );
  NOR U395 ( .A(n879), .B(n885), .Z(n258) );
  ANDN U396 ( .B(x[126]), .A(y[126]), .Z(n897) );
  ANDN U397 ( .B(n258), .A(n897), .Z(n259) );
  NANDN U398 ( .A(n891), .B(n259), .Z(n271) );
  ANDN U399 ( .B(x[108]), .A(y[108]), .Z(n843) );
  ANDN U400 ( .B(x[104]), .A(y[104]), .Z(n831) );
  ANDN U401 ( .B(x[106]), .A(y[106]), .Z(n837) );
  NOR U402 ( .A(n831), .B(n837), .Z(n260) );
  ANDN U403 ( .B(x[110]), .A(y[110]), .Z(n849) );
  ANDN U404 ( .B(n260), .A(n849), .Z(n261) );
  NANDN U405 ( .A(n843), .B(n261), .Z(n265) );
  ANDN U406 ( .B(x[100]), .A(y[100]), .Z(n819) );
  ANDN U407 ( .B(x[96]), .A(y[96]), .Z(n807) );
  ANDN U408 ( .B(x[98]), .A(y[98]), .Z(n813) );
  NOR U409 ( .A(n807), .B(n813), .Z(n262) );
  ANDN U410 ( .B(x[102]), .A(y[102]), .Z(n825) );
  ANDN U411 ( .B(n262), .A(n825), .Z(n263) );
  NANDN U412 ( .A(n819), .B(n263), .Z(n264) );
  NOR U413 ( .A(n265), .B(n264), .Z(n269) );
  ANDN U414 ( .B(x[116]), .A(y[116]), .Z(n867) );
  ANDN U415 ( .B(x[112]), .A(y[112]), .Z(n855) );
  ANDN U416 ( .B(x[114]), .A(y[114]), .Z(n861) );
  NOR U417 ( .A(n855), .B(n861), .Z(n266) );
  ANDN U418 ( .B(x[118]), .A(y[118]), .Z(n873) );
  ANDN U419 ( .B(n266), .A(n873), .Z(n267) );
  NANDN U420 ( .A(n867), .B(n267), .Z(n268) );
  ANDN U421 ( .B(n269), .A(n268), .Z(n270) );
  NANDN U422 ( .A(n271), .B(n270), .Z(n319) );
  ANDN U423 ( .B(x[60]), .A(y[60]), .Z(n699) );
  ANDN U424 ( .B(x[56]), .A(y[56]), .Z(n687) );
  ANDN U425 ( .B(x[58]), .A(y[58]), .Z(n693) );
  NOR U426 ( .A(n687), .B(n693), .Z(n272) );
  ANDN U427 ( .B(x[62]), .A(y[62]), .Z(n705) );
  ANDN U428 ( .B(n272), .A(n705), .Z(n273) );
  NANDN U429 ( .A(n699), .B(n273), .Z(n285) );
  ANDN U430 ( .B(x[44]), .A(y[44]), .Z(n651) );
  ANDN U431 ( .B(x[40]), .A(y[40]), .Z(n639) );
  ANDN U432 ( .B(x[42]), .A(y[42]), .Z(n645) );
  NOR U433 ( .A(n639), .B(n645), .Z(n274) );
  ANDN U434 ( .B(x[46]), .A(y[46]), .Z(n657) );
  ANDN U435 ( .B(n274), .A(n657), .Z(n275) );
  NANDN U436 ( .A(n651), .B(n275), .Z(n279) );
  ANDN U437 ( .B(x[36]), .A(y[36]), .Z(n627) );
  ANDN U438 ( .B(x[32]), .A(y[32]), .Z(n615) );
  ANDN U439 ( .B(x[34]), .A(y[34]), .Z(n621) );
  NOR U440 ( .A(n615), .B(n621), .Z(n276) );
  ANDN U441 ( .B(x[38]), .A(y[38]), .Z(n633) );
  ANDN U442 ( .B(n276), .A(n633), .Z(n277) );
  NANDN U443 ( .A(n627), .B(n277), .Z(n278) );
  NOR U444 ( .A(n279), .B(n278), .Z(n283) );
  ANDN U445 ( .B(x[52]), .A(y[52]), .Z(n675) );
  ANDN U446 ( .B(x[48]), .A(y[48]), .Z(n663) );
  ANDN U447 ( .B(x[50]), .A(y[50]), .Z(n669) );
  NOR U448 ( .A(n663), .B(n669), .Z(n280) );
  ANDN U449 ( .B(x[54]), .A(y[54]), .Z(n681) );
  ANDN U450 ( .B(n280), .A(n681), .Z(n281) );
  NANDN U451 ( .A(n675), .B(n281), .Z(n282) );
  ANDN U452 ( .B(n283), .A(n282), .Z(n284) );
  NANDN U453 ( .A(n285), .B(n284), .Z(n301) );
  ANDN U454 ( .B(x[28]), .A(y[28]), .Z(n603) );
  ANDN U455 ( .B(x[24]), .A(y[24]), .Z(n591) );
  ANDN U456 ( .B(x[26]), .A(y[26]), .Z(n597) );
  NOR U457 ( .A(n591), .B(n597), .Z(n286) );
  ANDN U458 ( .B(x[30]), .A(y[30]), .Z(n609) );
  ANDN U459 ( .B(n286), .A(n609), .Z(n287) );
  NANDN U460 ( .A(n603), .B(n287), .Z(n299) );
  NANDN U461 ( .A(y[8]), .B(x[8]), .Z(n525) );
  ANDN U462 ( .B(x[10]), .A(y[10]), .Z(n522) );
  ANDN U463 ( .B(n525), .A(n522), .Z(n288) );
  ANDN U464 ( .B(x[14]), .A(y[14]), .Z(n561) );
  ANDN U465 ( .B(n288), .A(n561), .Z(n289) );
  NANDN U466 ( .A(y[12]), .B(x[12]), .Z(n521) );
  NAND U467 ( .A(n289), .B(n521), .Z(n293) );
  NANDN U468 ( .A(y[6]), .B(x[6]), .Z(n527) );
  NANDN U469 ( .A(y[0]), .B(x[0]), .Z(n530) );
  NANDN U470 ( .A(y[4]), .B(x[4]), .Z(n529) );
  AND U471 ( .A(n530), .B(n529), .Z(n290) );
  AND U472 ( .A(n527), .B(n290), .Z(n291) );
  NANDN U473 ( .A(y[2]), .B(x[2]), .Z(n535) );
  NAND U474 ( .A(n291), .B(n535), .Z(n292) );
  NOR U475 ( .A(n293), .B(n292), .Z(n297) );
  ANDN U476 ( .B(x[20]), .A(y[20]), .Z(n579) );
  ANDN U477 ( .B(x[16]), .A(y[16]), .Z(n567) );
  ANDN U478 ( .B(x[18]), .A(y[18]), .Z(n573) );
  NOR U479 ( .A(n567), .B(n573), .Z(n294) );
  ANDN U480 ( .B(x[22]), .A(y[22]), .Z(n585) );
  ANDN U481 ( .B(n294), .A(n585), .Z(n295) );
  NANDN U482 ( .A(n579), .B(n295), .Z(n296) );
  ANDN U483 ( .B(n297), .A(n296), .Z(n298) );
  NANDN U484 ( .A(n299), .B(n298), .Z(n300) );
  NOR U485 ( .A(n301), .B(n300), .Z(n317) );
  ANDN U486 ( .B(x[92]), .A(y[92]), .Z(n795) );
  ANDN U487 ( .B(x[88]), .A(y[88]), .Z(n783) );
  ANDN U488 ( .B(x[90]), .A(y[90]), .Z(n789) );
  NOR U489 ( .A(n783), .B(n789), .Z(n302) );
  ANDN U490 ( .B(x[94]), .A(y[94]), .Z(n801) );
  ANDN U491 ( .B(n302), .A(n801), .Z(n303) );
  NANDN U492 ( .A(n795), .B(n303), .Z(n315) );
  ANDN U493 ( .B(x[76]), .A(y[76]), .Z(n747) );
  ANDN U494 ( .B(x[72]), .A(y[72]), .Z(n735) );
  ANDN U495 ( .B(x[74]), .A(y[74]), .Z(n741) );
  NOR U496 ( .A(n735), .B(n741), .Z(n304) );
  ANDN U497 ( .B(x[78]), .A(y[78]), .Z(n753) );
  ANDN U498 ( .B(n304), .A(n753), .Z(n305) );
  NANDN U499 ( .A(n747), .B(n305), .Z(n309) );
  ANDN U500 ( .B(x[68]), .A(y[68]), .Z(n723) );
  ANDN U501 ( .B(x[64]), .A(y[64]), .Z(n711) );
  ANDN U502 ( .B(x[66]), .A(y[66]), .Z(n717) );
  NOR U503 ( .A(n711), .B(n717), .Z(n306) );
  ANDN U504 ( .B(x[70]), .A(y[70]), .Z(n729) );
  ANDN U505 ( .B(n306), .A(n729), .Z(n307) );
  NANDN U506 ( .A(n723), .B(n307), .Z(n308) );
  NOR U507 ( .A(n309), .B(n308), .Z(n313) );
  ANDN U508 ( .B(x[84]), .A(y[84]), .Z(n771) );
  ANDN U509 ( .B(x[80]), .A(y[80]), .Z(n759) );
  ANDN U510 ( .B(x[82]), .A(y[82]), .Z(n765) );
  NOR U511 ( .A(n759), .B(n765), .Z(n310) );
  ANDN U512 ( .B(x[86]), .A(y[86]), .Z(n777) );
  ANDN U513 ( .B(n310), .A(n777), .Z(n311) );
  NANDN U514 ( .A(n771), .B(n311), .Z(n312) );
  ANDN U515 ( .B(n313), .A(n312), .Z(n314) );
  NANDN U516 ( .A(n315), .B(n314), .Z(n316) );
  ANDN U517 ( .B(n317), .A(n316), .Z(n318) );
  NANDN U518 ( .A(n319), .B(n318), .Z(n320) );
  ANDN U519 ( .B(n321), .A(n320), .Z(n322) );
  NANDN U520 ( .A(n323), .B(n322), .Z(n324) );
  ANDN U521 ( .B(n325), .A(n324), .Z(n518) );
  XNOR U522 ( .A(y[85]), .B(x[85]), .Z(n327) );
  NANDN U523 ( .A(x[84]), .B(y[84]), .Z(n326) );
  NAND U524 ( .A(n327), .B(n326), .Z(n773) );
  XNOR U525 ( .A(y[81]), .B(x[81]), .Z(n329) );
  NANDN U526 ( .A(x[80]), .B(y[80]), .Z(n328) );
  NAND U527 ( .A(n329), .B(n328), .Z(n761) );
  XNOR U528 ( .A(y[83]), .B(x[83]), .Z(n331) );
  NANDN U529 ( .A(x[82]), .B(y[82]), .Z(n330) );
  NAND U530 ( .A(n331), .B(n330), .Z(n767) );
  NOR U531 ( .A(n761), .B(n767), .Z(n334) );
  XNOR U532 ( .A(y[87]), .B(x[87]), .Z(n333) );
  NANDN U533 ( .A(x[86]), .B(y[86]), .Z(n332) );
  NAND U534 ( .A(n333), .B(n332), .Z(n779) );
  ANDN U535 ( .B(n334), .A(n779), .Z(n335) );
  NANDN U536 ( .A(n773), .B(n335), .Z(n371) );
  XNOR U537 ( .A(y[69]), .B(x[69]), .Z(n337) );
  NANDN U538 ( .A(x[68]), .B(y[68]), .Z(n336) );
  NAND U539 ( .A(n337), .B(n336), .Z(n725) );
  XNOR U540 ( .A(y[65]), .B(x[65]), .Z(n339) );
  NANDN U541 ( .A(x[64]), .B(y[64]), .Z(n338) );
  NAND U542 ( .A(n339), .B(n338), .Z(n713) );
  XNOR U543 ( .A(y[67]), .B(x[67]), .Z(n341) );
  NANDN U544 ( .A(x[66]), .B(y[66]), .Z(n340) );
  NAND U545 ( .A(n341), .B(n340), .Z(n719) );
  NOR U546 ( .A(n713), .B(n719), .Z(n344) );
  XNOR U547 ( .A(y[71]), .B(x[71]), .Z(n343) );
  NANDN U548 ( .A(x[70]), .B(y[70]), .Z(n342) );
  NAND U549 ( .A(n343), .B(n342), .Z(n731) );
  ANDN U550 ( .B(n344), .A(n731), .Z(n345) );
  NANDN U551 ( .A(n725), .B(n345), .Z(n357) );
  XNOR U552 ( .A(y[77]), .B(x[77]), .Z(n347) );
  NANDN U553 ( .A(x[76]), .B(y[76]), .Z(n346) );
  NAND U554 ( .A(n347), .B(n346), .Z(n749) );
  XNOR U555 ( .A(y[73]), .B(x[73]), .Z(n349) );
  NANDN U556 ( .A(x[72]), .B(y[72]), .Z(n348) );
  NAND U557 ( .A(n349), .B(n348), .Z(n737) );
  XNOR U558 ( .A(y[75]), .B(x[75]), .Z(n351) );
  NANDN U559 ( .A(x[74]), .B(y[74]), .Z(n350) );
  NAND U560 ( .A(n351), .B(n350), .Z(n743) );
  NOR U561 ( .A(n737), .B(n743), .Z(n354) );
  XNOR U562 ( .A(y[79]), .B(x[79]), .Z(n353) );
  NANDN U563 ( .A(x[78]), .B(y[78]), .Z(n352) );
  NAND U564 ( .A(n353), .B(n352), .Z(n755) );
  ANDN U565 ( .B(n354), .A(n755), .Z(n355) );
  NANDN U566 ( .A(n749), .B(n355), .Z(n356) );
  NOR U567 ( .A(n357), .B(n356), .Z(n369) );
  XNOR U568 ( .A(y[93]), .B(x[93]), .Z(n359) );
  NANDN U569 ( .A(x[92]), .B(y[92]), .Z(n358) );
  NAND U570 ( .A(n359), .B(n358), .Z(n797) );
  XNOR U571 ( .A(y[89]), .B(x[89]), .Z(n361) );
  NANDN U572 ( .A(x[88]), .B(y[88]), .Z(n360) );
  NAND U573 ( .A(n361), .B(n360), .Z(n785) );
  XNOR U574 ( .A(y[91]), .B(x[91]), .Z(n363) );
  NANDN U575 ( .A(x[90]), .B(y[90]), .Z(n362) );
  NAND U576 ( .A(n363), .B(n362), .Z(n791) );
  NOR U577 ( .A(n785), .B(n791), .Z(n366) );
  XNOR U578 ( .A(y[95]), .B(x[95]), .Z(n365) );
  NANDN U579 ( .A(x[94]), .B(y[94]), .Z(n364) );
  NAND U580 ( .A(n365), .B(n364), .Z(n803) );
  ANDN U581 ( .B(n366), .A(n803), .Z(n367) );
  NANDN U582 ( .A(n797), .B(n367), .Z(n368) );
  ANDN U583 ( .B(n369), .A(n368), .Z(n370) );
  NANDN U584 ( .A(n371), .B(n370), .Z(n516) );
  XNOR U585 ( .A(y[21]), .B(x[21]), .Z(n373) );
  NANDN U586 ( .A(x[20]), .B(y[20]), .Z(n372) );
  NAND U587 ( .A(n373), .B(n372), .Z(n581) );
  XNOR U588 ( .A(y[17]), .B(x[17]), .Z(n375) );
  NANDN U589 ( .A(x[16]), .B(y[16]), .Z(n374) );
  NAND U590 ( .A(n375), .B(n374), .Z(n569) );
  XNOR U591 ( .A(y[19]), .B(x[19]), .Z(n377) );
  NANDN U592 ( .A(x[18]), .B(y[18]), .Z(n376) );
  NAND U593 ( .A(n377), .B(n376), .Z(n575) );
  NOR U594 ( .A(n569), .B(n575), .Z(n380) );
  XNOR U595 ( .A(y[23]), .B(x[23]), .Z(n379) );
  NANDN U596 ( .A(x[22]), .B(y[22]), .Z(n378) );
  NAND U597 ( .A(n379), .B(n378), .Z(n587) );
  ANDN U598 ( .B(n380), .A(n587), .Z(n381) );
  NANDN U599 ( .A(n581), .B(n381), .Z(n418) );
  XNOR U600 ( .A(y[7]), .B(x[7]), .Z(n383) );
  NANDN U601 ( .A(x[6]), .B(y[6]), .Z(n382) );
  NAND U602 ( .A(n383), .B(n382), .Z(n545) );
  XNOR U603 ( .A(y[3]), .B(x[3]), .Z(n385) );
  NANDN U604 ( .A(x[2]), .B(y[2]), .Z(n384) );
  NAND U605 ( .A(n385), .B(n384), .Z(n537) );
  XNOR U606 ( .A(y[5]), .B(x[5]), .Z(n387) );
  NANDN U607 ( .A(x[4]), .B(y[4]), .Z(n386) );
  NAND U608 ( .A(n387), .B(n386), .Z(n541) );
  NOR U609 ( .A(n537), .B(n541), .Z(n391) );
  XNOR U610 ( .A(y[1]), .B(x[1]), .Z(n389) );
  NANDN U611 ( .A(x[0]), .B(y[0]), .Z(n388) );
  NAND U612 ( .A(n389), .B(n388), .Z(n390) );
  ANDN U613 ( .B(n391), .A(n390), .Z(n392) );
  NANDN U614 ( .A(n545), .B(n392), .Z(n404) );
  XNOR U615 ( .A(y[13]), .B(x[13]), .Z(n394) );
  NANDN U616 ( .A(x[12]), .B(y[12]), .Z(n393) );
  NAND U617 ( .A(n394), .B(n393), .Z(n557) );
  XNOR U618 ( .A(y[9]), .B(x[9]), .Z(n396) );
  NANDN U619 ( .A(x[8]), .B(y[8]), .Z(n395) );
  NAND U620 ( .A(n396), .B(n395), .Z(n549) );
  XNOR U621 ( .A(y[11]), .B(x[11]), .Z(n398) );
  NANDN U622 ( .A(x[10]), .B(y[10]), .Z(n397) );
  NAND U623 ( .A(n398), .B(n397), .Z(n553) );
  NOR U624 ( .A(n549), .B(n553), .Z(n401) );
  XNOR U625 ( .A(y[15]), .B(x[15]), .Z(n400) );
  NANDN U626 ( .A(x[14]), .B(y[14]), .Z(n399) );
  NAND U627 ( .A(n400), .B(n399), .Z(n563) );
  ANDN U628 ( .B(n401), .A(n563), .Z(n402) );
  NANDN U629 ( .A(n557), .B(n402), .Z(n403) );
  NOR U630 ( .A(n404), .B(n403), .Z(n416) );
  XNOR U631 ( .A(y[29]), .B(x[29]), .Z(n406) );
  NANDN U632 ( .A(x[28]), .B(y[28]), .Z(n405) );
  NAND U633 ( .A(n406), .B(n405), .Z(n605) );
  XNOR U634 ( .A(y[25]), .B(x[25]), .Z(n408) );
  NANDN U635 ( .A(x[24]), .B(y[24]), .Z(n407) );
  NAND U636 ( .A(n408), .B(n407), .Z(n593) );
  XNOR U637 ( .A(y[27]), .B(x[27]), .Z(n410) );
  NANDN U638 ( .A(x[26]), .B(y[26]), .Z(n409) );
  NAND U639 ( .A(n410), .B(n409), .Z(n599) );
  NOR U640 ( .A(n593), .B(n599), .Z(n413) );
  XNOR U641 ( .A(y[31]), .B(x[31]), .Z(n412) );
  NANDN U642 ( .A(x[30]), .B(y[30]), .Z(n411) );
  NAND U643 ( .A(n412), .B(n411), .Z(n611) );
  ANDN U644 ( .B(n413), .A(n611), .Z(n414) );
  NANDN U645 ( .A(n605), .B(n414), .Z(n415) );
  ANDN U646 ( .B(n416), .A(n415), .Z(n417) );
  NANDN U647 ( .A(n418), .B(n417), .Z(n466) );
  XNOR U648 ( .A(y[53]), .B(x[53]), .Z(n420) );
  NANDN U649 ( .A(x[52]), .B(y[52]), .Z(n419) );
  NAND U650 ( .A(n420), .B(n419), .Z(n677) );
  XNOR U651 ( .A(y[49]), .B(x[49]), .Z(n422) );
  NANDN U652 ( .A(x[48]), .B(y[48]), .Z(n421) );
  NAND U653 ( .A(n422), .B(n421), .Z(n665) );
  XNOR U654 ( .A(y[51]), .B(x[51]), .Z(n424) );
  NANDN U655 ( .A(x[50]), .B(y[50]), .Z(n423) );
  NAND U656 ( .A(n424), .B(n423), .Z(n671) );
  NOR U657 ( .A(n665), .B(n671), .Z(n427) );
  XNOR U658 ( .A(y[55]), .B(x[55]), .Z(n426) );
  NANDN U659 ( .A(x[54]), .B(y[54]), .Z(n425) );
  NAND U660 ( .A(n426), .B(n425), .Z(n683) );
  ANDN U661 ( .B(n427), .A(n683), .Z(n428) );
  NANDN U662 ( .A(n677), .B(n428), .Z(n464) );
  XNOR U663 ( .A(y[37]), .B(x[37]), .Z(n430) );
  NANDN U664 ( .A(x[36]), .B(y[36]), .Z(n429) );
  NAND U665 ( .A(n430), .B(n429), .Z(n629) );
  XNOR U666 ( .A(y[33]), .B(x[33]), .Z(n432) );
  NANDN U667 ( .A(x[32]), .B(y[32]), .Z(n431) );
  NAND U668 ( .A(n432), .B(n431), .Z(n617) );
  XNOR U669 ( .A(y[35]), .B(x[35]), .Z(n434) );
  NANDN U670 ( .A(x[34]), .B(y[34]), .Z(n433) );
  NAND U671 ( .A(n434), .B(n433), .Z(n623) );
  NOR U672 ( .A(n617), .B(n623), .Z(n437) );
  XNOR U673 ( .A(y[39]), .B(x[39]), .Z(n436) );
  NANDN U674 ( .A(x[38]), .B(y[38]), .Z(n435) );
  NAND U675 ( .A(n436), .B(n435), .Z(n635) );
  ANDN U676 ( .B(n437), .A(n635), .Z(n438) );
  NANDN U677 ( .A(n629), .B(n438), .Z(n450) );
  XNOR U678 ( .A(y[45]), .B(x[45]), .Z(n440) );
  NANDN U679 ( .A(x[44]), .B(y[44]), .Z(n439) );
  NAND U680 ( .A(n440), .B(n439), .Z(n653) );
  XNOR U681 ( .A(y[41]), .B(x[41]), .Z(n442) );
  NANDN U682 ( .A(x[40]), .B(y[40]), .Z(n441) );
  NAND U683 ( .A(n442), .B(n441), .Z(n641) );
  XNOR U684 ( .A(y[43]), .B(x[43]), .Z(n444) );
  NANDN U685 ( .A(x[42]), .B(y[42]), .Z(n443) );
  NAND U686 ( .A(n444), .B(n443), .Z(n647) );
  NOR U687 ( .A(n641), .B(n647), .Z(n447) );
  XNOR U688 ( .A(y[47]), .B(x[47]), .Z(n446) );
  NANDN U689 ( .A(x[46]), .B(y[46]), .Z(n445) );
  NAND U690 ( .A(n446), .B(n445), .Z(n659) );
  ANDN U691 ( .B(n447), .A(n659), .Z(n448) );
  NANDN U692 ( .A(n653), .B(n448), .Z(n449) );
  NOR U693 ( .A(n450), .B(n449), .Z(n462) );
  XNOR U694 ( .A(y[61]), .B(x[61]), .Z(n452) );
  NANDN U695 ( .A(x[60]), .B(y[60]), .Z(n451) );
  NAND U696 ( .A(n452), .B(n451), .Z(n701) );
  XNOR U697 ( .A(y[57]), .B(x[57]), .Z(n454) );
  NANDN U698 ( .A(x[56]), .B(y[56]), .Z(n453) );
  NAND U699 ( .A(n454), .B(n453), .Z(n689) );
  XNOR U700 ( .A(y[59]), .B(x[59]), .Z(n456) );
  NANDN U701 ( .A(x[58]), .B(y[58]), .Z(n455) );
  NAND U702 ( .A(n456), .B(n455), .Z(n695) );
  NOR U703 ( .A(n689), .B(n695), .Z(n459) );
  XNOR U704 ( .A(y[63]), .B(x[63]), .Z(n458) );
  NANDN U705 ( .A(x[62]), .B(y[62]), .Z(n457) );
  NAND U706 ( .A(n458), .B(n457), .Z(n707) );
  ANDN U707 ( .B(n459), .A(n707), .Z(n460) );
  NANDN U708 ( .A(n701), .B(n460), .Z(n461) );
  ANDN U709 ( .B(n462), .A(n461), .Z(n463) );
  NANDN U710 ( .A(n464), .B(n463), .Z(n465) );
  NOR U711 ( .A(n466), .B(n465), .Z(n514) );
  XNOR U712 ( .A(y[117]), .B(x[117]), .Z(n468) );
  NANDN U713 ( .A(x[116]), .B(y[116]), .Z(n467) );
  NAND U714 ( .A(n468), .B(n467), .Z(n869) );
  XNOR U715 ( .A(y[113]), .B(x[113]), .Z(n470) );
  NANDN U716 ( .A(x[112]), .B(y[112]), .Z(n469) );
  NAND U717 ( .A(n470), .B(n469), .Z(n857) );
  XNOR U718 ( .A(y[115]), .B(x[115]), .Z(n472) );
  NANDN U719 ( .A(x[114]), .B(y[114]), .Z(n471) );
  NAND U720 ( .A(n472), .B(n471), .Z(n863) );
  NOR U721 ( .A(n857), .B(n863), .Z(n475) );
  XNOR U722 ( .A(y[119]), .B(x[119]), .Z(n474) );
  NANDN U723 ( .A(x[118]), .B(y[118]), .Z(n473) );
  NAND U724 ( .A(n474), .B(n473), .Z(n875) );
  ANDN U725 ( .B(n475), .A(n875), .Z(n476) );
  NANDN U726 ( .A(n869), .B(n476), .Z(n512) );
  XNOR U727 ( .A(y[101]), .B(x[101]), .Z(n478) );
  NANDN U728 ( .A(x[100]), .B(y[100]), .Z(n477) );
  NAND U729 ( .A(n478), .B(n477), .Z(n821) );
  XNOR U730 ( .A(y[97]), .B(x[97]), .Z(n480) );
  NANDN U731 ( .A(x[96]), .B(y[96]), .Z(n479) );
  NAND U732 ( .A(n480), .B(n479), .Z(n809) );
  XNOR U733 ( .A(y[99]), .B(x[99]), .Z(n482) );
  NANDN U734 ( .A(x[98]), .B(y[98]), .Z(n481) );
  NAND U735 ( .A(n482), .B(n481), .Z(n815) );
  NOR U736 ( .A(n809), .B(n815), .Z(n485) );
  XNOR U737 ( .A(y[103]), .B(x[103]), .Z(n484) );
  NANDN U738 ( .A(x[102]), .B(y[102]), .Z(n483) );
  NAND U739 ( .A(n484), .B(n483), .Z(n827) );
  ANDN U740 ( .B(n485), .A(n827), .Z(n486) );
  NANDN U741 ( .A(n821), .B(n486), .Z(n498) );
  XNOR U742 ( .A(y[109]), .B(x[109]), .Z(n488) );
  NANDN U743 ( .A(x[108]), .B(y[108]), .Z(n487) );
  NAND U744 ( .A(n488), .B(n487), .Z(n845) );
  XNOR U745 ( .A(y[105]), .B(x[105]), .Z(n490) );
  NANDN U746 ( .A(x[104]), .B(y[104]), .Z(n489) );
  NAND U747 ( .A(n490), .B(n489), .Z(n833) );
  XNOR U748 ( .A(y[107]), .B(x[107]), .Z(n492) );
  NANDN U749 ( .A(x[106]), .B(y[106]), .Z(n491) );
  NAND U750 ( .A(n492), .B(n491), .Z(n839) );
  NOR U751 ( .A(n833), .B(n839), .Z(n495) );
  XNOR U752 ( .A(y[111]), .B(x[111]), .Z(n494) );
  NANDN U753 ( .A(x[110]), .B(y[110]), .Z(n493) );
  NAND U754 ( .A(n494), .B(n493), .Z(n851) );
  ANDN U755 ( .B(n495), .A(n851), .Z(n496) );
  NANDN U756 ( .A(n845), .B(n496), .Z(n497) );
  NOR U757 ( .A(n498), .B(n497), .Z(n510) );
  XNOR U758 ( .A(y[125]), .B(x[125]), .Z(n500) );
  NANDN U759 ( .A(x[124]), .B(y[124]), .Z(n499) );
  NAND U760 ( .A(n500), .B(n499), .Z(n893) );
  XNOR U761 ( .A(y[121]), .B(x[121]), .Z(n502) );
  NANDN U762 ( .A(x[120]), .B(y[120]), .Z(n501) );
  NAND U763 ( .A(n502), .B(n501), .Z(n881) );
  XNOR U764 ( .A(y[123]), .B(x[123]), .Z(n504) );
  NANDN U765 ( .A(x[122]), .B(y[122]), .Z(n503) );
  NAND U766 ( .A(n504), .B(n503), .Z(n887) );
  NOR U767 ( .A(n881), .B(n887), .Z(n507) );
  XNOR U768 ( .A(y[127]), .B(x[127]), .Z(n506) );
  NANDN U769 ( .A(x[126]), .B(y[126]), .Z(n505) );
  NAND U770 ( .A(n506), .B(n505), .Z(n899) );
  ANDN U771 ( .B(n507), .A(n899), .Z(n508) );
  NANDN U772 ( .A(n893), .B(n508), .Z(n509) );
  ANDN U773 ( .B(n510), .A(n509), .Z(n511) );
  NANDN U774 ( .A(n512), .B(n511), .Z(n513) );
  ANDN U775 ( .B(n514), .A(n513), .Z(n515) );
  NANDN U776 ( .A(n516), .B(n515), .Z(n517) );
  ANDN U777 ( .B(n518), .A(n517), .Z(n519) );
  NAND U778 ( .A(e), .B(n519), .Z(n5) );
  NANDN U779 ( .A(n519), .B(e), .Z(n1287) );
  ANDN U780 ( .B(x[255]), .A(y[255]), .Z(n1285) );
  ANDN U781 ( .B(x[127]), .A(y[127]), .Z(n901) );
  ANDN U782 ( .B(x[125]), .A(y[125]), .Z(n895) );
  ANDN U783 ( .B(x[123]), .A(y[123]), .Z(n889) );
  ANDN U784 ( .B(x[121]), .A(y[121]), .Z(n883) );
  ANDN U785 ( .B(x[119]), .A(y[119]), .Z(n877) );
  ANDN U786 ( .B(x[117]), .A(y[117]), .Z(n871) );
  ANDN U787 ( .B(x[115]), .A(y[115]), .Z(n865) );
  ANDN U788 ( .B(x[113]), .A(y[113]), .Z(n859) );
  ANDN U789 ( .B(x[111]), .A(y[111]), .Z(n853) );
  ANDN U790 ( .B(x[109]), .A(y[109]), .Z(n847) );
  ANDN U791 ( .B(x[107]), .A(y[107]), .Z(n841) );
  ANDN U792 ( .B(x[105]), .A(y[105]), .Z(n835) );
  ANDN U793 ( .B(x[103]), .A(y[103]), .Z(n829) );
  ANDN U794 ( .B(x[101]), .A(y[101]), .Z(n823) );
  ANDN U795 ( .B(x[99]), .A(y[99]), .Z(n817) );
  ANDN U796 ( .B(x[97]), .A(y[97]), .Z(n811) );
  ANDN U797 ( .B(x[95]), .A(y[95]), .Z(n805) );
  ANDN U798 ( .B(x[93]), .A(y[93]), .Z(n799) );
  ANDN U799 ( .B(x[91]), .A(y[91]), .Z(n793) );
  ANDN U800 ( .B(x[89]), .A(y[89]), .Z(n787) );
  ANDN U801 ( .B(x[87]), .A(y[87]), .Z(n781) );
  ANDN U802 ( .B(x[85]), .A(y[85]), .Z(n775) );
  ANDN U803 ( .B(x[83]), .A(y[83]), .Z(n769) );
  ANDN U804 ( .B(x[81]), .A(y[81]), .Z(n763) );
  ANDN U805 ( .B(x[79]), .A(y[79]), .Z(n757) );
  ANDN U806 ( .B(x[77]), .A(y[77]), .Z(n751) );
  ANDN U807 ( .B(x[75]), .A(y[75]), .Z(n745) );
  ANDN U808 ( .B(x[73]), .A(y[73]), .Z(n739) );
  ANDN U809 ( .B(x[71]), .A(y[71]), .Z(n733) );
  ANDN U810 ( .B(x[69]), .A(y[69]), .Z(n727) );
  ANDN U811 ( .B(x[67]), .A(y[67]), .Z(n721) );
  ANDN U812 ( .B(x[65]), .A(y[65]), .Z(n715) );
  ANDN U813 ( .B(x[63]), .A(y[63]), .Z(n709) );
  ANDN U814 ( .B(x[61]), .A(y[61]), .Z(n703) );
  ANDN U815 ( .B(x[59]), .A(y[59]), .Z(n697) );
  ANDN U816 ( .B(x[57]), .A(y[57]), .Z(n691) );
  ANDN U817 ( .B(x[55]), .A(y[55]), .Z(n685) );
  ANDN U818 ( .B(x[53]), .A(y[53]), .Z(n679) );
  ANDN U819 ( .B(x[51]), .A(y[51]), .Z(n673) );
  ANDN U820 ( .B(x[49]), .A(y[49]), .Z(n667) );
  ANDN U821 ( .B(x[47]), .A(y[47]), .Z(n661) );
  ANDN U822 ( .B(x[45]), .A(y[45]), .Z(n655) );
  ANDN U823 ( .B(x[43]), .A(y[43]), .Z(n649) );
  ANDN U824 ( .B(x[41]), .A(y[41]), .Z(n643) );
  ANDN U825 ( .B(x[39]), .A(y[39]), .Z(n637) );
  ANDN U826 ( .B(x[37]), .A(y[37]), .Z(n631) );
  ANDN U827 ( .B(x[35]), .A(y[35]), .Z(n625) );
  ANDN U828 ( .B(x[33]), .A(y[33]), .Z(n619) );
  ANDN U829 ( .B(x[31]), .A(y[31]), .Z(n613) );
  ANDN U830 ( .B(x[29]), .A(y[29]), .Z(n607) );
  ANDN U831 ( .B(x[27]), .A(y[27]), .Z(n601) );
  ANDN U832 ( .B(x[25]), .A(y[25]), .Z(n595) );
  ANDN U833 ( .B(x[23]), .A(y[23]), .Z(n589) );
  ANDN U834 ( .B(x[21]), .A(y[21]), .Z(n583) );
  ANDN U835 ( .B(x[19]), .A(y[19]), .Z(n577) );
  ANDN U836 ( .B(x[17]), .A(y[17]), .Z(n571) );
  ANDN U837 ( .B(x[15]), .A(y[15]), .Z(n565) );
  NANDN U838 ( .A(y[13]), .B(x[13]), .Z(n559) );
  NANDN U839 ( .A(y[11]), .B(x[11]), .Z(n520) );
  AND U840 ( .A(n521), .B(n520), .Z(n555) );
  NANDN U841 ( .A(y[9]), .B(x[9]), .Z(n523) );
  ANDN U842 ( .B(n523), .A(n522), .Z(n551) );
  NANDN U843 ( .A(y[7]), .B(x[7]), .Z(n524) );
  AND U844 ( .A(n525), .B(n524), .Z(n547) );
  NANDN U845 ( .A(y[5]), .B(x[5]), .Z(n526) );
  AND U846 ( .A(n527), .B(n526), .Z(n543) );
  NANDN U847 ( .A(y[3]), .B(x[3]), .Z(n528) );
  AND U848 ( .A(n529), .B(n528), .Z(n539) );
  NANDN U849 ( .A(x[1]), .B(n530), .Z(n533) );
  XNOR U850 ( .A(n530), .B(x[1]), .Z(n531) );
  NAND U851 ( .A(n531), .B(y[1]), .Z(n532) );
  NAND U852 ( .A(n533), .B(n532), .Z(n534) );
  AND U853 ( .A(n535), .B(n534), .Z(n536) );
  OR U854 ( .A(n537), .B(n536), .Z(n538) );
  AND U855 ( .A(n539), .B(n538), .Z(n540) );
  OR U856 ( .A(n541), .B(n540), .Z(n542) );
  AND U857 ( .A(n543), .B(n542), .Z(n544) );
  OR U858 ( .A(n545), .B(n544), .Z(n546) );
  AND U859 ( .A(n547), .B(n546), .Z(n548) );
  OR U860 ( .A(n549), .B(n548), .Z(n550) );
  AND U861 ( .A(n551), .B(n550), .Z(n552) );
  OR U862 ( .A(n553), .B(n552), .Z(n554) );
  AND U863 ( .A(n555), .B(n554), .Z(n556) );
  OR U864 ( .A(n557), .B(n556), .Z(n558) );
  AND U865 ( .A(n559), .B(n558), .Z(n560) );
  NANDN U866 ( .A(n561), .B(n560), .Z(n562) );
  NANDN U867 ( .A(n563), .B(n562), .Z(n564) );
  NANDN U868 ( .A(n565), .B(n564), .Z(n566) );
  OR U869 ( .A(n567), .B(n566), .Z(n568) );
  NANDN U870 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U871 ( .A(n571), .B(n570), .Z(n572) );
  OR U872 ( .A(n573), .B(n572), .Z(n574) );
  NANDN U873 ( .A(n575), .B(n574), .Z(n576) );
  NANDN U874 ( .A(n577), .B(n576), .Z(n578) );
  OR U875 ( .A(n579), .B(n578), .Z(n580) );
  NANDN U876 ( .A(n581), .B(n580), .Z(n582) );
  NANDN U877 ( .A(n583), .B(n582), .Z(n584) );
  OR U878 ( .A(n585), .B(n584), .Z(n586) );
  NANDN U879 ( .A(n587), .B(n586), .Z(n588) );
  NANDN U880 ( .A(n589), .B(n588), .Z(n590) );
  OR U881 ( .A(n591), .B(n590), .Z(n592) );
  NANDN U882 ( .A(n593), .B(n592), .Z(n594) );
  NANDN U883 ( .A(n595), .B(n594), .Z(n596) );
  OR U884 ( .A(n597), .B(n596), .Z(n598) );
  NANDN U885 ( .A(n599), .B(n598), .Z(n600) );
  NANDN U886 ( .A(n601), .B(n600), .Z(n602) );
  OR U887 ( .A(n603), .B(n602), .Z(n604) );
  NANDN U888 ( .A(n605), .B(n604), .Z(n606) );
  NANDN U889 ( .A(n607), .B(n606), .Z(n608) );
  OR U890 ( .A(n609), .B(n608), .Z(n610) );
  NANDN U891 ( .A(n611), .B(n610), .Z(n612) );
  NANDN U892 ( .A(n613), .B(n612), .Z(n614) );
  OR U893 ( .A(n615), .B(n614), .Z(n616) );
  NANDN U894 ( .A(n617), .B(n616), .Z(n618) );
  NANDN U895 ( .A(n619), .B(n618), .Z(n620) );
  OR U896 ( .A(n621), .B(n620), .Z(n622) );
  NANDN U897 ( .A(n623), .B(n622), .Z(n624) );
  NANDN U898 ( .A(n625), .B(n624), .Z(n626) );
  OR U899 ( .A(n627), .B(n626), .Z(n628) );
  NANDN U900 ( .A(n629), .B(n628), .Z(n630) );
  NANDN U901 ( .A(n631), .B(n630), .Z(n632) );
  OR U902 ( .A(n633), .B(n632), .Z(n634) );
  NANDN U903 ( .A(n635), .B(n634), .Z(n636) );
  NANDN U904 ( .A(n637), .B(n636), .Z(n638) );
  OR U905 ( .A(n639), .B(n638), .Z(n640) );
  NANDN U906 ( .A(n641), .B(n640), .Z(n642) );
  NANDN U907 ( .A(n643), .B(n642), .Z(n644) );
  OR U908 ( .A(n645), .B(n644), .Z(n646) );
  NANDN U909 ( .A(n647), .B(n646), .Z(n648) );
  NANDN U910 ( .A(n649), .B(n648), .Z(n650) );
  OR U911 ( .A(n651), .B(n650), .Z(n652) );
  NANDN U912 ( .A(n653), .B(n652), .Z(n654) );
  NANDN U913 ( .A(n655), .B(n654), .Z(n656) );
  OR U914 ( .A(n657), .B(n656), .Z(n658) );
  NANDN U915 ( .A(n659), .B(n658), .Z(n660) );
  NANDN U916 ( .A(n661), .B(n660), .Z(n662) );
  OR U917 ( .A(n663), .B(n662), .Z(n664) );
  NANDN U918 ( .A(n665), .B(n664), .Z(n666) );
  NANDN U919 ( .A(n667), .B(n666), .Z(n668) );
  OR U920 ( .A(n669), .B(n668), .Z(n670) );
  NANDN U921 ( .A(n671), .B(n670), .Z(n672) );
  NANDN U922 ( .A(n673), .B(n672), .Z(n674) );
  OR U923 ( .A(n675), .B(n674), .Z(n676) );
  NANDN U924 ( .A(n677), .B(n676), .Z(n678) );
  NANDN U925 ( .A(n679), .B(n678), .Z(n680) );
  OR U926 ( .A(n681), .B(n680), .Z(n682) );
  NANDN U927 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U928 ( .A(n685), .B(n684), .Z(n686) );
  OR U929 ( .A(n687), .B(n686), .Z(n688) );
  NANDN U930 ( .A(n689), .B(n688), .Z(n690) );
  NANDN U931 ( .A(n691), .B(n690), .Z(n692) );
  OR U932 ( .A(n693), .B(n692), .Z(n694) );
  NANDN U933 ( .A(n695), .B(n694), .Z(n696) );
  NANDN U934 ( .A(n697), .B(n696), .Z(n698) );
  OR U935 ( .A(n699), .B(n698), .Z(n700) );
  NANDN U936 ( .A(n701), .B(n700), .Z(n702) );
  NANDN U937 ( .A(n703), .B(n702), .Z(n704) );
  OR U938 ( .A(n705), .B(n704), .Z(n706) );
  NANDN U939 ( .A(n707), .B(n706), .Z(n708) );
  NANDN U940 ( .A(n709), .B(n708), .Z(n710) );
  OR U941 ( .A(n711), .B(n710), .Z(n712) );
  NANDN U942 ( .A(n713), .B(n712), .Z(n714) );
  NANDN U943 ( .A(n715), .B(n714), .Z(n716) );
  OR U944 ( .A(n717), .B(n716), .Z(n718) );
  NANDN U945 ( .A(n719), .B(n718), .Z(n720) );
  NANDN U946 ( .A(n721), .B(n720), .Z(n722) );
  OR U947 ( .A(n723), .B(n722), .Z(n724) );
  NANDN U948 ( .A(n725), .B(n724), .Z(n726) );
  NANDN U949 ( .A(n727), .B(n726), .Z(n728) );
  OR U950 ( .A(n729), .B(n728), .Z(n730) );
  NANDN U951 ( .A(n731), .B(n730), .Z(n732) );
  NANDN U952 ( .A(n733), .B(n732), .Z(n734) );
  OR U953 ( .A(n735), .B(n734), .Z(n736) );
  NANDN U954 ( .A(n737), .B(n736), .Z(n738) );
  NANDN U955 ( .A(n739), .B(n738), .Z(n740) );
  OR U956 ( .A(n741), .B(n740), .Z(n742) );
  NANDN U957 ( .A(n743), .B(n742), .Z(n744) );
  NANDN U958 ( .A(n745), .B(n744), .Z(n746) );
  OR U959 ( .A(n747), .B(n746), .Z(n748) );
  NANDN U960 ( .A(n749), .B(n748), .Z(n750) );
  NANDN U961 ( .A(n751), .B(n750), .Z(n752) );
  OR U962 ( .A(n753), .B(n752), .Z(n754) );
  NANDN U963 ( .A(n755), .B(n754), .Z(n756) );
  NANDN U964 ( .A(n757), .B(n756), .Z(n758) );
  OR U965 ( .A(n759), .B(n758), .Z(n760) );
  NANDN U966 ( .A(n761), .B(n760), .Z(n762) );
  NANDN U967 ( .A(n763), .B(n762), .Z(n764) );
  OR U968 ( .A(n765), .B(n764), .Z(n766) );
  NANDN U969 ( .A(n767), .B(n766), .Z(n768) );
  NANDN U970 ( .A(n769), .B(n768), .Z(n770) );
  OR U971 ( .A(n771), .B(n770), .Z(n772) );
  NANDN U972 ( .A(n773), .B(n772), .Z(n774) );
  NANDN U973 ( .A(n775), .B(n774), .Z(n776) );
  OR U974 ( .A(n777), .B(n776), .Z(n778) );
  NANDN U975 ( .A(n779), .B(n778), .Z(n780) );
  NANDN U976 ( .A(n781), .B(n780), .Z(n782) );
  OR U977 ( .A(n783), .B(n782), .Z(n784) );
  NANDN U978 ( .A(n785), .B(n784), .Z(n786) );
  NANDN U979 ( .A(n787), .B(n786), .Z(n788) );
  OR U980 ( .A(n789), .B(n788), .Z(n790) );
  NANDN U981 ( .A(n791), .B(n790), .Z(n792) );
  NANDN U982 ( .A(n793), .B(n792), .Z(n794) );
  OR U983 ( .A(n795), .B(n794), .Z(n796) );
  NANDN U984 ( .A(n797), .B(n796), .Z(n798) );
  NANDN U985 ( .A(n799), .B(n798), .Z(n800) );
  OR U986 ( .A(n801), .B(n800), .Z(n802) );
  NANDN U987 ( .A(n803), .B(n802), .Z(n804) );
  NANDN U988 ( .A(n805), .B(n804), .Z(n806) );
  OR U989 ( .A(n807), .B(n806), .Z(n808) );
  NANDN U990 ( .A(n809), .B(n808), .Z(n810) );
  NANDN U991 ( .A(n811), .B(n810), .Z(n812) );
  OR U992 ( .A(n813), .B(n812), .Z(n814) );
  NANDN U993 ( .A(n815), .B(n814), .Z(n816) );
  NANDN U994 ( .A(n817), .B(n816), .Z(n818) );
  OR U995 ( .A(n819), .B(n818), .Z(n820) );
  NANDN U996 ( .A(n821), .B(n820), .Z(n822) );
  NANDN U997 ( .A(n823), .B(n822), .Z(n824) );
  OR U998 ( .A(n825), .B(n824), .Z(n826) );
  NANDN U999 ( .A(n827), .B(n826), .Z(n828) );
  NANDN U1000 ( .A(n829), .B(n828), .Z(n830) );
  OR U1001 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U1002 ( .A(n833), .B(n832), .Z(n834) );
  NANDN U1003 ( .A(n835), .B(n834), .Z(n836) );
  OR U1004 ( .A(n837), .B(n836), .Z(n838) );
  NANDN U1005 ( .A(n839), .B(n838), .Z(n840) );
  NANDN U1006 ( .A(n841), .B(n840), .Z(n842) );
  OR U1007 ( .A(n843), .B(n842), .Z(n844) );
  NANDN U1008 ( .A(n845), .B(n844), .Z(n846) );
  NANDN U1009 ( .A(n847), .B(n846), .Z(n848) );
  OR U1010 ( .A(n849), .B(n848), .Z(n850) );
  NANDN U1011 ( .A(n851), .B(n850), .Z(n852) );
  NANDN U1012 ( .A(n853), .B(n852), .Z(n854) );
  OR U1013 ( .A(n855), .B(n854), .Z(n856) );
  NANDN U1014 ( .A(n857), .B(n856), .Z(n858) );
  NANDN U1015 ( .A(n859), .B(n858), .Z(n860) );
  OR U1016 ( .A(n861), .B(n860), .Z(n862) );
  NANDN U1017 ( .A(n863), .B(n862), .Z(n864) );
  NANDN U1018 ( .A(n865), .B(n864), .Z(n866) );
  OR U1019 ( .A(n867), .B(n866), .Z(n868) );
  NANDN U1020 ( .A(n869), .B(n868), .Z(n870) );
  NANDN U1021 ( .A(n871), .B(n870), .Z(n872) );
  OR U1022 ( .A(n873), .B(n872), .Z(n874) );
  NANDN U1023 ( .A(n875), .B(n874), .Z(n876) );
  NANDN U1024 ( .A(n877), .B(n876), .Z(n878) );
  OR U1025 ( .A(n879), .B(n878), .Z(n880) );
  NANDN U1026 ( .A(n881), .B(n880), .Z(n882) );
  NANDN U1027 ( .A(n883), .B(n882), .Z(n884) );
  OR U1028 ( .A(n885), .B(n884), .Z(n886) );
  NANDN U1029 ( .A(n887), .B(n886), .Z(n888) );
  NANDN U1030 ( .A(n889), .B(n888), .Z(n890) );
  OR U1031 ( .A(n891), .B(n890), .Z(n892) );
  NANDN U1032 ( .A(n893), .B(n892), .Z(n894) );
  NANDN U1033 ( .A(n895), .B(n894), .Z(n896) );
  OR U1034 ( .A(n897), .B(n896), .Z(n898) );
  NANDN U1035 ( .A(n899), .B(n898), .Z(n900) );
  NANDN U1036 ( .A(n901), .B(n900), .Z(n902) );
  OR U1037 ( .A(n903), .B(n902), .Z(n904) );
  NANDN U1038 ( .A(n905), .B(n904), .Z(n906) );
  NANDN U1039 ( .A(n907), .B(n906), .Z(n909) );
  ANDN U1040 ( .B(x[129]), .A(y[129]), .Z(n908) );
  OR U1041 ( .A(n909), .B(n908), .Z(n910) );
  NANDN U1042 ( .A(n911), .B(n910), .Z(n912) );
  NANDN U1043 ( .A(n913), .B(n912), .Z(n915) );
  ANDN U1044 ( .B(x[131]), .A(y[131]), .Z(n914) );
  OR U1045 ( .A(n915), .B(n914), .Z(n916) );
  NANDN U1046 ( .A(n917), .B(n916), .Z(n918) );
  NANDN U1047 ( .A(n919), .B(n918), .Z(n921) );
  ANDN U1048 ( .B(x[133]), .A(y[133]), .Z(n920) );
  OR U1049 ( .A(n921), .B(n920), .Z(n922) );
  NANDN U1050 ( .A(n923), .B(n922), .Z(n924) );
  NANDN U1051 ( .A(n925), .B(n924), .Z(n927) );
  ANDN U1052 ( .B(x[135]), .A(y[135]), .Z(n926) );
  OR U1053 ( .A(n927), .B(n926), .Z(n928) );
  NANDN U1054 ( .A(n929), .B(n928), .Z(n930) );
  NANDN U1055 ( .A(n931), .B(n930), .Z(n933) );
  ANDN U1056 ( .B(x[137]), .A(y[137]), .Z(n932) );
  OR U1057 ( .A(n933), .B(n932), .Z(n934) );
  NANDN U1058 ( .A(n935), .B(n934), .Z(n936) );
  NANDN U1059 ( .A(n937), .B(n936), .Z(n939) );
  ANDN U1060 ( .B(x[139]), .A(y[139]), .Z(n938) );
  OR U1061 ( .A(n939), .B(n938), .Z(n940) );
  NANDN U1062 ( .A(n941), .B(n940), .Z(n942) );
  NANDN U1063 ( .A(n943), .B(n942), .Z(n945) );
  ANDN U1064 ( .B(x[141]), .A(y[141]), .Z(n944) );
  OR U1065 ( .A(n945), .B(n944), .Z(n946) );
  NANDN U1066 ( .A(n947), .B(n946), .Z(n948) );
  NANDN U1067 ( .A(n949), .B(n948), .Z(n951) );
  ANDN U1068 ( .B(x[143]), .A(y[143]), .Z(n950) );
  OR U1069 ( .A(n951), .B(n950), .Z(n952) );
  NANDN U1070 ( .A(n953), .B(n952), .Z(n954) );
  NANDN U1071 ( .A(n955), .B(n954), .Z(n957) );
  ANDN U1072 ( .B(x[145]), .A(y[145]), .Z(n956) );
  OR U1073 ( .A(n957), .B(n956), .Z(n958) );
  NANDN U1074 ( .A(n959), .B(n958), .Z(n960) );
  NANDN U1075 ( .A(n961), .B(n960), .Z(n963) );
  ANDN U1076 ( .B(x[147]), .A(y[147]), .Z(n962) );
  OR U1077 ( .A(n963), .B(n962), .Z(n964) );
  NANDN U1078 ( .A(n965), .B(n964), .Z(n966) );
  NANDN U1079 ( .A(n967), .B(n966), .Z(n969) );
  ANDN U1080 ( .B(x[149]), .A(y[149]), .Z(n968) );
  OR U1081 ( .A(n969), .B(n968), .Z(n970) );
  NANDN U1082 ( .A(n971), .B(n970), .Z(n972) );
  NANDN U1083 ( .A(n973), .B(n972), .Z(n975) );
  ANDN U1084 ( .B(x[151]), .A(y[151]), .Z(n974) );
  OR U1085 ( .A(n975), .B(n974), .Z(n976) );
  NANDN U1086 ( .A(n977), .B(n976), .Z(n978) );
  NANDN U1087 ( .A(n979), .B(n978), .Z(n981) );
  ANDN U1088 ( .B(x[153]), .A(y[153]), .Z(n980) );
  OR U1089 ( .A(n981), .B(n980), .Z(n982) );
  NANDN U1090 ( .A(n983), .B(n982), .Z(n984) );
  NANDN U1091 ( .A(n985), .B(n984), .Z(n987) );
  ANDN U1092 ( .B(x[155]), .A(y[155]), .Z(n986) );
  OR U1093 ( .A(n987), .B(n986), .Z(n988) );
  NANDN U1094 ( .A(n989), .B(n988), .Z(n990) );
  NANDN U1095 ( .A(n991), .B(n990), .Z(n993) );
  ANDN U1096 ( .B(x[157]), .A(y[157]), .Z(n992) );
  OR U1097 ( .A(n993), .B(n992), .Z(n994) );
  NANDN U1098 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U1099 ( .A(n997), .B(n996), .Z(n999) );
  ANDN U1100 ( .B(x[159]), .A(y[159]), .Z(n998) );
  OR U1101 ( .A(n999), .B(n998), .Z(n1000) );
  NANDN U1102 ( .A(n1001), .B(n1000), .Z(n1002) );
  NANDN U1103 ( .A(n1003), .B(n1002), .Z(n1005) );
  ANDN U1104 ( .B(x[161]), .A(y[161]), .Z(n1004) );
  OR U1105 ( .A(n1005), .B(n1004), .Z(n1006) );
  NANDN U1106 ( .A(n1007), .B(n1006), .Z(n1008) );
  NANDN U1107 ( .A(n1009), .B(n1008), .Z(n1011) );
  ANDN U1108 ( .B(x[163]), .A(y[163]), .Z(n1010) );
  OR U1109 ( .A(n1011), .B(n1010), .Z(n1012) );
  NANDN U1110 ( .A(n1013), .B(n1012), .Z(n1014) );
  NANDN U1111 ( .A(n1015), .B(n1014), .Z(n1017) );
  ANDN U1112 ( .B(x[165]), .A(y[165]), .Z(n1016) );
  OR U1113 ( .A(n1017), .B(n1016), .Z(n1018) );
  NANDN U1114 ( .A(n1019), .B(n1018), .Z(n1020) );
  NANDN U1115 ( .A(n1021), .B(n1020), .Z(n1023) );
  ANDN U1116 ( .B(x[167]), .A(y[167]), .Z(n1022) );
  OR U1117 ( .A(n1023), .B(n1022), .Z(n1024) );
  NANDN U1118 ( .A(n1025), .B(n1024), .Z(n1026) );
  NANDN U1119 ( .A(n1027), .B(n1026), .Z(n1029) );
  ANDN U1120 ( .B(x[169]), .A(y[169]), .Z(n1028) );
  OR U1121 ( .A(n1029), .B(n1028), .Z(n1030) );
  NANDN U1122 ( .A(n1031), .B(n1030), .Z(n1032) );
  NANDN U1123 ( .A(n1033), .B(n1032), .Z(n1035) );
  ANDN U1124 ( .B(x[171]), .A(y[171]), .Z(n1034) );
  OR U1125 ( .A(n1035), .B(n1034), .Z(n1036) );
  NANDN U1126 ( .A(n1037), .B(n1036), .Z(n1038) );
  NANDN U1127 ( .A(n1039), .B(n1038), .Z(n1041) );
  ANDN U1128 ( .B(x[173]), .A(y[173]), .Z(n1040) );
  OR U1129 ( .A(n1041), .B(n1040), .Z(n1042) );
  NANDN U1130 ( .A(n1043), .B(n1042), .Z(n1044) );
  NANDN U1131 ( .A(n1045), .B(n1044), .Z(n1047) );
  ANDN U1132 ( .B(x[175]), .A(y[175]), .Z(n1046) );
  OR U1133 ( .A(n1047), .B(n1046), .Z(n1048) );
  NANDN U1134 ( .A(n1049), .B(n1048), .Z(n1050) );
  NANDN U1135 ( .A(n1051), .B(n1050), .Z(n1053) );
  ANDN U1136 ( .B(x[177]), .A(y[177]), .Z(n1052) );
  OR U1137 ( .A(n1053), .B(n1052), .Z(n1054) );
  NANDN U1138 ( .A(n1055), .B(n1054), .Z(n1056) );
  NANDN U1139 ( .A(n1057), .B(n1056), .Z(n1059) );
  ANDN U1140 ( .B(x[179]), .A(y[179]), .Z(n1058) );
  OR U1141 ( .A(n1059), .B(n1058), .Z(n1060) );
  NANDN U1142 ( .A(n1061), .B(n1060), .Z(n1062) );
  NANDN U1143 ( .A(n1063), .B(n1062), .Z(n1065) );
  ANDN U1144 ( .B(x[181]), .A(y[181]), .Z(n1064) );
  OR U1145 ( .A(n1065), .B(n1064), .Z(n1066) );
  NANDN U1146 ( .A(n1067), .B(n1066), .Z(n1068) );
  NANDN U1147 ( .A(n1069), .B(n1068), .Z(n1071) );
  ANDN U1148 ( .B(x[183]), .A(y[183]), .Z(n1070) );
  OR U1149 ( .A(n1071), .B(n1070), .Z(n1072) );
  NANDN U1150 ( .A(n1073), .B(n1072), .Z(n1074) );
  NANDN U1151 ( .A(n1075), .B(n1074), .Z(n1077) );
  ANDN U1152 ( .B(x[185]), .A(y[185]), .Z(n1076) );
  OR U1153 ( .A(n1077), .B(n1076), .Z(n1078) );
  NANDN U1154 ( .A(n1079), .B(n1078), .Z(n1080) );
  NANDN U1155 ( .A(n1081), .B(n1080), .Z(n1083) );
  ANDN U1156 ( .B(x[187]), .A(y[187]), .Z(n1082) );
  OR U1157 ( .A(n1083), .B(n1082), .Z(n1084) );
  NANDN U1158 ( .A(n1085), .B(n1084), .Z(n1086) );
  NANDN U1159 ( .A(n1087), .B(n1086), .Z(n1089) );
  ANDN U1160 ( .B(x[189]), .A(y[189]), .Z(n1088) );
  OR U1161 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U1162 ( .A(n1091), .B(n1090), .Z(n1092) );
  NANDN U1163 ( .A(n1093), .B(n1092), .Z(n1095) );
  ANDN U1164 ( .B(x[191]), .A(y[191]), .Z(n1094) );
  OR U1165 ( .A(n1095), .B(n1094), .Z(n1096) );
  NANDN U1166 ( .A(n1097), .B(n1096), .Z(n1098) );
  NANDN U1167 ( .A(n1099), .B(n1098), .Z(n1101) );
  ANDN U1168 ( .B(x[193]), .A(y[193]), .Z(n1100) );
  OR U1169 ( .A(n1101), .B(n1100), .Z(n1102) );
  NANDN U1170 ( .A(n1103), .B(n1102), .Z(n1104) );
  NANDN U1171 ( .A(n1105), .B(n1104), .Z(n1107) );
  ANDN U1172 ( .B(x[195]), .A(y[195]), .Z(n1106) );
  OR U1173 ( .A(n1107), .B(n1106), .Z(n1108) );
  NANDN U1174 ( .A(n1109), .B(n1108), .Z(n1110) );
  NANDN U1175 ( .A(n1111), .B(n1110), .Z(n1113) );
  ANDN U1176 ( .B(x[197]), .A(y[197]), .Z(n1112) );
  OR U1177 ( .A(n1113), .B(n1112), .Z(n1114) );
  NANDN U1178 ( .A(n1115), .B(n1114), .Z(n1116) );
  NANDN U1179 ( .A(n1117), .B(n1116), .Z(n1119) );
  ANDN U1180 ( .B(x[199]), .A(y[199]), .Z(n1118) );
  OR U1181 ( .A(n1119), .B(n1118), .Z(n1120) );
  NANDN U1182 ( .A(n1121), .B(n1120), .Z(n1122) );
  NANDN U1183 ( .A(n1123), .B(n1122), .Z(n1125) );
  ANDN U1184 ( .B(x[201]), .A(y[201]), .Z(n1124) );
  OR U1185 ( .A(n1125), .B(n1124), .Z(n1126) );
  NANDN U1186 ( .A(n1127), .B(n1126), .Z(n1128) );
  NANDN U1187 ( .A(n1129), .B(n1128), .Z(n1131) );
  ANDN U1188 ( .B(x[203]), .A(y[203]), .Z(n1130) );
  OR U1189 ( .A(n1131), .B(n1130), .Z(n1132) );
  NANDN U1190 ( .A(n1133), .B(n1132), .Z(n1134) );
  NANDN U1191 ( .A(n1135), .B(n1134), .Z(n1137) );
  ANDN U1192 ( .B(x[205]), .A(y[205]), .Z(n1136) );
  OR U1193 ( .A(n1137), .B(n1136), .Z(n1138) );
  NANDN U1194 ( .A(n1139), .B(n1138), .Z(n1140) );
  NANDN U1195 ( .A(n1141), .B(n1140), .Z(n1143) );
  ANDN U1196 ( .B(x[207]), .A(y[207]), .Z(n1142) );
  OR U1197 ( .A(n1143), .B(n1142), .Z(n1144) );
  NANDN U1198 ( .A(n1145), .B(n1144), .Z(n1146) );
  NANDN U1199 ( .A(n1147), .B(n1146), .Z(n1149) );
  ANDN U1200 ( .B(x[209]), .A(y[209]), .Z(n1148) );
  OR U1201 ( .A(n1149), .B(n1148), .Z(n1150) );
  NANDN U1202 ( .A(n1151), .B(n1150), .Z(n1152) );
  NANDN U1203 ( .A(n1153), .B(n1152), .Z(n1155) );
  ANDN U1204 ( .B(x[211]), .A(y[211]), .Z(n1154) );
  OR U1205 ( .A(n1155), .B(n1154), .Z(n1156) );
  NANDN U1206 ( .A(n1157), .B(n1156), .Z(n1158) );
  NANDN U1207 ( .A(n1159), .B(n1158), .Z(n1161) );
  ANDN U1208 ( .B(x[213]), .A(y[213]), .Z(n1160) );
  OR U1209 ( .A(n1161), .B(n1160), .Z(n1162) );
  NANDN U1210 ( .A(n1163), .B(n1162), .Z(n1164) );
  NANDN U1211 ( .A(n1165), .B(n1164), .Z(n1167) );
  ANDN U1212 ( .B(x[215]), .A(y[215]), .Z(n1166) );
  OR U1213 ( .A(n1167), .B(n1166), .Z(n1168) );
  NANDN U1214 ( .A(n1169), .B(n1168), .Z(n1170) );
  NANDN U1215 ( .A(n1171), .B(n1170), .Z(n1173) );
  ANDN U1216 ( .B(x[217]), .A(y[217]), .Z(n1172) );
  OR U1217 ( .A(n1173), .B(n1172), .Z(n1174) );
  NANDN U1218 ( .A(n1175), .B(n1174), .Z(n1176) );
  NANDN U1219 ( .A(n1177), .B(n1176), .Z(n1179) );
  ANDN U1220 ( .B(x[219]), .A(y[219]), .Z(n1178) );
  OR U1221 ( .A(n1179), .B(n1178), .Z(n1180) );
  NANDN U1222 ( .A(n1181), .B(n1180), .Z(n1182) );
  NANDN U1223 ( .A(n1183), .B(n1182), .Z(n1185) );
  ANDN U1224 ( .B(x[221]), .A(y[221]), .Z(n1184) );
  OR U1225 ( .A(n1185), .B(n1184), .Z(n1186) );
  NANDN U1226 ( .A(n1187), .B(n1186), .Z(n1188) );
  NANDN U1227 ( .A(n1189), .B(n1188), .Z(n1191) );
  ANDN U1228 ( .B(x[223]), .A(y[223]), .Z(n1190) );
  OR U1229 ( .A(n1191), .B(n1190), .Z(n1192) );
  NANDN U1230 ( .A(n1193), .B(n1192), .Z(n1194) );
  NANDN U1231 ( .A(n1195), .B(n1194), .Z(n1197) );
  ANDN U1232 ( .B(x[225]), .A(y[225]), .Z(n1196) );
  OR U1233 ( .A(n1197), .B(n1196), .Z(n1198) );
  NANDN U1234 ( .A(n1199), .B(n1198), .Z(n1200) );
  NANDN U1235 ( .A(n1201), .B(n1200), .Z(n1203) );
  ANDN U1236 ( .B(x[227]), .A(y[227]), .Z(n1202) );
  OR U1237 ( .A(n1203), .B(n1202), .Z(n1204) );
  NANDN U1238 ( .A(n1205), .B(n1204), .Z(n1206) );
  NANDN U1239 ( .A(n1207), .B(n1206), .Z(n1209) );
  ANDN U1240 ( .B(x[229]), .A(y[229]), .Z(n1208) );
  OR U1241 ( .A(n1209), .B(n1208), .Z(n1210) );
  NANDN U1242 ( .A(n1211), .B(n1210), .Z(n1212) );
  NANDN U1243 ( .A(n1213), .B(n1212), .Z(n1215) );
  ANDN U1244 ( .B(x[231]), .A(y[231]), .Z(n1214) );
  OR U1245 ( .A(n1215), .B(n1214), .Z(n1216) );
  NANDN U1246 ( .A(n1217), .B(n1216), .Z(n1218) );
  NANDN U1247 ( .A(n1219), .B(n1218), .Z(n1221) );
  ANDN U1248 ( .B(x[233]), .A(y[233]), .Z(n1220) );
  OR U1249 ( .A(n1221), .B(n1220), .Z(n1222) );
  NANDN U1250 ( .A(n1223), .B(n1222), .Z(n1224) );
  NANDN U1251 ( .A(n1225), .B(n1224), .Z(n1227) );
  ANDN U1252 ( .B(x[235]), .A(y[235]), .Z(n1226) );
  OR U1253 ( .A(n1227), .B(n1226), .Z(n1228) );
  NANDN U1254 ( .A(n1229), .B(n1228), .Z(n1230) );
  NANDN U1255 ( .A(n1231), .B(n1230), .Z(n1233) );
  ANDN U1256 ( .B(x[237]), .A(y[237]), .Z(n1232) );
  OR U1257 ( .A(n1233), .B(n1232), .Z(n1234) );
  NANDN U1258 ( .A(n1235), .B(n1234), .Z(n1236) );
  NANDN U1259 ( .A(n1237), .B(n1236), .Z(n1239) );
  ANDN U1260 ( .B(x[239]), .A(y[239]), .Z(n1238) );
  OR U1261 ( .A(n1239), .B(n1238), .Z(n1240) );
  NANDN U1262 ( .A(n1241), .B(n1240), .Z(n1242) );
  NANDN U1263 ( .A(n1243), .B(n1242), .Z(n1245) );
  ANDN U1264 ( .B(x[241]), .A(y[241]), .Z(n1244) );
  OR U1265 ( .A(n1245), .B(n1244), .Z(n1246) );
  NANDN U1266 ( .A(n1247), .B(n1246), .Z(n1248) );
  NANDN U1267 ( .A(n1249), .B(n1248), .Z(n1251) );
  ANDN U1268 ( .B(x[243]), .A(y[243]), .Z(n1250) );
  OR U1269 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U1270 ( .A(n1253), .B(n1252), .Z(n1254) );
  NANDN U1271 ( .A(n1255), .B(n1254), .Z(n1257) );
  ANDN U1272 ( .B(x[245]), .A(y[245]), .Z(n1256) );
  OR U1273 ( .A(n1257), .B(n1256), .Z(n1258) );
  NANDN U1274 ( .A(n1259), .B(n1258), .Z(n1260) );
  NANDN U1275 ( .A(n1261), .B(n1260), .Z(n1263) );
  ANDN U1276 ( .B(x[247]), .A(y[247]), .Z(n1262) );
  OR U1277 ( .A(n1263), .B(n1262), .Z(n1264) );
  NANDN U1278 ( .A(n1265), .B(n1264), .Z(n1266) );
  NANDN U1279 ( .A(n1267), .B(n1266), .Z(n1269) );
  ANDN U1280 ( .B(x[249]), .A(y[249]), .Z(n1268) );
  OR U1281 ( .A(n1269), .B(n1268), .Z(n1270) );
  NANDN U1282 ( .A(n1271), .B(n1270), .Z(n1272) );
  NANDN U1283 ( .A(n1273), .B(n1272), .Z(n1275) );
  ANDN U1284 ( .B(x[251]), .A(y[251]), .Z(n1274) );
  OR U1285 ( .A(n1275), .B(n1274), .Z(n1276) );
  NANDN U1286 ( .A(n1277), .B(n1276), .Z(n1278) );
  NANDN U1287 ( .A(n1279), .B(n1278), .Z(n1281) );
  ANDN U1288 ( .B(x[253]), .A(y[253]), .Z(n1280) );
  OR U1289 ( .A(n1281), .B(n1280), .Z(n1282) );
  NANDN U1290 ( .A(n1283), .B(n1282), .Z(n1284) );
  NANDN U1291 ( .A(n1285), .B(n1284), .Z(n1286) );
  NANDN U1292 ( .A(n1287), .B(n1286), .Z(n1289) );
  NAND U1293 ( .A(n1287), .B(g), .Z(n1288) );
  NAND U1294 ( .A(n1289), .B(n1288), .Z(n4) );
endmodule

