
module hamming_N160_CC2 ( clk, rst, x, y, o );
  input [79:0] x;
  input [79:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U83 ( .A(n130), .B(n129), .Z(n1) );
  NANDN U84 ( .A(n128), .B(n127), .Z(n2) );
  NAND U85 ( .A(n1), .B(n2), .Z(n361) );
  NAND U86 ( .A(n202), .B(n201), .Z(n3) );
  NANDN U87 ( .A(n200), .B(n199), .Z(n4) );
  AND U88 ( .A(n3), .B(n4), .Z(n334) );
  NAND U89 ( .A(n337), .B(n336), .Z(n5) );
  XOR U90 ( .A(n336), .B(n337), .Z(n6) );
  NAND U91 ( .A(n6), .B(n335), .Z(n7) );
  NAND U92 ( .A(n5), .B(n7), .Z(n425) );
  NANDN U93 ( .A(n124), .B(n123), .Z(n8) );
  NANDN U94 ( .A(n126), .B(n125), .Z(n9) );
  NAND U95 ( .A(n8), .B(n9), .Z(n366) );
  NANDN U96 ( .A(n282), .B(n281), .Z(n10) );
  NANDN U97 ( .A(n284), .B(n283), .Z(n11) );
  AND U98 ( .A(n10), .B(n11), .Z(n363) );
  NANDN U99 ( .A(n224), .B(n223), .Z(n12) );
  NANDN U100 ( .A(n226), .B(n225), .Z(n13) );
  AND U101 ( .A(n12), .B(n13), .Z(n337) );
  NAND U102 ( .A(n361), .B(n359), .Z(n14) );
  XOR U103 ( .A(n359), .B(n361), .Z(n15) );
  NANDN U104 ( .A(n360), .B(n15), .Z(n16) );
  NAND U105 ( .A(n14), .B(n16), .Z(n437) );
  NANDN U106 ( .A(n235), .B(n234), .Z(n17) );
  NANDN U107 ( .A(n237), .B(n236), .Z(n18) );
  NAND U108 ( .A(n17), .B(n18), .Z(n328) );
  OR U109 ( .A(n331), .B(n332), .Z(n19) );
  NANDN U110 ( .A(n334), .B(n333), .Z(n20) );
  NAND U111 ( .A(n19), .B(n20), .Z(n427) );
  XOR U112 ( .A(n423), .B(n422), .Z(n21) );
  NANDN U113 ( .A(n421), .B(n21), .Z(n22) );
  NAND U114 ( .A(n423), .B(n422), .Z(n23) );
  AND U115 ( .A(n22), .B(n23), .Z(n476) );
  NANDN U116 ( .A(n120), .B(n119), .Z(n24) );
  NANDN U117 ( .A(n122), .B(n121), .Z(n25) );
  NAND U118 ( .A(n24), .B(n25), .Z(n365) );
  NAND U119 ( .A(n274), .B(n273), .Z(n26) );
  NANDN U120 ( .A(n272), .B(n271), .Z(n27) );
  NAND U121 ( .A(n26), .B(n27), .Z(n364) );
  NANDN U122 ( .A(n297), .B(n296), .Z(n28) );
  NANDN U123 ( .A(n299), .B(n298), .Z(n29) );
  AND U124 ( .A(n28), .B(n29), .Z(n355) );
  NANDN U125 ( .A(n138), .B(n137), .Z(n30) );
  NANDN U126 ( .A(n140), .B(n139), .Z(n31) );
  AND U127 ( .A(n30), .B(n31), .Z(n360) );
  NANDN U128 ( .A(n220), .B(n219), .Z(n32) );
  NANDN U129 ( .A(n222), .B(n221), .Z(n33) );
  AND U130 ( .A(n32), .B(n33), .Z(n336) );
  NANDN U131 ( .A(n251), .B(n250), .Z(n34) );
  NANDN U132 ( .A(n253), .B(n252), .Z(n35) );
  AND U133 ( .A(n34), .B(n35), .Z(n396) );
  NANDN U134 ( .A(n143), .B(n142), .Z(n36) );
  NANDN U135 ( .A(n145), .B(n144), .Z(n37) );
  AND U136 ( .A(n36), .B(n37), .Z(n345) );
  XOR U137 ( .A(n404), .B(n403), .Z(n38) );
  NANDN U138 ( .A(n402), .B(n38), .Z(n39) );
  NAND U139 ( .A(n404), .B(n403), .Z(n40) );
  AND U140 ( .A(n39), .B(n40), .Z(n446) );
  NAND U141 ( .A(n434), .B(n433), .Z(n41) );
  NANDN U142 ( .A(n432), .B(n431), .Z(n42) );
  NAND U143 ( .A(n41), .B(n42), .Z(n468) );
  NAND U144 ( .A(n478), .B(n476), .Z(n43) );
  XOR U145 ( .A(n476), .B(n478), .Z(n44) );
  NANDN U146 ( .A(n477), .B(n44), .Z(n45) );
  NAND U147 ( .A(n43), .B(n45), .Z(n481) );
  NANDN U148 ( .A(n264), .B(n263), .Z(n46) );
  NANDN U149 ( .A(n266), .B(n265), .Z(n47) );
  AND U150 ( .A(n46), .B(n47), .Z(n349) );
  NANDN U151 ( .A(n287), .B(n286), .Z(n48) );
  NANDN U152 ( .A(n289), .B(n288), .Z(n49) );
  NAND U153 ( .A(n48), .B(n49), .Z(n356) );
  XOR U154 ( .A(n358), .B(oglobal[1]), .Z(n50) );
  XNOR U155 ( .A(n357), .B(n50), .Z(n387) );
  XOR U156 ( .A(n364), .B(n362), .Z(n51) );
  NANDN U157 ( .A(n363), .B(n51), .Z(n52) );
  NAND U158 ( .A(n364), .B(n362), .Z(n53) );
  AND U159 ( .A(n52), .B(n53), .Z(n436) );
  XOR U160 ( .A(n240), .B(n239), .Z(n54) );
  NANDN U161 ( .A(n238), .B(n54), .Z(n55) );
  NAND U162 ( .A(n240), .B(n239), .Z(n56) );
  AND U163 ( .A(n55), .B(n56), .Z(n325) );
  XOR U164 ( .A(n155), .B(n154), .Z(n57) );
  NANDN U165 ( .A(n153), .B(n57), .Z(n58) );
  NAND U166 ( .A(n155), .B(n154), .Z(n59) );
  AND U167 ( .A(n58), .B(n59), .Z(n381) );
  XOR U168 ( .A(n394), .B(n392), .Z(n60) );
  NANDN U169 ( .A(n393), .B(n60), .Z(n61) );
  NAND U170 ( .A(n394), .B(n392), .Z(n62) );
  AND U171 ( .A(n61), .B(n62), .Z(n421) );
  NAND U172 ( .A(n346), .B(n344), .Z(n63) );
  XOR U173 ( .A(n344), .B(n346), .Z(n64) );
  NANDN U174 ( .A(n345), .B(n64), .Z(n65) );
  NAND U175 ( .A(n63), .B(n65), .Z(n443) );
  NAND U176 ( .A(n317), .B(n316), .Z(n66) );
  XOR U177 ( .A(n316), .B(n317), .Z(n67) );
  NANDN U178 ( .A(n318), .B(n67), .Z(n68) );
  NAND U179 ( .A(n66), .B(n68), .Z(n412) );
  NAND U180 ( .A(n457), .B(n456), .Z(n69) );
  XOR U181 ( .A(n456), .B(n457), .Z(n70) );
  NANDN U182 ( .A(n458), .B(n70), .Z(n71) );
  NAND U183 ( .A(n69), .B(n71), .Z(n484) );
  XOR U184 ( .A(n483), .B(n481), .Z(n72) );
  NAND U185 ( .A(n72), .B(n482), .Z(n73) );
  NAND U186 ( .A(n483), .B(n481), .Z(n74) );
  AND U187 ( .A(n73), .B(n74), .Z(n494) );
  NANDN U188 ( .A(n260), .B(n259), .Z(n75) );
  NANDN U189 ( .A(n262), .B(n261), .Z(n76) );
  AND U190 ( .A(n75), .B(n76), .Z(n348) );
  NANDN U191 ( .A(n228), .B(n227), .Z(n77) );
  NANDN U192 ( .A(n230), .B(n229), .Z(n78) );
  AND U193 ( .A(n77), .B(n78), .Z(n335) );
  NAND U194 ( .A(n248), .B(n247), .Z(n79) );
  XOR U195 ( .A(n247), .B(n248), .Z(n80) );
  NANDN U196 ( .A(n249), .B(n80), .Z(n81) );
  NAND U197 ( .A(n79), .B(n81), .Z(n395) );
  NAND U198 ( .A(n218), .B(n217), .Z(n82) );
  XOR U199 ( .A(n217), .B(n218), .Z(n83) );
  NAND U200 ( .A(n83), .B(n216), .Z(n84) );
  NAND U201 ( .A(n82), .B(n84), .Z(n393) );
  NAND U202 ( .A(n356), .B(n354), .Z(n85) );
  XOR U203 ( .A(n354), .B(n356), .Z(n86) );
  NANDN U204 ( .A(n355), .B(n86), .Z(n87) );
  NAND U205 ( .A(n85), .B(n87), .Z(n438) );
  NANDN U206 ( .A(n268), .B(n267), .Z(n88) );
  NANDN U207 ( .A(n270), .B(n269), .Z(n89) );
  NAND U208 ( .A(n88), .B(n89), .Z(n375) );
  NAND U209 ( .A(n358), .B(oglobal[1]), .Z(n90) );
  XOR U210 ( .A(oglobal[1]), .B(n358), .Z(n91) );
  NANDN U211 ( .A(n357), .B(n91), .Z(n92) );
  NAND U212 ( .A(n90), .B(n92), .Z(n415) );
  XOR U213 ( .A(n436), .B(n435), .Z(n93) );
  NANDN U214 ( .A(n437), .B(n93), .Z(n94) );
  NAND U215 ( .A(n436), .B(n435), .Z(n95) );
  AND U216 ( .A(n94), .B(n95), .Z(n471) );
  NAND U217 ( .A(n445), .B(n444), .Z(n96) );
  XOR U218 ( .A(n444), .B(n445), .Z(n97) );
  NAND U219 ( .A(n97), .B(n443), .Z(n98) );
  NAND U220 ( .A(n96), .B(n98), .Z(n465) );
  XOR U221 ( .A(n446), .B(n447), .Z(n99) );
  NANDN U222 ( .A(n448), .B(n99), .Z(n100) );
  NAND U223 ( .A(n446), .B(n447), .Z(n101) );
  AND U224 ( .A(n100), .B(n101), .Z(n457) );
  NAND U225 ( .A(n414), .B(n413), .Z(n102) );
  XOR U226 ( .A(n413), .B(n414), .Z(n103) );
  NAND U227 ( .A(n103), .B(n412), .Z(n104) );
  NAND U228 ( .A(n102), .B(n104), .Z(n459) );
  ANDN U229 ( .B(n495), .A(n496), .Z(n105) );
  NANDN U230 ( .A(n494), .B(n493), .Z(n106) );
  AND U231 ( .A(n105), .B(n106), .Z(n498) );
  XNOR U232 ( .A(x[22]), .B(y[22]), .Z(n140) );
  XNOR U233 ( .A(x[26]), .B(y[26]), .Z(n138) );
  XOR U234 ( .A(x[24]), .B(y[24]), .Z(n137) );
  XNOR U235 ( .A(n138), .B(n137), .Z(n139) );
  XNOR U236 ( .A(n140), .B(n139), .Z(n267) );
  XNOR U237 ( .A(x[16]), .B(y[16]), .Z(n122) );
  XNOR U238 ( .A(x[20]), .B(y[20]), .Z(n120) );
  XOR U239 ( .A(x[18]), .B(y[18]), .Z(n119) );
  XNOR U240 ( .A(n120), .B(n119), .Z(n121) );
  XOR U241 ( .A(n122), .B(n121), .Z(n268) );
  XNOR U242 ( .A(n267), .B(n268), .Z(n269) );
  XNOR U243 ( .A(x[10]), .B(y[10]), .Z(n126) );
  XNOR U244 ( .A(x[14]), .B(y[14]), .Z(n124) );
  XOR U245 ( .A(x[12]), .B(y[12]), .Z(n123) );
  XNOR U246 ( .A(n124), .B(n123), .Z(n125) );
  XOR U247 ( .A(n126), .B(n125), .Z(n270) );
  XOR U248 ( .A(n269), .B(n270), .Z(n306) );
  XNOR U249 ( .A(x[74]), .B(y[74]), .Z(n299) );
  XNOR U250 ( .A(x[78]), .B(y[78]), .Z(n297) );
  XOR U251 ( .A(x[76]), .B(y[76]), .Z(n296) );
  XNOR U252 ( .A(n297), .B(n296), .Z(n298) );
  XOR U253 ( .A(n299), .B(n298), .Z(n240) );
  XNOR U254 ( .A(x[46]), .B(y[46]), .Z(n145) );
  XNOR U255 ( .A(x[50]), .B(y[50]), .Z(n143) );
  XOR U256 ( .A(x[48]), .B(y[48]), .Z(n142) );
  XNOR U257 ( .A(n143), .B(n142), .Z(n144) );
  XNOR U258 ( .A(n145), .B(n144), .Z(n238) );
  XNOR U259 ( .A(x[56]), .B(y[56]), .Z(n282) );
  XOR U260 ( .A(x[54]), .B(y[54]), .Z(n281) );
  XNOR U261 ( .A(n282), .B(n281), .Z(n283) );
  XNOR U262 ( .A(x[52]), .B(y[52]), .Z(n284) );
  XOR U263 ( .A(n283), .B(n284), .Z(n239) );
  XOR U264 ( .A(n238), .B(n239), .Z(n107) );
  XOR U265 ( .A(n240), .B(n107), .Z(n304) );
  IV U266 ( .A(n304), .Z(n302) );
  XNOR U267 ( .A(x[44]), .B(y[44]), .Z(n272) );
  XOR U268 ( .A(x[42]), .B(y[42]), .Z(n271) );
  XNOR U269 ( .A(n272), .B(n271), .Z(n273) );
  XOR U270 ( .A(x[40]), .B(y[40]), .Z(n274) );
  XNOR U271 ( .A(n273), .B(n274), .Z(n241) );
  XNOR U272 ( .A(x[34]), .B(y[34]), .Z(n278) );
  XNOR U273 ( .A(x[38]), .B(y[38]), .Z(n276) );
  XNOR U274 ( .A(x[36]), .B(y[36]), .Z(n275) );
  XOR U275 ( .A(n276), .B(n275), .Z(n277) );
  XOR U276 ( .A(n278), .B(n277), .Z(n242) );
  XOR U277 ( .A(n241), .B(n242), .Z(n243) );
  XNOR U278 ( .A(x[32]), .B(y[32]), .Z(n128) );
  XOR U279 ( .A(x[30]), .B(y[30]), .Z(n127) );
  XNOR U280 ( .A(n128), .B(n127), .Z(n129) );
  XOR U281 ( .A(x[28]), .B(y[28]), .Z(n130) );
  XNOR U282 ( .A(n129), .B(n130), .Z(n244) );
  XNOR U283 ( .A(n243), .B(n244), .Z(n303) );
  XOR U284 ( .A(n302), .B(n303), .Z(n108) );
  XNOR U285 ( .A(n306), .B(n108), .Z(n311) );
  XNOR U286 ( .A(x[55]), .B(y[55]), .Z(n177) );
  XNOR U287 ( .A(x[75]), .B(y[75]), .Z(n175) );
  XNOR U288 ( .A(x[53]), .B(y[53]), .Z(n174) );
  XNOR U289 ( .A(n175), .B(n174), .Z(n176) );
  XOR U290 ( .A(n177), .B(n176), .Z(n218) );
  XNOR U291 ( .A(x[63]), .B(y[63]), .Z(n190) );
  XNOR U292 ( .A(x[71]), .B(y[71]), .Z(n188) );
  XNOR U293 ( .A(x[61]), .B(y[61]), .Z(n187) );
  XNOR U294 ( .A(n188), .B(n187), .Z(n189) );
  XOR U295 ( .A(n190), .B(n189), .Z(n217) );
  XNOR U296 ( .A(x[59]), .B(y[59]), .Z(n196) );
  XNOR U297 ( .A(x[73]), .B(y[73]), .Z(n194) );
  XNOR U298 ( .A(x[57]), .B(y[57]), .Z(n193) );
  XNOR U299 ( .A(n194), .B(n193), .Z(n195) );
  XOR U300 ( .A(n196), .B(n195), .Z(n216) );
  XNOR U301 ( .A(n217), .B(n216), .Z(n109) );
  XOR U302 ( .A(n218), .B(n109), .Z(n155) );
  XNOR U303 ( .A(x[31]), .B(y[31]), .Z(n213) );
  XNOR U304 ( .A(x[29]), .B(y[29]), .Z(n211) );
  XOR U305 ( .A(x[27]), .B(y[27]), .Z(n209) );
  XNOR U306 ( .A(n211), .B(n209), .Z(n212) );
  XNOR U307 ( .A(n213), .B(n212), .Z(n250) );
  XNOR U308 ( .A(x[37]), .B(y[37]), .Z(n226) );
  XNOR U309 ( .A(x[35]), .B(y[35]), .Z(n224) );
  XOR U310 ( .A(x[33]), .B(y[33]), .Z(n223) );
  XNOR U311 ( .A(n224), .B(n223), .Z(n225) );
  XOR U312 ( .A(n226), .B(n225), .Z(n251) );
  XNOR U313 ( .A(n250), .B(n251), .Z(n252) );
  XNOR U314 ( .A(x[43]), .B(y[43]), .Z(n230) );
  XNOR U315 ( .A(x[41]), .B(y[41]), .Z(n228) );
  XOR U316 ( .A(x[39]), .B(y[39]), .Z(n227) );
  XNOR U317 ( .A(n228), .B(n227), .Z(n229) );
  XOR U318 ( .A(n230), .B(n229), .Z(n253) );
  XNOR U319 ( .A(n252), .B(n253), .Z(n153) );
  XNOR U320 ( .A(x[47]), .B(y[47]), .Z(n222) );
  XNOR U321 ( .A(x[79]), .B(y[79]), .Z(n220) );
  XOR U322 ( .A(x[45]), .B(y[45]), .Z(n219) );
  XNOR U323 ( .A(n220), .B(n219), .Z(n221) );
  XOR U324 ( .A(n222), .B(n221), .Z(n249) );
  XNOR U325 ( .A(x[51]), .B(y[51]), .Z(n171) );
  XNOR U326 ( .A(x[77]), .B(y[77]), .Z(n169) );
  XNOR U327 ( .A(x[49]), .B(y[49]), .Z(n168) );
  XNOR U328 ( .A(n169), .B(n168), .Z(n170) );
  XOR U329 ( .A(n171), .B(n170), .Z(n248) );
  XNOR U330 ( .A(x[67]), .B(y[67]), .Z(n165) );
  XNOR U331 ( .A(x[69]), .B(y[69]), .Z(n163) );
  XNOR U332 ( .A(x[65]), .B(y[65]), .Z(n162) );
  XNOR U333 ( .A(n163), .B(n162), .Z(n164) );
  XOR U334 ( .A(n165), .B(n164), .Z(n247) );
  XNOR U335 ( .A(n248), .B(n247), .Z(n110) );
  XNOR U336 ( .A(n249), .B(n110), .Z(n154) );
  XOR U337 ( .A(n153), .B(n154), .Z(n111) );
  XOR U338 ( .A(n155), .B(n111), .Z(n310) );
  XOR U339 ( .A(n311), .B(n310), .Z(n313) );
  XNOR U340 ( .A(x[64]), .B(y[64]), .Z(n116) );
  XNOR U341 ( .A(x[68]), .B(y[68]), .Z(n114) );
  XNOR U342 ( .A(x[66]), .B(y[66]), .Z(n113) );
  XNOR U343 ( .A(n114), .B(n113), .Z(n115) );
  XOR U344 ( .A(n116), .B(n115), .Z(n183) );
  XNOR U345 ( .A(x[58]), .B(y[58]), .Z(n134) );
  XNOR U346 ( .A(x[62]), .B(y[62]), .Z(n132) );
  XNOR U347 ( .A(x[60]), .B(y[60]), .Z(n131) );
  XNOR U348 ( .A(n132), .B(n131), .Z(n133) );
  XOR U349 ( .A(n134), .B(n133), .Z(n182) );
  IV U350 ( .A(n182), .Z(n180) );
  XNOR U351 ( .A(x[70]), .B(y[70]), .Z(n256) );
  XOR U352 ( .A(x[72]), .B(y[72]), .Z(n254) );
  XNOR U353 ( .A(oglobal[0]), .B(n254), .Z(n255) );
  XOR U354 ( .A(n256), .B(n255), .Z(n181) );
  XOR U355 ( .A(n180), .B(n181), .Z(n112) );
  XOR U356 ( .A(n183), .B(n112), .Z(n150) );
  XNOR U357 ( .A(x[13]), .B(y[13]), .Z(n293) );
  XNOR U358 ( .A(x[11]), .B(y[11]), .Z(n291) );
  XNOR U359 ( .A(x[9]), .B(y[9]), .Z(n290) );
  XOR U360 ( .A(n291), .B(n290), .Z(n292) );
  XNOR U361 ( .A(n293), .B(n292), .Z(n234) );
  XNOR U362 ( .A(x[19]), .B(y[19]), .Z(n206) );
  XNOR U363 ( .A(x[17]), .B(y[17]), .Z(n204) );
  XNOR U364 ( .A(x[15]), .B(y[15]), .Z(n203) );
  XOR U365 ( .A(n204), .B(n203), .Z(n205) );
  XOR U366 ( .A(n206), .B(n205), .Z(n235) );
  XNOR U367 ( .A(n234), .B(n235), .Z(n236) );
  XNOR U368 ( .A(x[23]), .B(y[23]), .Z(n200) );
  XOR U369 ( .A(x[21]), .B(y[21]), .Z(n199) );
  XNOR U370 ( .A(n200), .B(n199), .Z(n201) );
  XOR U371 ( .A(x[25]), .B(y[25]), .Z(n202) );
  XNOR U372 ( .A(n201), .B(n202), .Z(n237) );
  XOR U373 ( .A(n236), .B(n237), .Z(n147) );
  XNOR U374 ( .A(x[7]), .B(y[7]), .Z(n289) );
  XNOR U375 ( .A(x[5]), .B(y[5]), .Z(n287) );
  XOR U376 ( .A(x[3]), .B(y[3]), .Z(n286) );
  XNOR U377 ( .A(n287), .B(n286), .Z(n288) );
  XOR U378 ( .A(n289), .B(n288), .Z(n159) );
  XNOR U379 ( .A(x[4]), .B(y[4]), .Z(n266) );
  XNOR U380 ( .A(x[8]), .B(y[8]), .Z(n264) );
  XOR U381 ( .A(x[6]), .B(y[6]), .Z(n263) );
  XNOR U382 ( .A(n264), .B(n263), .Z(n265) );
  XOR U383 ( .A(n266), .B(n265), .Z(n156) );
  XNOR U384 ( .A(x[1]), .B(y[1]), .Z(n262) );
  XNOR U385 ( .A(x[2]), .B(y[2]), .Z(n260) );
  XOR U386 ( .A(x[0]), .B(y[0]), .Z(n259) );
  XNOR U387 ( .A(n260), .B(n259), .Z(n261) );
  XNOR U388 ( .A(n262), .B(n261), .Z(n157) );
  XNOR U389 ( .A(n156), .B(n157), .Z(n158) );
  XNOR U390 ( .A(n159), .B(n158), .Z(n148) );
  XNOR U391 ( .A(n147), .B(n148), .Z(n149) );
  XOR U392 ( .A(n150), .B(n149), .Z(n312) );
  XOR U393 ( .A(n313), .B(n312), .Z(o[0]) );
  OR U394 ( .A(n114), .B(n113), .Z(n118) );
  OR U395 ( .A(n116), .B(n115), .Z(n117) );
  NAND U396 ( .A(n118), .B(n117), .Z(n367) );
  XOR U397 ( .A(n365), .B(n366), .Z(n368) );
  XOR U398 ( .A(n367), .B(n368), .Z(n346) );
  OR U399 ( .A(n132), .B(n131), .Z(n136) );
  OR U400 ( .A(n134), .B(n133), .Z(n135) );
  NAND U401 ( .A(n136), .B(n135), .Z(n359) );
  XOR U402 ( .A(n359), .B(n360), .Z(n141) );
  XNOR U403 ( .A(n361), .B(n141), .Z(n344) );
  XOR U404 ( .A(n344), .B(n345), .Z(n146) );
  XOR U405 ( .A(n346), .B(n146), .Z(n383) );
  NANDN U406 ( .A(n148), .B(n147), .Z(n152) );
  NAND U407 ( .A(n150), .B(n149), .Z(n151) );
  NAND U408 ( .A(n152), .B(n151), .Z(n380) );
  XNOR U409 ( .A(n380), .B(n381), .Z(n382) );
  XOR U410 ( .A(n383), .B(n382), .Z(n407) );
  NANDN U411 ( .A(n157), .B(n156), .Z(n161) );
  NAND U412 ( .A(n159), .B(n158), .Z(n160) );
  AND U413 ( .A(n161), .B(n160), .Z(n403) );
  OR U414 ( .A(n163), .B(n162), .Z(n167) );
  OR U415 ( .A(n165), .B(n164), .Z(n166) );
  NAND U416 ( .A(n167), .B(n166), .Z(n339) );
  OR U417 ( .A(n169), .B(n168), .Z(n173) );
  OR U418 ( .A(n171), .B(n170), .Z(n172) );
  NAND U419 ( .A(n173), .B(n172), .Z(n338) );
  XNOR U420 ( .A(n339), .B(n338), .Z(n341) );
  OR U421 ( .A(n175), .B(n174), .Z(n179) );
  OR U422 ( .A(n177), .B(n176), .Z(n178) );
  NAND U423 ( .A(n179), .B(n178), .Z(n340) );
  XNOR U424 ( .A(n341), .B(n340), .Z(n389) );
  NANDN U425 ( .A(n180), .B(n181), .Z(n186) );
  NOR U426 ( .A(n182), .B(n181), .Z(n184) );
  NANDN U427 ( .A(n184), .B(n183), .Z(n185) );
  NAND U428 ( .A(n186), .B(n185), .Z(n386) );
  OR U429 ( .A(n188), .B(n187), .Z(n192) );
  OR U430 ( .A(n190), .B(n189), .Z(n191) );
  NAND U431 ( .A(n192), .B(n191), .Z(n358) );
  OR U432 ( .A(n194), .B(n193), .Z(n198) );
  OR U433 ( .A(n196), .B(n195), .Z(n197) );
  AND U434 ( .A(n198), .B(n197), .Z(n357) );
  XOR U435 ( .A(n386), .B(n387), .Z(n388) );
  XOR U436 ( .A(n389), .B(n388), .Z(n404) );
  OR U437 ( .A(n204), .B(n203), .Z(n208) );
  NANDN U438 ( .A(n206), .B(n205), .Z(n207) );
  AND U439 ( .A(n208), .B(n207), .Z(n331) );
  IV U440 ( .A(n209), .Z(n210) );
  OR U441 ( .A(n211), .B(n210), .Z(n215) );
  NANDN U442 ( .A(n213), .B(n212), .Z(n214) );
  AND U443 ( .A(n215), .B(n214), .Z(n332) );
  XOR U444 ( .A(n331), .B(n332), .Z(n333) );
  XOR U445 ( .A(n334), .B(n333), .Z(n392) );
  XNOR U446 ( .A(n337), .B(n335), .Z(n231) );
  XNOR U447 ( .A(n336), .B(n231), .Z(n394) );
  XNOR U448 ( .A(n393), .B(n394), .Z(n232) );
  XOR U449 ( .A(n392), .B(n232), .Z(n402) );
  XNOR U450 ( .A(n404), .B(n402), .Z(n233) );
  XNOR U451 ( .A(n403), .B(n233), .Z(n318) );
  OR U452 ( .A(n242), .B(n241), .Z(n246) );
  NANDN U453 ( .A(n244), .B(n243), .Z(n245) );
  AND U454 ( .A(n246), .B(n245), .Z(n326) );
  XNOR U455 ( .A(n325), .B(n326), .Z(n327) );
  XNOR U456 ( .A(n328), .B(n327), .Z(n322) );
  XOR U457 ( .A(n395), .B(n396), .Z(n398) );
  NAND U458 ( .A(n254), .B(oglobal[0]), .Z(n258) );
  OR U459 ( .A(n256), .B(n255), .Z(n257) );
  AND U460 ( .A(n258), .B(n257), .Z(n350) );
  XNOR U461 ( .A(n348), .B(n349), .Z(n351) );
  XNOR U462 ( .A(n350), .B(n351), .Z(n397) );
  XOR U463 ( .A(n398), .B(n397), .Z(n319) );
  OR U464 ( .A(n276), .B(n275), .Z(n280) );
  NANDN U465 ( .A(n278), .B(n277), .Z(n279) );
  NAND U466 ( .A(n280), .B(n279), .Z(n362) );
  XOR U467 ( .A(n362), .B(n363), .Z(n285) );
  XNOR U468 ( .A(n364), .B(n285), .Z(n373) );
  IV U469 ( .A(n373), .Z(n372) );
  OR U470 ( .A(n291), .B(n290), .Z(n295) );
  NANDN U471 ( .A(n293), .B(n292), .Z(n294) );
  NAND U472 ( .A(n295), .B(n294), .Z(n354) );
  XOR U473 ( .A(n354), .B(n355), .Z(n300) );
  XOR U474 ( .A(n356), .B(n300), .Z(n374) );
  XNOR U475 ( .A(n372), .B(n374), .Z(n301) );
  XOR U476 ( .A(n375), .B(n301), .Z(n320) );
  XOR U477 ( .A(n319), .B(n320), .Z(n321) );
  XOR U478 ( .A(n322), .B(n321), .Z(n317) );
  NANDN U479 ( .A(n302), .B(n303), .Z(n308) );
  NOR U480 ( .A(n304), .B(n303), .Z(n305) );
  OR U481 ( .A(n306), .B(n305), .Z(n307) );
  NAND U482 ( .A(n308), .B(n307), .Z(n316) );
  XOR U483 ( .A(n317), .B(n316), .Z(n309) );
  XNOR U484 ( .A(n318), .B(n309), .Z(n406) );
  XOR U485 ( .A(n407), .B(n406), .Z(n409) );
  NANDN U486 ( .A(n311), .B(n310), .Z(n315) );
  OR U487 ( .A(n313), .B(n312), .Z(n314) );
  AND U488 ( .A(n315), .B(n314), .Z(n408) );
  XOR U489 ( .A(n409), .B(n408), .Z(o[1]) );
  NANDN U490 ( .A(n320), .B(n319), .Z(n324) );
  OR U491 ( .A(n322), .B(n321), .Z(n323) );
  NAND U492 ( .A(n324), .B(n323), .Z(n413) );
  NANDN U493 ( .A(n326), .B(n325), .Z(n330) );
  NAND U494 ( .A(n328), .B(n327), .Z(n329) );
  NAND U495 ( .A(n330), .B(n329), .Z(n445) );
  OR U496 ( .A(n339), .B(n338), .Z(n343) );
  OR U497 ( .A(n341), .B(n340), .Z(n342) );
  NAND U498 ( .A(n343), .B(n342), .Z(n424) );
  XOR U499 ( .A(n425), .B(n424), .Z(n426) );
  XOR U500 ( .A(n427), .B(n426), .Z(n444) );
  XOR U501 ( .A(n444), .B(n443), .Z(n347) );
  XOR U502 ( .A(n445), .B(n347), .Z(n434) );
  OR U503 ( .A(n349), .B(n348), .Z(n353) );
  OR U504 ( .A(n351), .B(n350), .Z(n352) );
  AND U505 ( .A(n353), .B(n352), .Z(n439) );
  XNOR U506 ( .A(n438), .B(oglobal[2]), .Z(n440) );
  XNOR U507 ( .A(n439), .B(n440), .Z(n416) );
  XNOR U508 ( .A(n416), .B(n415), .Z(n417) );
  NAND U509 ( .A(n366), .B(n365), .Z(n370) );
  NAND U510 ( .A(n368), .B(n367), .Z(n369) );
  AND U511 ( .A(n370), .B(n369), .Z(n435) );
  XNOR U512 ( .A(n436), .B(n435), .Z(n371) );
  XNOR U513 ( .A(n437), .B(n371), .Z(n418) );
  XNOR U514 ( .A(n417), .B(n418), .Z(n432) );
  OR U515 ( .A(n374), .B(n372), .Z(n378) );
  ANDN U516 ( .B(n374), .A(n373), .Z(n376) );
  NANDN U517 ( .A(n376), .B(n375), .Z(n377) );
  NAND U518 ( .A(n378), .B(n377), .Z(n431) );
  XNOR U519 ( .A(n432), .B(n431), .Z(n433) );
  XOR U520 ( .A(n434), .B(n433), .Z(n414) );
  XOR U521 ( .A(n413), .B(n414), .Z(n379) );
  XNOR U522 ( .A(n412), .B(n379), .Z(n451) );
  NANDN U523 ( .A(n381), .B(n380), .Z(n385) );
  NAND U524 ( .A(n383), .B(n382), .Z(n384) );
  AND U525 ( .A(n385), .B(n384), .Z(n448) );
  NAND U526 ( .A(n387), .B(n386), .Z(n391) );
  NAND U527 ( .A(n389), .B(n388), .Z(n390) );
  AND U528 ( .A(n391), .B(n390), .Z(n423) );
  NANDN U529 ( .A(n396), .B(n395), .Z(n400) );
  OR U530 ( .A(n398), .B(n397), .Z(n399) );
  AND U531 ( .A(n400), .B(n399), .Z(n422) );
  XOR U532 ( .A(n421), .B(n422), .Z(n401) );
  XNOR U533 ( .A(n423), .B(n401), .Z(n447) );
  XOR U534 ( .A(n447), .B(n446), .Z(n405) );
  XOR U535 ( .A(n448), .B(n405), .Z(n450) );
  XOR U536 ( .A(n451), .B(n450), .Z(n453) );
  NANDN U537 ( .A(n407), .B(n406), .Z(n411) );
  OR U538 ( .A(n409), .B(n408), .Z(n410) );
  AND U539 ( .A(n411), .B(n410), .Z(n452) );
  XOR U540 ( .A(n453), .B(n452), .Z(o[2]) );
  NANDN U541 ( .A(n416), .B(n415), .Z(n420) );
  NAND U542 ( .A(n418), .B(n417), .Z(n419) );
  NAND U543 ( .A(n420), .B(n419), .Z(n478) );
  OR U544 ( .A(n425), .B(n424), .Z(n429) );
  NAND U545 ( .A(n427), .B(n426), .Z(n428) );
  AND U546 ( .A(n429), .B(n428), .Z(n477) );
  XOR U547 ( .A(n476), .B(n477), .Z(n430) );
  XNOR U548 ( .A(n478), .B(n430), .Z(n456) );
  XNOR U549 ( .A(n471), .B(oglobal[3]), .Z(n473) );
  NAND U550 ( .A(n438), .B(oglobal[2]), .Z(n442) );
  OR U551 ( .A(n440), .B(n439), .Z(n441) );
  NAND U552 ( .A(n442), .B(n441), .Z(n472) );
  XOR U553 ( .A(n473), .B(n472), .Z(n466) );
  XNOR U554 ( .A(n466), .B(n465), .Z(n467) );
  XNOR U555 ( .A(n468), .B(n467), .Z(n458) );
  XOR U556 ( .A(n458), .B(n457), .Z(n449) );
  XNOR U557 ( .A(n456), .B(n449), .Z(n460) );
  XOR U558 ( .A(n459), .B(n460), .Z(n461) );
  NANDN U559 ( .A(n451), .B(n450), .Z(n455) );
  OR U560 ( .A(n453), .B(n452), .Z(n454) );
  AND U561 ( .A(n455), .B(n454), .Z(n462) );
  XNOR U562 ( .A(n461), .B(n462), .Z(o[3]) );
  NAND U563 ( .A(n460), .B(n459), .Z(n464) );
  NANDN U564 ( .A(n462), .B(n461), .Z(n463) );
  AND U565 ( .A(n464), .B(n463), .Z(n485) );
  XNOR U566 ( .A(n484), .B(n485), .Z(n486) );
  NANDN U567 ( .A(n466), .B(n465), .Z(n470) );
  NAND U568 ( .A(n468), .B(n467), .Z(n469) );
  NAND U569 ( .A(n470), .B(n469), .Z(n483) );
  NAND U570 ( .A(oglobal[3]), .B(n471), .Z(n475) );
  NANDN U571 ( .A(n473), .B(n472), .Z(n474) );
  AND U572 ( .A(n475), .B(n474), .Z(n480) );
  XNOR U573 ( .A(oglobal[4]), .B(n480), .Z(n482) );
  XOR U574 ( .A(n482), .B(n481), .Z(n479) );
  XOR U575 ( .A(n483), .B(n479), .Z(n487) );
  XOR U576 ( .A(n486), .B(n487), .Z(o[4]) );
  ANDN U577 ( .B(oglobal[4]), .A(n480), .Z(n490) );
  XOR U578 ( .A(oglobal[5]), .B(n490), .Z(n493) );
  XOR U579 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U580 ( .A(n485), .B(n484), .Z(n489) );
  NAND U581 ( .A(n487), .B(n486), .Z(n488) );
  AND U582 ( .A(n489), .B(n488), .Z(n491) );
  XOR U583 ( .A(n492), .B(n491), .Z(o[5]) );
  AND U584 ( .A(n490), .B(oglobal[5]), .Z(n496) );
  OR U585 ( .A(n492), .B(n491), .Z(n495) );
  ANDN U586 ( .B(n496), .A(n495), .Z(n500) );
  OR U587 ( .A(n500), .B(n498), .Z(n497) );
  XNOR U588 ( .A(oglobal[6]), .B(n497), .Z(o[6]) );
  NANDN U589 ( .A(n498), .B(oglobal[6]), .Z(n499) );
  NANDN U590 ( .A(n500), .B(n499), .Z(n501) );
  XOR U591 ( .A(oglobal[7]), .B(n501), .Z(o[7]) );
endmodule

