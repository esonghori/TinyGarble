
module mult_N1024_CC256 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [3:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2043]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2043]) );
  DFF \sreg_reg[2042]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2042]) );
  DFF \sreg_reg[2041]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2041]) );
  DFF \sreg_reg[2040]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2040]) );
  DFF \sreg_reg[2039]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U7 ( .A(n3246), .B(n3245), .Z(n1) );
  NANDN U8 ( .A(n3247), .B(n3248), .Z(n2) );
  NAND U9 ( .A(n1), .B(n2), .Z(n3256) );
  NANDN U10 ( .A(n7788), .B(n7787), .Z(n3) );
  NANDN U11 ( .A(n7789), .B(n7790), .Z(n4) );
  NAND U12 ( .A(n3), .B(n4), .Z(n7798) );
  NAND U13 ( .A(n8083), .B(n8081), .Z(n5) );
  XOR U14 ( .A(n8081), .B(n8083), .Z(n6) );
  NANDN U15 ( .A(n8082), .B(n6), .Z(n7) );
  NAND U16 ( .A(n5), .B(n7), .Z(n8104) );
  NANDN U17 ( .A(n14064), .B(n14063), .Z(n8) );
  NANDN U18 ( .A(n14065), .B(n14066), .Z(n9) );
  NAND U19 ( .A(n8), .B(n9), .Z(n14091) );
  NANDN U20 ( .A(n16856), .B(n16855), .Z(n10) );
  NANDN U21 ( .A(n16857), .B(n16858), .Z(n11) );
  NAND U22 ( .A(n10), .B(n11), .Z(n16866) );
  NANDN U23 ( .A(n19305), .B(n19306), .Z(n12) );
  NANDN U24 ( .A(n19304), .B(n19303), .Z(n13) );
  AND U25 ( .A(n12), .B(n13), .Z(n19314) );
  NANDN U26 ( .A(n23136), .B(n23135), .Z(n14) );
  NANDN U27 ( .A(n23137), .B(n23138), .Z(n15) );
  NAND U28 ( .A(n14), .B(n15), .Z(n23163) );
  NAND U29 ( .A(n16788), .B(n16786), .Z(n16) );
  XOR U30 ( .A(n16786), .B(n16788), .Z(n17) );
  NANDN U31 ( .A(n16787), .B(n17), .Z(n18) );
  NAND U32 ( .A(n16), .B(n18), .Z(n16807) );
  NAND U33 ( .A(n2492), .B(sreg[1053]), .Z(n19) );
  XOR U34 ( .A(sreg[1053]), .B(n2492), .Z(n20) );
  NAND U35 ( .A(n20), .B(n2491), .Z(n21) );
  NAND U36 ( .A(n19), .B(n21), .Z(n2512) );
  NAND U37 ( .A(sreg[1099]), .B(n3489), .Z(n22) );
  XOR U38 ( .A(n3489), .B(sreg[1099]), .Z(n23) );
  NANDN U39 ( .A(n3490), .B(n23), .Z(n24) );
  NAND U40 ( .A(n22), .B(n24), .Z(n3510) );
  NAND U41 ( .A(n3641), .B(sreg[1106]), .Z(n25) );
  XOR U42 ( .A(sreg[1106]), .B(n3641), .Z(n26) );
  NAND U43 ( .A(n26), .B(n3640), .Z(n27) );
  NAND U44 ( .A(n25), .B(n27), .Z(n3661) );
  NAND U45 ( .A(sreg[1117]), .B(n3881), .Z(n28) );
  XOR U46 ( .A(n3881), .B(sreg[1117]), .Z(n29) );
  NANDN U47 ( .A(n3882), .B(n29), .Z(n30) );
  NAND U48 ( .A(n28), .B(n30), .Z(n3902) );
  NAND U49 ( .A(sreg[1140]), .B(n4382), .Z(n31) );
  XOR U50 ( .A(n4382), .B(sreg[1140]), .Z(n32) );
  NANDN U51 ( .A(n4383), .B(n32), .Z(n33) );
  NAND U52 ( .A(n31), .B(n33), .Z(n4403) );
  XOR U53 ( .A(n5600), .B(n5599), .Z(n34) );
  NAND U54 ( .A(n34), .B(sreg[1195]), .Z(n35) );
  NAND U55 ( .A(n5600), .B(n5599), .Z(n36) );
  AND U56 ( .A(n35), .B(n36), .Z(n5620) );
  NAND U57 ( .A(sreg[1213]), .B(n5989), .Z(n37) );
  XOR U58 ( .A(n5989), .B(sreg[1213]), .Z(n38) );
  NANDN U59 ( .A(n5990), .B(n38), .Z(n39) );
  NAND U60 ( .A(n37), .B(n39), .Z(n6010) );
  NAND U61 ( .A(sreg[1247]), .B(n6733), .Z(n40) );
  XOR U62 ( .A(n6733), .B(sreg[1247]), .Z(n41) );
  NANDN U63 ( .A(n6734), .B(n41), .Z(n42) );
  NAND U64 ( .A(n40), .B(n42), .Z(n6754) );
  NAND U65 ( .A(n7145), .B(sreg[1266]), .Z(n43) );
  XOR U66 ( .A(sreg[1266]), .B(n7145), .Z(n44) );
  NANDN U67 ( .A(n7144), .B(n44), .Z(n45) );
  NAND U68 ( .A(n43), .B(n45), .Z(n7165) );
  NAND U69 ( .A(sreg[1282]), .B(n7494), .Z(n46) );
  XOR U70 ( .A(n7494), .B(sreg[1282]), .Z(n47) );
  NANDN U71 ( .A(n7495), .B(n47), .Z(n48) );
  NAND U72 ( .A(n46), .B(n48), .Z(n7515) );
  NAND U73 ( .A(sreg[1315]), .B(n8199), .Z(n49) );
  XOR U74 ( .A(n8199), .B(sreg[1315]), .Z(n50) );
  NANDN U75 ( .A(n8200), .B(n50), .Z(n51) );
  NAND U76 ( .A(n49), .B(n51), .Z(n8220) );
  NAND U77 ( .A(sreg[1330]), .B(n8518), .Z(n52) );
  XOR U78 ( .A(n8518), .B(sreg[1330]), .Z(n53) );
  NANDN U79 ( .A(n8519), .B(n53), .Z(n54) );
  NAND U80 ( .A(n52), .B(n54), .Z(n8539) );
  NAND U81 ( .A(n8603), .B(n8602), .Z(n55) );
  XOR U82 ( .A(n8602), .B(n8603), .Z(n56) );
  NAND U83 ( .A(n56), .B(sreg[1334]), .Z(n57) );
  NAND U84 ( .A(n55), .B(n57), .Z(n8623) );
  NAND U85 ( .A(sreg[1373]), .B(n9459), .Z(n58) );
  XOR U86 ( .A(n9459), .B(sreg[1373]), .Z(n59) );
  NANDN U87 ( .A(n9460), .B(n59), .Z(n60) );
  NAND U88 ( .A(n58), .B(n60), .Z(n9480) );
  XOR U89 ( .A(n9605), .B(n9604), .Z(n61) );
  NANDN U90 ( .A(sreg[1380]), .B(n61), .Z(n62) );
  NAND U91 ( .A(n9605), .B(n9604), .Z(n63) );
  AND U92 ( .A(n62), .B(n63), .Z(n9625) );
  NAND U93 ( .A(n11550), .B(sreg[1469]), .Z(n64) );
  XOR U94 ( .A(sreg[1469]), .B(n11550), .Z(n65) );
  NAND U95 ( .A(n65), .B(n11549), .Z(n66) );
  NAND U96 ( .A(n64), .B(n66), .Z(n11570) );
  NAND U97 ( .A(n11988), .B(n11987), .Z(n67) );
  XOR U98 ( .A(n11987), .B(n11988), .Z(n68) );
  NAND U99 ( .A(n68), .B(sreg[1489]), .Z(n69) );
  NAND U100 ( .A(n67), .B(n69), .Z(n12008) );
  NAND U101 ( .A(sreg[1655]), .B(n15629), .Z(n70) );
  XOR U102 ( .A(n15629), .B(sreg[1655]), .Z(n71) );
  NANDN U103 ( .A(n15630), .B(n71), .Z(n72) );
  NAND U104 ( .A(n70), .B(n72), .Z(n15650) );
  NAND U105 ( .A(sreg[1684]), .B(n16256), .Z(n73) );
  XOR U106 ( .A(n16256), .B(sreg[1684]), .Z(n74) );
  NANDN U107 ( .A(n16257), .B(n74), .Z(n75) );
  NAND U108 ( .A(n73), .B(n75), .Z(n16277) );
  XOR U109 ( .A(n17234), .B(n17233), .Z(n76) );
  NAND U110 ( .A(n76), .B(sreg[1729]), .Z(n77) );
  NAND U111 ( .A(n17234), .B(n17233), .Z(n78) );
  AND U112 ( .A(n77), .B(n78), .Z(n17254) );
  XOR U113 ( .A(n17362), .B(n17361), .Z(n79) );
  NAND U114 ( .A(n79), .B(sreg[1735]), .Z(n80) );
  NAND U115 ( .A(n17362), .B(n17361), .Z(n81) );
  AND U116 ( .A(n80), .B(n81), .Z(n17382) );
  NAND U117 ( .A(sreg[1782]), .B(n18402), .Z(n82) );
  XOR U118 ( .A(n18402), .B(sreg[1782]), .Z(n83) );
  NANDN U119 ( .A(n18403), .B(n83), .Z(n84) );
  NAND U120 ( .A(n82), .B(n84), .Z(n18423) );
  NAND U121 ( .A(sreg[1789]), .B(n18553), .Z(n85) );
  XOR U122 ( .A(n18553), .B(sreg[1789]), .Z(n86) );
  NANDN U123 ( .A(n18554), .B(n86), .Z(n87) );
  NAND U124 ( .A(n85), .B(n87), .Z(n18574) );
  NAND U125 ( .A(sreg[1809]), .B(n18989), .Z(n88) );
  XOR U126 ( .A(n18989), .B(sreg[1809]), .Z(n89) );
  NANDN U127 ( .A(n18990), .B(n89), .Z(n90) );
  NAND U128 ( .A(n88), .B(n90), .Z(n19010) );
  NAND U129 ( .A(sreg[1832]), .B(n19482), .Z(n91) );
  XOR U130 ( .A(n19482), .B(sreg[1832]), .Z(n92) );
  NANDN U131 ( .A(n19483), .B(n92), .Z(n93) );
  NAND U132 ( .A(n91), .B(n93), .Z(n19503) );
  XOR U133 ( .A(n21526), .B(sreg[1926]), .Z(n94) );
  NANDN U134 ( .A(n21527), .B(n94), .Z(n95) );
  NAND U135 ( .A(n21526), .B(sreg[1926]), .Z(n96) );
  AND U136 ( .A(n95), .B(n96), .Z(n21547) );
  NAND U137 ( .A(n22914), .B(sreg[1989]), .Z(n97) );
  XOR U138 ( .A(sreg[1989]), .B(n22914), .Z(n98) );
  NAND U139 ( .A(n98), .B(n22913), .Z(n99) );
  NAND U140 ( .A(n97), .B(n99), .Z(n22934) );
  NAND U141 ( .A(b[1]), .B(a[1021]), .Z(n24059) );
  OR U142 ( .A(n24079), .B(n24039), .Z(n100) );
  NANDN U143 ( .A(n24041), .B(n24040), .Z(n101) );
  AND U144 ( .A(n100), .B(n101), .Z(n24067) );
  NAND U145 ( .A(n2541), .B(n2540), .Z(n102) );
  XOR U146 ( .A(n2540), .B(n2541), .Z(n103) );
  NAND U147 ( .A(n103), .B(n2539), .Z(n104) );
  NAND U148 ( .A(n102), .B(n104), .Z(n2567) );
  NAND U149 ( .A(n3930), .B(n3929), .Z(n105) );
  XOR U150 ( .A(n3929), .B(n3930), .Z(n106) );
  NANDN U151 ( .A(n3931), .B(n106), .Z(n107) );
  NAND U152 ( .A(n105), .B(n107), .Z(n3944) );
  NAND U153 ( .A(n5649), .B(n5647), .Z(n108) );
  XOR U154 ( .A(n5647), .B(n5649), .Z(n109) );
  NANDN U155 ( .A(n5648), .B(n109), .Z(n110) );
  NAND U156 ( .A(n108), .B(n110), .Z(n5682) );
  NANDN U157 ( .A(n5717), .B(n5716), .Z(n111) );
  NANDN U158 ( .A(n5718), .B(n5719), .Z(n112) );
  NAND U159 ( .A(n111), .B(n112), .Z(n5729) );
  NAND U160 ( .A(n6636), .B(n6635), .Z(n113) );
  XOR U161 ( .A(n6635), .B(n6636), .Z(n114) );
  NAND U162 ( .A(n114), .B(n6634), .Z(n115) );
  NAND U163 ( .A(n113), .B(n115), .Z(n6649) );
  NANDN U164 ( .A(n7093), .B(n7092), .Z(n116) );
  NANDN U165 ( .A(n7094), .B(n7095), .Z(n117) );
  NAND U166 ( .A(n116), .B(n117), .Z(n7117) );
  NAND U167 ( .A(n8124), .B(n8123), .Z(n118) );
  XOR U168 ( .A(n8123), .B(n8124), .Z(n119) );
  NANDN U169 ( .A(n8125), .B(n119), .Z(n120) );
  NAND U170 ( .A(n118), .B(n120), .Z(n8151) );
  NANDN U171 ( .A(n9517), .B(n9516), .Z(n121) );
  NANDN U172 ( .A(n9518), .B(n9519), .Z(n122) );
  NAND U173 ( .A(n121), .B(n122), .Z(n9521) );
  NANDN U174 ( .A(n9944), .B(n9943), .Z(n123) );
  NANDN U175 ( .A(n9945), .B(n9946), .Z(n124) );
  NAND U176 ( .A(n123), .B(n124), .Z(n9956) );
  NANDN U177 ( .A(n10198), .B(n10197), .Z(n125) );
  NANDN U178 ( .A(n10199), .B(n10200), .Z(n126) );
  NAND U179 ( .A(n125), .B(n126), .Z(n10212) );
  NANDN U180 ( .A(n13002), .B(n13001), .Z(n127) );
  NANDN U181 ( .A(n13003), .B(n13004), .Z(n128) );
  NAND U182 ( .A(n127), .B(n128), .Z(n13016) );
  NAND U183 ( .A(n16035), .B(n16034), .Z(n129) );
  XOR U184 ( .A(n16034), .B(n16035), .Z(n130) );
  NAND U185 ( .A(n130), .B(n16033), .Z(n131) );
  NAND U186 ( .A(n129), .B(n131), .Z(n16060) );
  NAND U187 ( .A(n16158), .B(n16157), .Z(n132) );
  XOR U188 ( .A(n16157), .B(n16158), .Z(n133) );
  NANDN U189 ( .A(n16159), .B(n133), .Z(n134) );
  NAND U190 ( .A(n132), .B(n134), .Z(n16185) );
  XOR U191 ( .A(n19238), .B(n19237), .Z(n135) );
  NANDN U192 ( .A(n19236), .B(n135), .Z(n136) );
  NAND U193 ( .A(n19238), .B(n19237), .Z(n137) );
  AND U194 ( .A(n136), .B(n137), .Z(n19254) );
  NANDN U195 ( .A(n19323), .B(n19322), .Z(n138) );
  NANDN U196 ( .A(n19324), .B(n19325), .Z(n139) );
  NAND U197 ( .A(n138), .B(n139), .Z(n19335) );
  NAND U198 ( .A(n19295), .B(n19294), .Z(n140) );
  XOR U199 ( .A(n19294), .B(n19295), .Z(n141) );
  NANDN U200 ( .A(n19296), .B(n141), .Z(n142) );
  NAND U201 ( .A(n140), .B(n142), .Z(n19315) );
  NAND U202 ( .A(n20564), .B(n20563), .Z(n143) );
  XOR U203 ( .A(n20563), .B(n20564), .Z(n144) );
  NANDN U204 ( .A(n20565), .B(n144), .Z(n145) );
  NAND U205 ( .A(n143), .B(n145), .Z(n20578) );
  NAND U206 ( .A(n20689), .B(n20688), .Z(n146) );
  XOR U207 ( .A(n20688), .B(n20689), .Z(n147) );
  NAND U208 ( .A(n147), .B(n20687), .Z(n148) );
  NAND U209 ( .A(n146), .B(n148), .Z(n20715) );
  NAND U210 ( .A(n3176), .B(n3174), .Z(n149) );
  XOR U211 ( .A(n3174), .B(n3176), .Z(n150) );
  NANDN U212 ( .A(n3175), .B(n150), .Z(n151) );
  NAND U213 ( .A(n149), .B(n151), .Z(n3197) );
  XOR U214 ( .A(n8421), .B(n8420), .Z(n152) );
  NANDN U215 ( .A(n8419), .B(n152), .Z(n153) );
  NAND U216 ( .A(n8421), .B(n8420), .Z(n154) );
  AND U217 ( .A(n153), .B(n154), .Z(n8442) );
  NAND U218 ( .A(n10064), .B(n10063), .Z(n155) );
  XOR U219 ( .A(n10063), .B(n10064), .Z(n156) );
  NANDN U220 ( .A(n10065), .B(n156), .Z(n157) );
  NAND U221 ( .A(n155), .B(n157), .Z(n10083) );
  NAND U222 ( .A(n12294), .B(n12293), .Z(n158) );
  XOR U223 ( .A(n12293), .B(n12294), .Z(n159) );
  NANDN U224 ( .A(n12295), .B(n159), .Z(n160) );
  NAND U225 ( .A(n158), .B(n160), .Z(n12313) );
  NAND U226 ( .A(n14062), .B(n14061), .Z(n161) );
  XOR U227 ( .A(n14061), .B(n14062), .Z(n162) );
  NAND U228 ( .A(n162), .B(n14060), .Z(n163) );
  NAND U229 ( .A(n161), .B(n163), .Z(n14094) );
  NAND U230 ( .A(n16847), .B(n16846), .Z(n164) );
  XOR U231 ( .A(n16846), .B(n16847), .Z(n165) );
  NANDN U232 ( .A(n16848), .B(n165), .Z(n166) );
  NAND U233 ( .A(n164), .B(n166), .Z(n16867) );
  NAND U234 ( .A(n23133), .B(n23132), .Z(n167) );
  XOR U235 ( .A(n23132), .B(n23133), .Z(n168) );
  NANDN U236 ( .A(n23134), .B(n168), .Z(n169) );
  NAND U237 ( .A(n167), .B(n169), .Z(n23166) );
  XOR U238 ( .A(n1880), .B(sreg[1025]), .Z(n170) );
  NANDN U239 ( .A(n1879), .B(n170), .Z(n171) );
  NAND U240 ( .A(n1880), .B(sreg[1025]), .Z(n172) );
  AND U241 ( .A(n171), .B(n172), .Z(n1900) );
  NAND U242 ( .A(sreg[1030]), .B(n1988), .Z(n173) );
  XOR U243 ( .A(n1988), .B(sreg[1030]), .Z(n174) );
  NANDN U244 ( .A(n1989), .B(n174), .Z(n175) );
  NAND U245 ( .A(n173), .B(n175), .Z(n1991) );
  NAND U246 ( .A(sreg[1048]), .B(n2384), .Z(n176) );
  XOR U247 ( .A(n2384), .B(sreg[1048]), .Z(n177) );
  NANDN U248 ( .A(n2385), .B(n177), .Z(n178) );
  NAND U249 ( .A(n176), .B(n178), .Z(n2387) );
  NAND U250 ( .A(sreg[1055]), .B(n2534), .Z(n179) );
  XOR U251 ( .A(n2534), .B(sreg[1055]), .Z(n180) );
  NANDN U252 ( .A(n2535), .B(n180), .Z(n181) );
  NAND U253 ( .A(n179), .B(n181), .Z(n2537) );
  XOR U254 ( .A(sreg[1060]), .B(n2620), .Z(n182) );
  NANDN U255 ( .A(n2621), .B(n182), .Z(n183) );
  NAND U256 ( .A(sreg[1060]), .B(n2620), .Z(n184) );
  AND U257 ( .A(n183), .B(n184), .Z(n2660) );
  XOR U258 ( .A(sreg[1079]), .B(n3041), .Z(n185) );
  NANDN U259 ( .A(n3042), .B(n185), .Z(n186) );
  NAND U260 ( .A(sreg[1079]), .B(n3041), .Z(n187) );
  AND U261 ( .A(n186), .B(n187), .Z(n3081) );
  NAND U262 ( .A(n3277), .B(n3276), .Z(n188) );
  XOR U263 ( .A(n3276), .B(n3277), .Z(n189) );
  NANDN U264 ( .A(sreg[1090]), .B(n189), .Z(n190) );
  NAND U265 ( .A(n188), .B(n190), .Z(n3298) );
  XOR U266 ( .A(n3404), .B(sreg[1095]), .Z(n191) );
  NANDN U267 ( .A(n3403), .B(n191), .Z(n192) );
  NAND U268 ( .A(n3404), .B(sreg[1095]), .Z(n193) );
  AND U269 ( .A(n192), .B(n193), .Z(n3406) );
  XOR U270 ( .A(n3532), .B(n3531), .Z(n194) );
  NAND U271 ( .A(n194), .B(sreg[1101]), .Z(n195) );
  NAND U272 ( .A(n3532), .B(n3531), .Z(n196) );
  AND U273 ( .A(n195), .B(n196), .Z(n3534) );
  NAND U274 ( .A(sreg[1107]), .B(n3661), .Z(n197) );
  XOR U275 ( .A(n3661), .B(sreg[1107]), .Z(n198) );
  NANDN U276 ( .A(n3662), .B(n198), .Z(n199) );
  NAND U277 ( .A(n197), .B(n199), .Z(n3682) );
  NAND U278 ( .A(sreg[1119]), .B(n3924), .Z(n200) );
  XOR U279 ( .A(n3924), .B(sreg[1119]), .Z(n201) );
  NANDN U280 ( .A(n3925), .B(n201), .Z(n202) );
  NAND U281 ( .A(n200), .B(n202), .Z(n3927) );
  XOR U282 ( .A(sreg[1127]), .B(n4077), .Z(n203) );
  NANDN U283 ( .A(n4078), .B(n203), .Z(n204) );
  NAND U284 ( .A(sreg[1127]), .B(n4077), .Z(n205) );
  AND U285 ( .A(n204), .B(n205), .Z(n4117) );
  NAND U286 ( .A(sreg[1139]), .B(n4361), .Z(n206) );
  XOR U287 ( .A(n4361), .B(sreg[1139]), .Z(n207) );
  NANDN U288 ( .A(n4362), .B(n207), .Z(n208) );
  NAND U289 ( .A(n206), .B(n208), .Z(n4382) );
  NAND U290 ( .A(n4428), .B(n4427), .Z(n209) );
  XOR U291 ( .A(n4427), .B(n4428), .Z(n210) );
  NAND U292 ( .A(n210), .B(sreg[1143]), .Z(n211) );
  NAND U293 ( .A(n209), .B(n211), .Z(n4448) );
  NAND U294 ( .A(n5029), .B(sreg[1170]), .Z(n212) );
  XOR U295 ( .A(sreg[1170]), .B(n5029), .Z(n213) );
  NANDN U296 ( .A(n5028), .B(n213), .Z(n214) );
  NAND U297 ( .A(n212), .B(n214), .Z(n5067) );
  XOR U298 ( .A(n5642), .B(sreg[1197]), .Z(n215) );
  NANDN U299 ( .A(n5643), .B(n215), .Z(n216) );
  NAND U300 ( .A(n5642), .B(sreg[1197]), .Z(n217) );
  AND U301 ( .A(n216), .B(n217), .Z(n5645) );
  NAND U302 ( .A(sreg[1215]), .B(n6031), .Z(n218) );
  XOR U303 ( .A(n6031), .B(sreg[1215]), .Z(n219) );
  NANDN U304 ( .A(n6032), .B(n219), .Z(n220) );
  NAND U305 ( .A(n218), .B(n220), .Z(n6034) );
  XOR U306 ( .A(sreg[1222]), .B(n6166), .Z(n221) );
  NANDN U307 ( .A(n6167), .B(n221), .Z(n222) );
  NAND U308 ( .A(sreg[1222]), .B(n6166), .Z(n223) );
  AND U309 ( .A(n222), .B(n223), .Z(n6206) );
  XOR U310 ( .A(n6776), .B(n6775), .Z(n224) );
  NAND U311 ( .A(n224), .B(sreg[1249]), .Z(n225) );
  NAND U312 ( .A(n6776), .B(n6775), .Z(n226) );
  AND U313 ( .A(n225), .B(n226), .Z(n6778) );
  XOR U314 ( .A(sreg[1264]), .B(n7102), .Z(n227) );
  NANDN U315 ( .A(n7103), .B(n227), .Z(n228) );
  NAND U316 ( .A(sreg[1264]), .B(n7102), .Z(n229) );
  AND U317 ( .A(n228), .B(n229), .Z(n7124) );
  NAND U318 ( .A(sreg[1268]), .B(n7186), .Z(n230) );
  XOR U319 ( .A(n7186), .B(sreg[1268]), .Z(n231) );
  NANDN U320 ( .A(n7187), .B(n231), .Z(n232) );
  NAND U321 ( .A(n230), .B(n232), .Z(n7189) );
  NAND U322 ( .A(sreg[1281]), .B(n7473), .Z(n233) );
  XOR U323 ( .A(n7473), .B(sreg[1281]), .Z(n234) );
  NANDN U324 ( .A(n7474), .B(n234), .Z(n235) );
  NAND U325 ( .A(n233), .B(n235), .Z(n7494) );
  NAND U326 ( .A(n7540), .B(n7539), .Z(n236) );
  XOR U327 ( .A(n7539), .B(n7540), .Z(n237) );
  NAND U328 ( .A(n237), .B(sreg[1285]), .Z(n238) );
  NAND U329 ( .A(n236), .B(n238), .Z(n7578) );
  XOR U330 ( .A(n7667), .B(sreg[1290]), .Z(n239) );
  NANDN U331 ( .A(n7666), .B(n239), .Z(n240) );
  NAND U332 ( .A(n7667), .B(sreg[1290]), .Z(n241) );
  AND U333 ( .A(n240), .B(n241), .Z(n7687) );
  NAND U334 ( .A(sreg[1297]), .B(n7815), .Z(n242) );
  XOR U335 ( .A(n7815), .B(sreg[1297]), .Z(n243) );
  NANDN U336 ( .A(n7816), .B(n243), .Z(n244) );
  NAND U337 ( .A(n242), .B(n244), .Z(n7818) );
  NAND U338 ( .A(n7948), .B(sreg[1303]), .Z(n245) );
  XOR U339 ( .A(sreg[1303]), .B(n7948), .Z(n246) );
  NANDN U340 ( .A(n7947), .B(n246), .Z(n247) );
  NAND U341 ( .A(n245), .B(n247), .Z(n7968) );
  XOR U342 ( .A(n8077), .B(n8076), .Z(n248) );
  NAND U343 ( .A(n248), .B(sreg[1309]), .Z(n249) );
  NAND U344 ( .A(n8077), .B(n8076), .Z(n250) );
  AND U345 ( .A(n249), .B(n250), .Z(n8079) );
  NAND U346 ( .A(n8220), .B(sreg[1316]), .Z(n251) );
  XOR U347 ( .A(sreg[1316]), .B(n8220), .Z(n252) );
  NANDN U348 ( .A(n8221), .B(n252), .Z(n253) );
  NAND U349 ( .A(n251), .B(n253), .Z(n8241) );
  NAND U350 ( .A(n8307), .B(sreg[1320]), .Z(n254) );
  XOR U351 ( .A(sreg[1320]), .B(n8307), .Z(n255) );
  NAND U352 ( .A(n255), .B(n8306), .Z(n256) );
  NAND U353 ( .A(n254), .B(n256), .Z(n8309) );
  NAND U354 ( .A(n8417), .B(n8416), .Z(n257) );
  XOR U355 ( .A(n8416), .B(n8417), .Z(n258) );
  NAND U356 ( .A(n258), .B(sreg[1325]), .Z(n259) );
  NAND U357 ( .A(n257), .B(n259), .Z(n8434) );
  XOR U358 ( .A(sreg[1331]), .B(n8539), .Z(n260) );
  NANDN U359 ( .A(n8540), .B(n260), .Z(n261) );
  NAND U360 ( .A(sreg[1331]), .B(n8539), .Z(n262) );
  AND U361 ( .A(n261), .B(n262), .Z(n8560) );
  XOR U362 ( .A(n8624), .B(n8623), .Z(n263) );
  NAND U363 ( .A(n263), .B(sreg[1335]), .Z(n264) );
  NAND U364 ( .A(n8624), .B(n8623), .Z(n265) );
  AND U365 ( .A(n264), .B(n265), .Z(n8644) );
  XOR U366 ( .A(n8844), .B(sreg[1345]), .Z(n266) );
  NAND U367 ( .A(n266), .B(n8843), .Z(n267) );
  NAND U368 ( .A(n8844), .B(sreg[1345]), .Z(n268) );
  AND U369 ( .A(n267), .B(n268), .Z(n8846) );
  NAND U370 ( .A(sreg[1357]), .B(n9109), .Z(n269) );
  XOR U371 ( .A(n9109), .B(sreg[1357]), .Z(n270) );
  NANDN U372 ( .A(n9110), .B(n270), .Z(n271) );
  NAND U373 ( .A(n269), .B(n271), .Z(n9112) );
  NAND U374 ( .A(n9219), .B(sreg[1362]), .Z(n272) );
  XOR U375 ( .A(sreg[1362]), .B(n9219), .Z(n273) );
  NAND U376 ( .A(n273), .B(n9218), .Z(n274) );
  NAND U377 ( .A(n272), .B(n274), .Z(n9239) );
  NAND U378 ( .A(sreg[1367]), .B(n9327), .Z(n275) );
  XOR U379 ( .A(n9327), .B(sreg[1367]), .Z(n276) );
  NANDN U380 ( .A(n9328), .B(n276), .Z(n277) );
  NAND U381 ( .A(n275), .B(n277), .Z(n9330) );
  NAND U382 ( .A(n9505), .B(sreg[1376]), .Z(n278) );
  XOR U383 ( .A(sreg[1376]), .B(n9505), .Z(n279) );
  NANDN U384 ( .A(n9506), .B(n279), .Z(n280) );
  NAND U385 ( .A(n278), .B(n280), .Z(n9539) );
  NAND U386 ( .A(sreg[1381]), .B(n9625), .Z(n281) );
  XOR U387 ( .A(n9625), .B(sreg[1381]), .Z(n282) );
  NANDN U388 ( .A(n9626), .B(n282), .Z(n283) );
  NAND U389 ( .A(n281), .B(n283), .Z(n9646) );
  XOR U390 ( .A(sreg[1387]), .B(n9739), .Z(n284) );
  NANDN U391 ( .A(n9740), .B(n284), .Z(n285) );
  NAND U392 ( .A(sreg[1387]), .B(n9739), .Z(n286) );
  AND U393 ( .A(n285), .B(n286), .Z(n9778) );
  XOR U394 ( .A(sreg[1401]), .B(n10041), .Z(n287) );
  NANDN U395 ( .A(n10042), .B(n287), .Z(n288) );
  NAND U396 ( .A(sreg[1401]), .B(n10041), .Z(n289) );
  AND U397 ( .A(n288), .B(n289), .Z(n10077) );
  NAND U398 ( .A(n10605), .B(sreg[1426]), .Z(n290) );
  XOR U399 ( .A(sreg[1426]), .B(n10605), .Z(n291) );
  NAND U400 ( .A(n291), .B(n10604), .Z(n292) );
  NAND U401 ( .A(n290), .B(n292), .Z(n10607) );
  XOR U402 ( .A(n11315), .B(sreg[1458]), .Z(n293) );
  NAND U403 ( .A(n293), .B(n11314), .Z(n294) );
  NAND U404 ( .A(n11315), .B(sreg[1458]), .Z(n295) );
  AND U405 ( .A(n294), .B(n295), .Z(n11317) );
  NAND U406 ( .A(n11571), .B(sreg[1470]), .Z(n296) );
  XOR U407 ( .A(sreg[1470]), .B(n11571), .Z(n297) );
  NAND U408 ( .A(n297), .B(n11570), .Z(n298) );
  NAND U409 ( .A(n296), .B(n298), .Z(n11592) );
  NAND U410 ( .A(n11884), .B(n11883), .Z(n299) );
  XOR U411 ( .A(n11883), .B(n11884), .Z(n300) );
  NAND U412 ( .A(n300), .B(sreg[1485]), .Z(n301) );
  NAND U413 ( .A(n299), .B(n301), .Z(n11923) );
  XOR U414 ( .A(n12009), .B(n12008), .Z(n302) );
  NAND U415 ( .A(n302), .B(sreg[1490]), .Z(n303) );
  NAND U416 ( .A(n12009), .B(n12008), .Z(n304) );
  AND U417 ( .A(n303), .B(n304), .Z(n12029) );
  NAND U418 ( .A(sreg[1495]), .B(n12117), .Z(n305) );
  XOR U419 ( .A(n12117), .B(sreg[1495]), .Z(n306) );
  NANDN U420 ( .A(n12118), .B(n306), .Z(n307) );
  NAND U421 ( .A(n305), .B(n307), .Z(n12138) );
  XOR U422 ( .A(n12249), .B(sreg[1502]), .Z(n308) );
  NANDN U423 ( .A(n12248), .B(n308), .Z(n309) );
  NAND U424 ( .A(n12249), .B(sreg[1502]), .Z(n310) );
  AND U425 ( .A(n309), .B(n310), .Z(n12270) );
  NAND U426 ( .A(sreg[1551]), .B(n13345), .Z(n311) );
  XOR U427 ( .A(n13345), .B(sreg[1551]), .Z(n312) );
  NANDN U428 ( .A(n13346), .B(n312), .Z(n313) );
  NAND U429 ( .A(n311), .B(n313), .Z(n13348) );
  NAND U430 ( .A(sreg[1559]), .B(n13521), .Z(n314) );
  XOR U431 ( .A(n13521), .B(sreg[1559]), .Z(n315) );
  NANDN U432 ( .A(n13522), .B(n315), .Z(n316) );
  NAND U433 ( .A(n314), .B(n316), .Z(n13542) );
  XOR U434 ( .A(sreg[1572]), .B(n13794), .Z(n317) );
  NANDN U435 ( .A(n13795), .B(n317), .Z(n318) );
  NAND U436 ( .A(sreg[1572]), .B(n13794), .Z(n319) );
  AND U437 ( .A(n318), .B(n319), .Z(n13834) );
  NAND U438 ( .A(sreg[1588]), .B(n14162), .Z(n320) );
  XOR U439 ( .A(n14162), .B(sreg[1588]), .Z(n321) );
  NANDN U440 ( .A(n14163), .B(n321), .Z(n322) );
  NAND U441 ( .A(n320), .B(n322), .Z(n14165) );
  NAND U442 ( .A(n14448), .B(n14447), .Z(n323) );
  XOR U443 ( .A(n14447), .B(n14448), .Z(n324) );
  NAND U444 ( .A(n324), .B(sreg[1601]), .Z(n325) );
  NAND U445 ( .A(n323), .B(n325), .Z(n14450) );
  NAND U446 ( .A(n14580), .B(sreg[1607]), .Z(n326) );
  XOR U447 ( .A(sreg[1607]), .B(n14580), .Z(n327) );
  NAND U448 ( .A(n327), .B(n14579), .Z(n328) );
  NAND U449 ( .A(n326), .B(n328), .Z(n14582) );
  NAND U450 ( .A(sreg[1613]), .B(n14711), .Z(n329) );
  XOR U451 ( .A(n14711), .B(sreg[1613]), .Z(n330) );
  NANDN U452 ( .A(n14712), .B(n330), .Z(n331) );
  NAND U453 ( .A(n329), .B(n331), .Z(n14714) );
  XOR U454 ( .A(n14886), .B(n14885), .Z(n332) );
  NANDN U455 ( .A(sreg[1621]), .B(n332), .Z(n333) );
  NAND U456 ( .A(n14886), .B(n14885), .Z(n334) );
  AND U457 ( .A(n333), .B(n334), .Z(n14888) );
  NAND U458 ( .A(sreg[1625]), .B(n14971), .Z(n335) );
  XOR U459 ( .A(n14971), .B(sreg[1625]), .Z(n336) );
  NANDN U460 ( .A(n14972), .B(n336), .Z(n337) );
  NAND U461 ( .A(n335), .B(n337), .Z(n14974) );
  NAND U462 ( .A(sreg[1631]), .B(n15101), .Z(n338) );
  XOR U463 ( .A(n15101), .B(sreg[1631]), .Z(n339) );
  NANDN U464 ( .A(n15102), .B(n339), .Z(n340) );
  NAND U465 ( .A(n338), .B(n340), .Z(n15104) );
  NAND U466 ( .A(n15349), .B(sreg[1643]), .Z(n341) );
  XOR U467 ( .A(sreg[1643]), .B(n15349), .Z(n342) );
  NANDN U468 ( .A(n15350), .B(n342), .Z(n343) );
  NAND U469 ( .A(n341), .B(n343), .Z(n15371) );
  XOR U470 ( .A(sreg[1647]), .B(n15435), .Z(n344) );
  NANDN U471 ( .A(n15436), .B(n344), .Z(n345) );
  NAND U472 ( .A(sreg[1647]), .B(n15435), .Z(n346) );
  AND U473 ( .A(n345), .B(n346), .Z(n15474) );
  XOR U474 ( .A(n15651), .B(n15650), .Z(n347) );
  NAND U475 ( .A(n347), .B(sreg[1656]), .Z(n348) );
  NAND U476 ( .A(n15651), .B(n15650), .Z(n349) );
  AND U477 ( .A(n348), .B(n349), .Z(n15671) );
  NAND U478 ( .A(n16108), .B(sreg[1677]), .Z(n350) );
  XOR U479 ( .A(sreg[1677]), .B(n16108), .Z(n351) );
  NANDN U480 ( .A(n16107), .B(n351), .Z(n352) );
  NAND U481 ( .A(n350), .B(n352), .Z(n16110) );
  NAND U482 ( .A(n16278), .B(sreg[1685]), .Z(n353) );
  XOR U483 ( .A(sreg[1685]), .B(n16278), .Z(n354) );
  NAND U484 ( .A(n354), .B(n16277), .Z(n355) );
  NAND U485 ( .A(n353), .B(n355), .Z(n16298) );
  NAND U486 ( .A(n16651), .B(n16650), .Z(n356) );
  XOR U487 ( .A(n16650), .B(n16651), .Z(n357) );
  NAND U488 ( .A(n357), .B(sreg[1702]), .Z(n358) );
  NAND U489 ( .A(n356), .B(n358), .Z(n16653) );
  XOR U490 ( .A(sreg[1707]), .B(n16741), .Z(n359) );
  NANDN U491 ( .A(n16742), .B(n359), .Z(n360) );
  NAND U492 ( .A(sreg[1707]), .B(n16741), .Z(n361) );
  AND U493 ( .A(n360), .B(n361), .Z(n16782) );
  NAND U494 ( .A(n16826), .B(n16825), .Z(n362) );
  XOR U495 ( .A(n16825), .B(n16826), .Z(n363) );
  NANDN U496 ( .A(sreg[1711]), .B(n363), .Z(n364) );
  NAND U497 ( .A(n362), .B(n364), .Z(n16861) );
  XOR U498 ( .A(sreg[1716]), .B(n16930), .Z(n365) );
  NANDN U499 ( .A(n16931), .B(n365), .Z(n366) );
  NAND U500 ( .A(sreg[1716]), .B(n16930), .Z(n367) );
  AND U501 ( .A(n366), .B(n367), .Z(n16969) );
  NAND U502 ( .A(n17017), .B(n17016), .Z(n368) );
  XOR U503 ( .A(n17016), .B(n17017), .Z(n369) );
  NANDN U504 ( .A(sreg[1720]), .B(n369), .Z(n370) );
  NAND U505 ( .A(n368), .B(n370), .Z(n17056) );
  NAND U506 ( .A(sreg[1731]), .B(n17275), .Z(n371) );
  XOR U507 ( .A(n17275), .B(sreg[1731]), .Z(n372) );
  NANDN U508 ( .A(n17276), .B(n372), .Z(n373) );
  NAND U509 ( .A(n371), .B(n373), .Z(n17278) );
  NAND U510 ( .A(sreg[1737]), .B(n17403), .Z(n374) );
  XOR U511 ( .A(n17403), .B(sreg[1737]), .Z(n375) );
  NANDN U512 ( .A(n17404), .B(n375), .Z(n376) );
  NAND U513 ( .A(n374), .B(n376), .Z(n17406) );
  XOR U514 ( .A(n18031), .B(sreg[1766]), .Z(n377) );
  NAND U515 ( .A(n377), .B(n18030), .Z(n378) );
  NAND U516 ( .A(n18031), .B(sreg[1766]), .Z(n379) );
  AND U517 ( .A(n378), .B(n379), .Z(n18052) );
  NAND U518 ( .A(n18445), .B(sreg[1784]), .Z(n380) );
  XOR U519 ( .A(sreg[1784]), .B(n18445), .Z(n381) );
  NAND U520 ( .A(n381), .B(n18444), .Z(n382) );
  NAND U521 ( .A(n380), .B(n382), .Z(n18447) );
  NAND U522 ( .A(n18574), .B(sreg[1790]), .Z(n383) );
  XOR U523 ( .A(sreg[1790]), .B(n18574), .Z(n384) );
  NANDN U524 ( .A(n18575), .B(n384), .Z(n385) );
  NAND U525 ( .A(n383), .B(n385), .Z(n18597) );
  NAND U526 ( .A(sreg[1798]), .B(n18746), .Z(n386) );
  XOR U527 ( .A(n18746), .B(sreg[1798]), .Z(n387) );
  NANDN U528 ( .A(n18747), .B(n387), .Z(n388) );
  NAND U529 ( .A(n386), .B(n388), .Z(n18749) );
  XOR U530 ( .A(n19011), .B(n19010), .Z(n389) );
  NAND U531 ( .A(n389), .B(sreg[1810]), .Z(n390) );
  NAND U532 ( .A(n19011), .B(n19010), .Z(n391) );
  AND U533 ( .A(n390), .B(n391), .Z(n19031) );
  NAND U534 ( .A(sreg[1815]), .B(n19119), .Z(n392) );
  XOR U535 ( .A(n19119), .B(sreg[1815]), .Z(n393) );
  NANDN U536 ( .A(n19120), .B(n393), .Z(n394) );
  NAND U537 ( .A(n392), .B(n394), .Z(n19122) );
  XOR U538 ( .A(n19504), .B(n19503), .Z(n395) );
  NAND U539 ( .A(n395), .B(sreg[1833]), .Z(n396) );
  NAND U540 ( .A(n19504), .B(n19503), .Z(n397) );
  AND U541 ( .A(n396), .B(n397), .Z(n19524) );
  NAND U542 ( .A(sreg[1837]), .B(n19589), .Z(n398) );
  XOR U543 ( .A(n19589), .B(sreg[1837]), .Z(n399) );
  NANDN U544 ( .A(n19590), .B(n399), .Z(n400) );
  NAND U545 ( .A(n398), .B(n400), .Z(n19592) );
  NAND U546 ( .A(n19681), .B(sreg[1842]), .Z(n401) );
  XOR U547 ( .A(sreg[1842]), .B(n19681), .Z(n402) );
  NANDN U548 ( .A(n19680), .B(n402), .Z(n403) );
  NAND U549 ( .A(n401), .B(n403), .Z(n19701) );
  NAND U550 ( .A(sreg[1847]), .B(n19807), .Z(n404) );
  XOR U551 ( .A(n19807), .B(sreg[1847]), .Z(n405) );
  NANDN U552 ( .A(n19808), .B(n405), .Z(n406) );
  NAND U553 ( .A(n404), .B(n406), .Z(n19810) );
  XOR U554 ( .A(n20007), .B(n20006), .Z(n407) );
  NAND U555 ( .A(n407), .B(sreg[1856]), .Z(n408) );
  NAND U556 ( .A(n20007), .B(n20006), .Z(n409) );
  AND U557 ( .A(n408), .B(n409), .Z(n20027) );
  NAND U558 ( .A(n20292), .B(sreg[1869]), .Z(n410) );
  XOR U559 ( .A(sreg[1869]), .B(n20292), .Z(n411) );
  NANDN U560 ( .A(n20291), .B(n411), .Z(n412) );
  NAND U561 ( .A(n410), .B(n412), .Z(n20294) );
  NAND U562 ( .A(sreg[1887]), .B(n20682), .Z(n413) );
  XOR U563 ( .A(n20682), .B(sreg[1887]), .Z(n414) );
  NANDN U564 ( .A(n20683), .B(n414), .Z(n415) );
  NAND U565 ( .A(n413), .B(n415), .Z(n20685) );
  NAND U566 ( .A(n20768), .B(sreg[1892]), .Z(n416) );
  XOR U567 ( .A(sreg[1892]), .B(n20768), .Z(n417) );
  NANDN U568 ( .A(n20769), .B(n417), .Z(n418) );
  NAND U569 ( .A(n416), .B(n418), .Z(n20790) );
  NAND U570 ( .A(sreg[1897]), .B(n20895), .Z(n419) );
  XOR U571 ( .A(n20895), .B(sreg[1897]), .Z(n420) );
  NANDN U572 ( .A(n20896), .B(n420), .Z(n421) );
  NAND U573 ( .A(n419), .B(n421), .Z(n20898) );
  NAND U574 ( .A(n21075), .B(n21074), .Z(n422) );
  XOR U575 ( .A(n21074), .B(n21075), .Z(n423) );
  NAND U576 ( .A(n423), .B(sreg[1906]), .Z(n424) );
  NAND U577 ( .A(n422), .B(n424), .Z(n21095) );
  NAND U578 ( .A(n21202), .B(sreg[1911]), .Z(n425) );
  XOR U579 ( .A(sreg[1911]), .B(n21202), .Z(n426) );
  NANDN U580 ( .A(n21201), .B(n426), .Z(n427) );
  NAND U581 ( .A(n425), .B(n427), .Z(n21204) );
  NAND U582 ( .A(sreg[1915]), .B(n21287), .Z(n428) );
  XOR U583 ( .A(n21287), .B(sreg[1915]), .Z(n429) );
  NANDN U584 ( .A(n21288), .B(n429), .Z(n430) );
  NAND U585 ( .A(n428), .B(n430), .Z(n21290) );
  NAND U586 ( .A(sreg[1922]), .B(n21440), .Z(n431) );
  XOR U587 ( .A(n21440), .B(sreg[1922]), .Z(n432) );
  NANDN U588 ( .A(n21441), .B(n432), .Z(n433) );
  NAND U589 ( .A(n431), .B(n433), .Z(n21443) );
  NAND U590 ( .A(n21548), .B(n21547), .Z(n434) );
  XOR U591 ( .A(n21547), .B(n21548), .Z(n435) );
  NANDN U592 ( .A(sreg[1927]), .B(n435), .Z(n436) );
  NAND U593 ( .A(n434), .B(n436), .Z(n21568) );
  NAND U594 ( .A(n21970), .B(n21969), .Z(n437) );
  XOR U595 ( .A(n21969), .B(n21970), .Z(n438) );
  NAND U596 ( .A(n438), .B(sreg[1947]), .Z(n439) );
  NAND U597 ( .A(n437), .B(n439), .Z(n22008) );
  NAND U598 ( .A(sreg[1960]), .B(n22270), .Z(n440) );
  XOR U599 ( .A(n22270), .B(sreg[1960]), .Z(n441) );
  NANDN U600 ( .A(n22271), .B(n441), .Z(n442) );
  NAND U601 ( .A(n440), .B(n442), .Z(n22291) );
  NAND U602 ( .A(n22955), .B(sreg[1991]), .Z(n443) );
  XOR U603 ( .A(sreg[1991]), .B(n22955), .Z(n444) );
  NANDN U604 ( .A(n22956), .B(n444), .Z(n445) );
  NAND U605 ( .A(n443), .B(n445), .Z(n22958) );
  NAND U606 ( .A(n23023), .B(sreg[1995]), .Z(n446) );
  XOR U607 ( .A(sreg[1995]), .B(n23023), .Z(n447) );
  NANDN U608 ( .A(n23024), .B(n447), .Z(n448) );
  NAND U609 ( .A(n446), .B(n448), .Z(n23044) );
  NAND U610 ( .A(sreg[2004]), .B(n23234), .Z(n449) );
  XOR U611 ( .A(n23234), .B(sreg[2004]), .Z(n450) );
  NANDN U612 ( .A(n23235), .B(n450), .Z(n451) );
  NAND U613 ( .A(n449), .B(n451), .Z(n23237) );
  XOR U614 ( .A(n23587), .B(sreg[2020]), .Z(n452) );
  NANDN U615 ( .A(n23586), .B(n452), .Z(n453) );
  NAND U616 ( .A(n23587), .B(sreg[2020]), .Z(n454) );
  AND U617 ( .A(n453), .B(n454), .Z(n23607) );
  NAND U618 ( .A(sreg[2024]), .B(n23672), .Z(n455) );
  XOR U619 ( .A(n23672), .B(sreg[2024]), .Z(n456) );
  NANDN U620 ( .A(n23673), .B(n456), .Z(n457) );
  NAND U621 ( .A(n455), .B(n457), .Z(n23693) );
  AND U622 ( .A(b[0]), .B(a[1]), .Z(n1843) );
  NANDN U623 ( .A(n18605), .B(n18604), .Z(n458) );
  NANDN U624 ( .A(n18606), .B(n18607), .Z(n459) );
  NAND U625 ( .A(n458), .B(n459), .Z(n18631) );
  NANDN U626 ( .A(n22112), .B(n22111), .Z(n460) );
  NANDN U627 ( .A(n22113), .B(n22114), .Z(n461) );
  NAND U628 ( .A(n460), .B(n461), .Z(n22116) );
  NANDN U629 ( .A(n2543), .B(n2542), .Z(n462) );
  NANDN U630 ( .A(n2544), .B(n2545), .Z(n463) );
  NAND U631 ( .A(n462), .B(n463), .Z(n2564) );
  NAND U632 ( .A(n7720), .B(n7718), .Z(n464) );
  XOR U633 ( .A(n7718), .B(n7720), .Z(n465) );
  NANDN U634 ( .A(n7719), .B(n465), .Z(n466) );
  NAND U635 ( .A(n464), .B(n466), .Z(n7736) );
  NANDN U636 ( .A(n8127), .B(n8126), .Z(n467) );
  NANDN U637 ( .A(n8128), .B(n8129), .Z(n468) );
  NAND U638 ( .A(n467), .B(n468), .Z(n8148) );
  NANDN U639 ( .A(n8491), .B(n8490), .Z(n469) );
  NANDN U640 ( .A(n8492), .B(n8493), .Z(n470) );
  NAND U641 ( .A(n469), .B(n470), .Z(n8501) );
  NANDN U642 ( .A(n10073), .B(n10072), .Z(n471) );
  NANDN U643 ( .A(n10074), .B(n10075), .Z(n472) );
  NAND U644 ( .A(n471), .B(n472), .Z(n10082) );
  NAND U645 ( .A(n10189), .B(n10188), .Z(n473) );
  XOR U646 ( .A(n10188), .B(n10189), .Z(n474) );
  NANDN U647 ( .A(n10190), .B(n474), .Z(n475) );
  NAND U648 ( .A(n473), .B(n475), .Z(n10213) );
  NAND U649 ( .A(n11474), .B(n11473), .Z(n476) );
  XOR U650 ( .A(n11473), .B(n11474), .Z(n477) );
  NANDN U651 ( .A(n11475), .B(n477), .Z(n478) );
  NAND U652 ( .A(n476), .B(n478), .Z(n11488) );
  NAND U653 ( .A(n11598), .B(n11597), .Z(n479) );
  XOR U654 ( .A(n11597), .B(n11598), .Z(n480) );
  NANDN U655 ( .A(n11599), .B(n480), .Z(n481) );
  NAND U656 ( .A(n479), .B(n481), .Z(n11625) );
  NANDN U657 ( .A(n12303), .B(n12302), .Z(n482) );
  NANDN U658 ( .A(n12304), .B(n12305), .Z(n483) );
  NAND U659 ( .A(n482), .B(n483), .Z(n12312) );
  NAND U660 ( .A(n12999), .B(n12998), .Z(n484) );
  XOR U661 ( .A(n12998), .B(n12999), .Z(n485) );
  NANDN U662 ( .A(n13000), .B(n485), .Z(n486) );
  NAND U663 ( .A(n484), .B(n486), .Z(n13019) );
  NANDN U664 ( .A(n16161), .B(n16160), .Z(n487) );
  NANDN U665 ( .A(n16162), .B(n16163), .Z(n488) );
  NAND U666 ( .A(n487), .B(n488), .Z(n16182) );
  XOR U667 ( .A(n17499), .B(n17498), .Z(n489) );
  NANDN U668 ( .A(n17497), .B(n489), .Z(n490) );
  NAND U669 ( .A(n17499), .B(n17498), .Z(n491) );
  AND U670 ( .A(n490), .B(n491), .Z(n17515) );
  NANDN U671 ( .A(n20691), .B(n20690), .Z(n492) );
  NANDN U672 ( .A(n20692), .B(n20693), .Z(n493) );
  NAND U673 ( .A(n492), .B(n493), .Z(n20712) );
  XOR U674 ( .A(n22039), .B(n22038), .Z(n494) );
  NANDN U675 ( .A(n22037), .B(n494), .Z(n495) );
  NAND U676 ( .A(n22039), .B(n22038), .Z(n496) );
  AND U677 ( .A(n495), .B(n496), .Z(n22055) );
  OR U678 ( .A(n24064), .B(n24065), .Z(n497) );
  NAND U679 ( .A(n24066), .B(n24067), .Z(n498) );
  AND U680 ( .A(n497), .B(n498), .Z(n24073) );
  NAND U681 ( .A(n2478), .B(n2476), .Z(n499) );
  XOR U682 ( .A(n2476), .B(n2478), .Z(n500) );
  NANDN U683 ( .A(n2477), .B(n500), .Z(n501) );
  NAND U684 ( .A(n499), .B(n501), .Z(n2497) );
  NAND U685 ( .A(n7090), .B(n7089), .Z(n502) );
  XOR U686 ( .A(n7089), .B(n7090), .Z(n503) );
  NANDN U687 ( .A(n7091), .B(n503), .Z(n504) );
  NAND U688 ( .A(n502), .B(n504), .Z(n7120) );
  XOR U689 ( .A(n8062), .B(n8061), .Z(n505) );
  NANDN U690 ( .A(n8060), .B(n505), .Z(n506) );
  NAND U691 ( .A(n8062), .B(n8061), .Z(n507) );
  AND U692 ( .A(n506), .B(n507), .Z(n8083) );
  NAND U693 ( .A(n9935), .B(n9934), .Z(n508) );
  XOR U694 ( .A(n9934), .B(n9935), .Z(n509) );
  NANDN U695 ( .A(n9936), .B(n509), .Z(n510) );
  NAND U696 ( .A(n508), .B(n510), .Z(n9957) );
  XOR U697 ( .A(n12232), .B(n12231), .Z(n511) );
  NANDN U698 ( .A(n12230), .B(n511), .Z(n512) );
  NAND U699 ( .A(n12232), .B(n12231), .Z(n513) );
  AND U700 ( .A(n512), .B(n513), .Z(n12253) );
  XOR U701 ( .A(sreg[1526]), .B(n12794), .Z(n514) );
  NANDN U702 ( .A(n12795), .B(n514), .Z(n515) );
  NAND U703 ( .A(sreg[1526]), .B(n12794), .Z(n516) );
  AND U704 ( .A(n515), .B(n516), .Z(n12816) );
  NAND U705 ( .A(n16094), .B(n16092), .Z(n517) );
  XOR U706 ( .A(n16092), .B(n16094), .Z(n518) );
  NANDN U707 ( .A(n16093), .B(n518), .Z(n519) );
  NAND U708 ( .A(n517), .B(n519), .Z(n16115) );
  NAND U709 ( .A(n19315), .B(n19314), .Z(n520) );
  XOR U710 ( .A(n19314), .B(n19315), .Z(n521) );
  NAND U711 ( .A(n521), .B(n19313), .Z(n522) );
  NAND U712 ( .A(n520), .B(n522), .Z(n19336) );
  NAND U713 ( .A(n20623), .B(n20621), .Z(n523) );
  XOR U714 ( .A(n20621), .B(n20623), .Z(n524) );
  NANDN U715 ( .A(n20622), .B(n524), .Z(n525) );
  NAND U716 ( .A(n523), .B(n525), .Z(n20645) );
  XOR U717 ( .A(n1901), .B(n1900), .Z(n526) );
  NANDN U718 ( .A(sreg[1026]), .B(n526), .Z(n527) );
  NAND U719 ( .A(n1901), .B(n1900), .Z(n528) );
  AND U720 ( .A(n527), .B(n528), .Z(n1903) );
  NAND U721 ( .A(n2036), .B(sreg[1033]), .Z(n529) );
  XOR U722 ( .A(sreg[1033]), .B(n2036), .Z(n530) );
  NANDN U723 ( .A(n2035), .B(n530), .Z(n531) );
  NAND U724 ( .A(n529), .B(n531), .Z(n2074) );
  XOR U725 ( .A(sreg[1038]), .B(n2146), .Z(n532) );
  NANDN U726 ( .A(n2147), .B(n532), .Z(n533) );
  NAND U727 ( .A(sreg[1038]), .B(n2146), .Z(n534) );
  AND U728 ( .A(n533), .B(n534), .Z(n2186) );
  XOR U729 ( .A(sreg[1043]), .B(n2257), .Z(n535) );
  NANDN U730 ( .A(n2258), .B(n535), .Z(n536) );
  NAND U731 ( .A(sreg[1043]), .B(n2257), .Z(n537) );
  AND U732 ( .A(n536), .B(n537), .Z(n2296) );
  NAND U733 ( .A(sreg[1047]), .B(n2363), .Z(n538) );
  XOR U734 ( .A(n2363), .B(sreg[1047]), .Z(n539) );
  NANDN U735 ( .A(n2364), .B(n539), .Z(n540) );
  NAND U736 ( .A(n538), .B(n540), .Z(n2384) );
  XOR U737 ( .A(sreg[1051]), .B(n2431), .Z(n541) );
  NANDN U738 ( .A(n2432), .B(n541), .Z(n542) );
  NAND U739 ( .A(sreg[1051]), .B(n2431), .Z(n543) );
  AND U740 ( .A(n542), .B(n543), .Z(n2471) );
  NAND U741 ( .A(n2537), .B(sreg[1056]), .Z(n544) );
  XOR U742 ( .A(sreg[1056]), .B(n2537), .Z(n545) );
  NANDN U743 ( .A(n2538), .B(n545), .Z(n546) );
  NAND U744 ( .A(n544), .B(n546), .Z(n2571) );
  NAND U745 ( .A(n2686), .B(n2685), .Z(n547) );
  XOR U746 ( .A(n2685), .B(n2686), .Z(n548) );
  NAND U747 ( .A(n548), .B(sreg[1063]), .Z(n549) );
  NAND U748 ( .A(n547), .B(n549), .Z(n2724) );
  XOR U749 ( .A(n2884), .B(sreg[1071]), .Z(n550) );
  NANDN U750 ( .A(n2883), .B(n550), .Z(n551) );
  NAND U751 ( .A(n2884), .B(sreg[1071]), .Z(n552) );
  AND U752 ( .A(n551), .B(n552), .Z(n2886) );
  XOR U753 ( .A(sreg[1075]), .B(n2953), .Z(n553) );
  NANDN U754 ( .A(n2954), .B(n553), .Z(n554) );
  NAND U755 ( .A(sreg[1075]), .B(n2953), .Z(n555) );
  AND U756 ( .A(n554), .B(n555), .Z(n2993) );
  NAND U757 ( .A(sreg[1081]), .B(n3103), .Z(n556) );
  XOR U758 ( .A(n3103), .B(sreg[1081]), .Z(n557) );
  NANDN U759 ( .A(n3104), .B(n557), .Z(n558) );
  NAND U760 ( .A(n556), .B(n558), .Z(n3106) );
  NAND U761 ( .A(n3190), .B(sreg[1085]), .Z(n559) );
  XOR U762 ( .A(sreg[1085]), .B(n3190), .Z(n560) );
  NAND U763 ( .A(n560), .B(n3189), .Z(n561) );
  NAND U764 ( .A(n559), .B(n561), .Z(n3192) );
  NAND U765 ( .A(n3274), .B(n3273), .Z(n562) );
  XOR U766 ( .A(n3273), .B(n3274), .Z(n563) );
  NANDN U767 ( .A(sreg[1089]), .B(n563), .Z(n564) );
  NAND U768 ( .A(n562), .B(n564), .Z(n3276) );
  XOR U769 ( .A(sreg[1093]), .B(n3341), .Z(n565) );
  NANDN U770 ( .A(n3342), .B(n565), .Z(n566) );
  NAND U771 ( .A(sreg[1093]), .B(n3341), .Z(n567) );
  AND U772 ( .A(n566), .B(n567), .Z(n3381) );
  NAND U773 ( .A(sreg[1098]), .B(n3468), .Z(n568) );
  XOR U774 ( .A(n3468), .B(sreg[1098]), .Z(n569) );
  NANDN U775 ( .A(n3469), .B(n569), .Z(n570) );
  NAND U776 ( .A(n568), .B(n570), .Z(n3489) );
  NAND U777 ( .A(n3535), .B(n3534), .Z(n571) );
  XOR U778 ( .A(n3534), .B(n3535), .Z(n572) );
  NANDN U779 ( .A(sreg[1102]), .B(n572), .Z(n573) );
  NAND U780 ( .A(n571), .B(n573), .Z(n3574) );
  NAND U781 ( .A(sreg[1108]), .B(n3682), .Z(n574) );
  XOR U782 ( .A(n3682), .B(sreg[1108]), .Z(n575) );
  NANDN U783 ( .A(n3683), .B(n575), .Z(n576) );
  NAND U784 ( .A(n574), .B(n576), .Z(n3685) );
  XOR U785 ( .A(n3753), .B(sreg[1112]), .Z(n577) );
  NAND U786 ( .A(n577), .B(n3752), .Z(n578) );
  NAND U787 ( .A(n3753), .B(sreg[1112]), .Z(n579) );
  AND U788 ( .A(n578), .B(n579), .Z(n3792) );
  NAND U789 ( .A(n3903), .B(sreg[1118]), .Z(n580) );
  XOR U790 ( .A(sreg[1118]), .B(n3903), .Z(n581) );
  NAND U791 ( .A(n581), .B(n3902), .Z(n582) );
  NAND U792 ( .A(n580), .B(n582), .Z(n3924) );
  XOR U793 ( .A(sreg[1122]), .B(n3966), .Z(n583) );
  NANDN U794 ( .A(n3967), .B(n583), .Z(n584) );
  NAND U795 ( .A(sreg[1122]), .B(n3966), .Z(n585) );
  AND U796 ( .A(n584), .B(n585), .Z(n4006) );
  XOR U797 ( .A(n4140), .B(sreg[1129]), .Z(n586) );
  NANDN U798 ( .A(n4139), .B(n586), .Z(n587) );
  NAND U799 ( .A(n4140), .B(sreg[1129]), .Z(n588) );
  AND U800 ( .A(n587), .B(n588), .Z(n4142) );
  XOR U801 ( .A(sreg[1136]), .B(n4278), .Z(n589) );
  NANDN U802 ( .A(n4279), .B(n589), .Z(n590) );
  NAND U803 ( .A(sreg[1136]), .B(n4278), .Z(n591) );
  AND U804 ( .A(n590), .B(n591), .Z(n4318) );
  NAND U805 ( .A(n4404), .B(sreg[1141]), .Z(n592) );
  XOR U806 ( .A(sreg[1141]), .B(n4404), .Z(n593) );
  NAND U807 ( .A(n593), .B(n4403), .Z(n594) );
  NAND U808 ( .A(n592), .B(n594), .Z(n4424) );
  NAND U809 ( .A(sreg[1145]), .B(n4489), .Z(n595) );
  XOR U810 ( .A(n4489), .B(sreg[1145]), .Z(n596) );
  NANDN U811 ( .A(n4490), .B(n596), .Z(n597) );
  NAND U812 ( .A(n595), .B(n597), .Z(n4492) );
  XOR U813 ( .A(sreg[1155]), .B(n4695), .Z(n598) );
  NANDN U814 ( .A(n4696), .B(n598), .Z(n599) );
  NAND U815 ( .A(sreg[1155]), .B(n4695), .Z(n600) );
  AND U816 ( .A(n599), .B(n600), .Z(n4735) );
  XOR U817 ( .A(sreg[1159]), .B(n4783), .Z(n601) );
  NANDN U818 ( .A(n4784), .B(n601), .Z(n602) );
  NAND U819 ( .A(sreg[1159]), .B(n4783), .Z(n603) );
  AND U820 ( .A(n602), .B(n603), .Z(n4823) );
  NAND U821 ( .A(n4959), .B(sreg[1166]), .Z(n604) );
  XOR U822 ( .A(sreg[1166]), .B(n4959), .Z(n605) );
  NAND U823 ( .A(n605), .B(n4958), .Z(n606) );
  NAND U824 ( .A(n604), .B(n606), .Z(n4961) );
  NAND U825 ( .A(n5094), .B(n5093), .Z(n607) );
  XOR U826 ( .A(n5093), .B(n5094), .Z(n608) );
  NAND U827 ( .A(n608), .B(sreg[1173]), .Z(n609) );
  NAND U828 ( .A(n607), .B(n609), .Z(n5115) );
  NAND U829 ( .A(n5182), .B(n5181), .Z(n610) );
  XOR U830 ( .A(n5181), .B(n5182), .Z(n611) );
  NAND U831 ( .A(n611), .B(sreg[1177]), .Z(n612) );
  NAND U832 ( .A(n610), .B(n612), .Z(n5220) );
  XOR U833 ( .A(sreg[1182]), .B(n5292), .Z(n613) );
  NANDN U834 ( .A(n5293), .B(n613), .Z(n614) );
  NAND U835 ( .A(sreg[1182]), .B(n5292), .Z(n615) );
  AND U836 ( .A(n614), .B(n615), .Z(n5332) );
  NAND U837 ( .A(n5381), .B(n5380), .Z(n616) );
  XOR U838 ( .A(n5380), .B(n5381), .Z(n617) );
  NAND U839 ( .A(n617), .B(sreg[1186]), .Z(n618) );
  NAND U840 ( .A(n616), .B(n618), .Z(n5419) );
  XOR U841 ( .A(sreg[1193]), .B(n5537), .Z(n619) );
  NANDN U842 ( .A(n5538), .B(n619), .Z(n620) );
  NAND U843 ( .A(sreg[1193]), .B(n5537), .Z(n621) );
  AND U844 ( .A(n620), .B(n621), .Z(n5559) );
  XOR U845 ( .A(n5646), .B(sreg[1198]), .Z(n622) );
  NANDN U846 ( .A(n5645), .B(n622), .Z(n623) );
  NAND U847 ( .A(n5646), .B(sreg[1198]), .Z(n624) );
  AND U848 ( .A(n623), .B(n624), .Z(n5664) );
  XOR U849 ( .A(n5727), .B(n5726), .Z(n625) );
  NANDN U850 ( .A(sreg[1202]), .B(n625), .Z(n626) );
  NAND U851 ( .A(n5727), .B(n5726), .Z(n627) );
  AND U852 ( .A(n626), .B(n627), .Z(n5748) );
  XOR U853 ( .A(sreg[1208]), .B(n5860), .Z(n628) );
  NANDN U854 ( .A(n5861), .B(n628), .Z(n629) );
  NAND U855 ( .A(sreg[1208]), .B(n5860), .Z(n630) );
  AND U856 ( .A(n629), .B(n630), .Z(n5900) );
  NAND U857 ( .A(sreg[1214]), .B(n6010), .Z(n631) );
  XOR U858 ( .A(n6010), .B(sreg[1214]), .Z(n632) );
  NANDN U859 ( .A(n6011), .B(n632), .Z(n633) );
  NAND U860 ( .A(n631), .B(n633), .Z(n6031) );
  XOR U861 ( .A(n6079), .B(sreg[1218]), .Z(n634) );
  NAND U862 ( .A(n634), .B(n6078), .Z(n635) );
  NAND U863 ( .A(n6079), .B(sreg[1218]), .Z(n636) );
  AND U864 ( .A(n635), .B(n636), .Z(n6118) );
  NAND U865 ( .A(n6232), .B(n6231), .Z(n637) );
  XOR U866 ( .A(n6231), .B(n6232), .Z(n638) );
  NANDN U867 ( .A(sreg[1225]), .B(n638), .Z(n639) );
  NAND U868 ( .A(n637), .B(n639), .Z(n6253) );
  XOR U869 ( .A(sreg[1230]), .B(n6344), .Z(n640) );
  NANDN U870 ( .A(n6345), .B(n640), .Z(n641) );
  NAND U871 ( .A(sreg[1230]), .B(n6344), .Z(n642) );
  AND U872 ( .A(n641), .B(n642), .Z(n6384) );
  NAND U873 ( .A(n6433), .B(n6432), .Z(n643) );
  XOR U874 ( .A(n6432), .B(n6433), .Z(n644) );
  NANDN U875 ( .A(sreg[1234]), .B(n644), .Z(n645) );
  NAND U876 ( .A(n643), .B(n645), .Z(n6472) );
  NAND U877 ( .A(n6587), .B(sreg[1241]), .Z(n646) );
  XOR U878 ( .A(sreg[1241]), .B(n6587), .Z(n647) );
  NANDN U879 ( .A(n6588), .B(n647), .Z(n648) );
  NAND U880 ( .A(n646), .B(n648), .Z(n6628) );
  XOR U881 ( .A(sreg[1245]), .B(n6671), .Z(n649) );
  NANDN U882 ( .A(n6672), .B(n649), .Z(n650) );
  NAND U883 ( .A(sreg[1245]), .B(n6671), .Z(n651) );
  AND U884 ( .A(n650), .B(n651), .Z(n6710) );
  NAND U885 ( .A(n6779), .B(n6778), .Z(n652) );
  XOR U886 ( .A(n6778), .B(n6779), .Z(n653) );
  NANDN U887 ( .A(sreg[1250]), .B(n653), .Z(n654) );
  NAND U888 ( .A(n652), .B(n654), .Z(n6818) );
  NAND U889 ( .A(n6977), .B(n6976), .Z(n655) );
  XOR U890 ( .A(n6976), .B(n6977), .Z(n656) );
  NAND U891 ( .A(n656), .B(sreg[1258]), .Z(n657) );
  NAND U892 ( .A(n655), .B(n657), .Z(n6979) );
  XOR U893 ( .A(n7045), .B(sreg[1262]), .Z(n658) );
  NAND U894 ( .A(n658), .B(n7044), .Z(n659) );
  NAND U895 ( .A(n7045), .B(sreg[1262]), .Z(n660) );
  AND U896 ( .A(n659), .B(n660), .Z(n7066) );
  NAND U897 ( .A(sreg[1267]), .B(n7165), .Z(n661) );
  XOR U898 ( .A(n7165), .B(sreg[1267]), .Z(n662) );
  NANDN U899 ( .A(n7166), .B(n662), .Z(n663) );
  NAND U900 ( .A(n661), .B(n663), .Z(n7186) );
  NAND U901 ( .A(n7234), .B(sreg[1271]), .Z(n664) );
  XOR U902 ( .A(sreg[1271]), .B(n7234), .Z(n665) );
  NANDN U903 ( .A(n7233), .B(n665), .Z(n666) );
  NAND U904 ( .A(n664), .B(n666), .Z(n7272) );
  NAND U905 ( .A(n7409), .B(sreg[1278]), .Z(n667) );
  XOR U906 ( .A(sreg[1278]), .B(n7409), .Z(n668) );
  NANDN U907 ( .A(n7408), .B(n668), .Z(n669) );
  NAND U908 ( .A(n667), .B(n669), .Z(n7411) );
  NAND U909 ( .A(sreg[1284]), .B(n7536), .Z(n670) );
  XOR U910 ( .A(n7536), .B(sreg[1284]), .Z(n671) );
  NANDN U911 ( .A(n7537), .B(n671), .Z(n672) );
  NAND U912 ( .A(n670), .B(n672), .Z(n7539) );
  NAND U913 ( .A(n7605), .B(n7604), .Z(n673) );
  XOR U914 ( .A(n7604), .B(n7605), .Z(n674) );
  NANDN U915 ( .A(sreg[1288]), .B(n674), .Z(n675) );
  NAND U916 ( .A(n673), .B(n675), .Z(n7644) );
  XOR U917 ( .A(sreg[1292]), .B(n7690), .Z(n676) );
  NANDN U918 ( .A(n7691), .B(n676), .Z(n677) );
  NAND U919 ( .A(sreg[1292]), .B(n7690), .Z(n678) );
  AND U920 ( .A(n677), .B(n678), .Z(n7714) );
  NAND U921 ( .A(n7819), .B(n7818), .Z(n679) );
  XOR U922 ( .A(n7818), .B(n7819), .Z(n680) );
  NAND U923 ( .A(n680), .B(sreg[1298]), .Z(n681) );
  NAND U924 ( .A(n679), .B(n681), .Z(n7857) );
  NAND U925 ( .A(n7969), .B(n7968), .Z(n682) );
  XOR U926 ( .A(n7968), .B(n7969), .Z(n683) );
  NAND U927 ( .A(n683), .B(sreg[1304]), .Z(n684) );
  NAND U928 ( .A(n682), .B(n684), .Z(n7971) );
  NAND U929 ( .A(sreg[1308]), .B(n8057), .Z(n685) );
  XOR U930 ( .A(n8057), .B(sreg[1308]), .Z(n686) );
  NANDN U931 ( .A(n8058), .B(n686), .Z(n687) );
  NAND U932 ( .A(n685), .B(n687), .Z(n8076) );
  XOR U933 ( .A(sreg[1312]), .B(n8121), .Z(n688) );
  NANDN U934 ( .A(n8122), .B(n688), .Z(n689) );
  NAND U935 ( .A(sreg[1312]), .B(n8121), .Z(n690) );
  AND U936 ( .A(n689), .B(n690), .Z(n8156) );
  NAND U937 ( .A(n8242), .B(n8241), .Z(n691) );
  XOR U938 ( .A(n8241), .B(n8242), .Z(n692) );
  NAND U939 ( .A(n692), .B(sreg[1317]), .Z(n693) );
  NAND U940 ( .A(n691), .B(n693), .Z(n8244) );
  XOR U941 ( .A(sreg[1321]), .B(n8309), .Z(n694) );
  NANDN U942 ( .A(n8310), .B(n694), .Z(n695) );
  NAND U943 ( .A(sreg[1321]), .B(n8309), .Z(n696) );
  AND U944 ( .A(n695), .B(n696), .Z(n8349) );
  NAND U945 ( .A(n8435), .B(n8434), .Z(n697) );
  XOR U946 ( .A(n8434), .B(n8435), .Z(n698) );
  NAND U947 ( .A(n698), .B(sreg[1326]), .Z(n699) );
  NAND U948 ( .A(n697), .B(n699), .Z(n8437) );
  NAND U949 ( .A(n8561), .B(sreg[1332]), .Z(n700) );
  XOR U950 ( .A(sreg[1332]), .B(n8561), .Z(n701) );
  NANDN U951 ( .A(n8560), .B(n701), .Z(n702) );
  NAND U952 ( .A(n700), .B(n702), .Z(n8581) );
  XOR U953 ( .A(n8645), .B(n8644), .Z(n703) );
  NANDN U954 ( .A(sreg[1336]), .B(n703), .Z(n704) );
  NAND U955 ( .A(n8645), .B(n8644), .Z(n705) );
  AND U956 ( .A(n704), .B(n705), .Z(n8647) );
  XOR U957 ( .A(sreg[1340]), .B(n8714), .Z(n706) );
  NANDN U958 ( .A(n8715), .B(n706), .Z(n707) );
  NAND U959 ( .A(sreg[1340]), .B(n8714), .Z(n708) );
  AND U960 ( .A(n707), .B(n708), .Z(n8754) );
  XOR U961 ( .A(n8847), .B(sreg[1346]), .Z(n709) );
  NANDN U962 ( .A(n8846), .B(n709), .Z(n710) );
  NAND U963 ( .A(n8847), .B(sreg[1346]), .Z(n711) );
  AND U964 ( .A(n710), .B(n711), .Z(n8886) );
  NAND U965 ( .A(sreg[1354]), .B(n9044), .Z(n712) );
  XOR U966 ( .A(n9044), .B(sreg[1354]), .Z(n713) );
  NANDN U967 ( .A(n9045), .B(n713), .Z(n714) );
  NAND U968 ( .A(n712), .B(n714), .Z(n9047) );
  NAND U969 ( .A(n9113), .B(n9112), .Z(n715) );
  XOR U970 ( .A(n9112), .B(n9113), .Z(n716) );
  NAND U971 ( .A(n716), .B(sreg[1358]), .Z(n717) );
  NAND U972 ( .A(n715), .B(n717), .Z(n9151) );
  XOR U973 ( .A(n9240), .B(n9239), .Z(n718) );
  NAND U974 ( .A(n718), .B(sreg[1363]), .Z(n719) );
  NAND U975 ( .A(n9240), .B(n9239), .Z(n720) );
  AND U976 ( .A(n719), .B(n720), .Z(n9242) );
  NAND U977 ( .A(n9330), .B(sreg[1368]), .Z(n721) );
  XOR U978 ( .A(sreg[1368]), .B(n9330), .Z(n722) );
  NANDN U979 ( .A(n9331), .B(n722), .Z(n723) );
  NAND U980 ( .A(n721), .B(n723), .Z(n9351) );
  NAND U981 ( .A(n9480), .B(sreg[1374]), .Z(n724) );
  XOR U982 ( .A(sreg[1374]), .B(n9480), .Z(n725) );
  NANDN U983 ( .A(n9481), .B(n725), .Z(n726) );
  NAND U984 ( .A(n724), .B(n726), .Z(n9503) );
  NAND U985 ( .A(sreg[1378]), .B(n9562), .Z(n727) );
  XOR U986 ( .A(n9562), .B(sreg[1378]), .Z(n728) );
  NANDN U987 ( .A(n9563), .B(n728), .Z(n729) );
  NAND U988 ( .A(n727), .B(n729), .Z(n9583) );
  XOR U989 ( .A(n9647), .B(n9646), .Z(n730) );
  NAND U990 ( .A(n730), .B(sreg[1382]), .Z(n731) );
  NAND U991 ( .A(n9647), .B(n9646), .Z(n732) );
  AND U992 ( .A(n731), .B(n732), .Z(n9649) );
  XOR U993 ( .A(sreg[1389]), .B(n9781), .Z(n733) );
  NANDN U994 ( .A(n9782), .B(n733), .Z(n734) );
  NAND U995 ( .A(sreg[1389]), .B(n9781), .Z(n735) );
  AND U996 ( .A(n734), .B(n735), .Z(n9821) );
  XOR U997 ( .A(n9891), .B(n9890), .Z(n736) );
  NANDN U998 ( .A(sreg[1394]), .B(n736), .Z(n737) );
  NAND U999 ( .A(n9891), .B(n9890), .Z(n738) );
  AND U1000 ( .A(n737), .B(n738), .Z(n9930) );
  NAND U1001 ( .A(sreg[1402]), .B(n10076), .Z(n739) );
  XOR U1002 ( .A(n10076), .B(sreg[1402]), .Z(n740) );
  NANDN U1003 ( .A(n10077), .B(n740), .Z(n741) );
  NAND U1004 ( .A(n739), .B(n741), .Z(n10079) );
  XOR U1005 ( .A(n10167), .B(sreg[1407]), .Z(n742) );
  NANDN U1006 ( .A(n10168), .B(n742), .Z(n743) );
  NAND U1007 ( .A(n10167), .B(sreg[1407]), .Z(n744) );
  AND U1008 ( .A(n743), .B(n744), .Z(n10203) );
  XOR U1009 ( .A(sreg[1413]), .B(n10297), .Z(n745) );
  NANDN U1010 ( .A(n10298), .B(n745), .Z(n746) );
  NAND U1011 ( .A(sreg[1413]), .B(n10297), .Z(n747) );
  AND U1012 ( .A(n746), .B(n747), .Z(n10337) );
  XOR U1013 ( .A(sreg[1422]), .B(n10498), .Z(n748) );
  NANDN U1014 ( .A(n10499), .B(n748), .Z(n749) );
  NAND U1015 ( .A(sreg[1422]), .B(n10498), .Z(n750) );
  AND U1016 ( .A(n749), .B(n750), .Z(n10537) );
  XOR U1017 ( .A(sreg[1427]), .B(n10607), .Z(n751) );
  NANDN U1018 ( .A(n10608), .B(n751), .Z(n752) );
  NAND U1019 ( .A(sreg[1427]), .B(n10607), .Z(n753) );
  AND U1020 ( .A(n752), .B(n753), .Z(n10647) );
  XOR U1021 ( .A(n10719), .B(sreg[1432]), .Z(n754) );
  NAND U1022 ( .A(n754), .B(n10718), .Z(n755) );
  NAND U1023 ( .A(n10719), .B(sreg[1432]), .Z(n756) );
  AND U1024 ( .A(n755), .B(n756), .Z(n10758) );
  XOR U1025 ( .A(sreg[1437]), .B(n10829), .Z(n757) );
  NANDN U1026 ( .A(n10830), .B(n757), .Z(n758) );
  NAND U1027 ( .A(sreg[1437]), .B(n10829), .Z(n759) );
  AND U1028 ( .A(n758), .B(n759), .Z(n10869) );
  XOR U1029 ( .A(sreg[1442]), .B(n10940), .Z(n760) );
  NANDN U1030 ( .A(n10941), .B(n760), .Z(n761) );
  NAND U1031 ( .A(sreg[1442]), .B(n10940), .Z(n762) );
  AND U1032 ( .A(n761), .B(n762), .Z(n10980) );
  NAND U1033 ( .A(n11075), .B(n11074), .Z(n763) );
  XOR U1034 ( .A(n11074), .B(n11075), .Z(n764) );
  NAND U1035 ( .A(n764), .B(sreg[1448]), .Z(n765) );
  NAND U1036 ( .A(n763), .B(n765), .Z(n11113) );
  XOR U1037 ( .A(sreg[1453]), .B(n11185), .Z(n766) );
  NANDN U1038 ( .A(n11186), .B(n766), .Z(n767) );
  NAND U1039 ( .A(sreg[1453]), .B(n11185), .Z(n768) );
  AND U1040 ( .A(n767), .B(n768), .Z(n11225) );
  NAND U1041 ( .A(n11318), .B(n11317), .Z(n769) );
  XOR U1042 ( .A(n11317), .B(n11318), .Z(n770) );
  NANDN U1043 ( .A(sreg[1459]), .B(n770), .Z(n771) );
  NAND U1044 ( .A(n769), .B(n771), .Z(n11356) );
  XOR U1045 ( .A(n11407), .B(sreg[1463]), .Z(n772) );
  NAND U1046 ( .A(n772), .B(n11406), .Z(n773) );
  NAND U1047 ( .A(n11407), .B(sreg[1463]), .Z(n774) );
  AND U1048 ( .A(n773), .B(n774), .Z(n11443) );
  NAND U1049 ( .A(sreg[1471]), .B(n11592), .Z(n775) );
  XOR U1050 ( .A(n11592), .B(sreg[1471]), .Z(n776) );
  NANDN U1051 ( .A(n11593), .B(n776), .Z(n777) );
  NAND U1052 ( .A(n775), .B(n777), .Z(n11595) );
  XOR U1053 ( .A(sreg[1475]), .B(n11657), .Z(n778) );
  NANDN U1054 ( .A(n11658), .B(n778), .Z(n779) );
  NAND U1055 ( .A(sreg[1475]), .B(n11657), .Z(n780) );
  AND U1056 ( .A(n779), .B(n780), .Z(n11697) );
  XOR U1057 ( .A(sreg[1487]), .B(n11927), .Z(n781) );
  NANDN U1058 ( .A(n11928), .B(n781), .Z(n782) );
  NAND U1059 ( .A(sreg[1487]), .B(n11927), .Z(n783) );
  AND U1060 ( .A(n782), .B(n783), .Z(n11967) );
  XOR U1061 ( .A(n12030), .B(n12029), .Z(n784) );
  NANDN U1062 ( .A(sreg[1491]), .B(n784), .Z(n785) );
  NAND U1063 ( .A(n12030), .B(n12029), .Z(n786) );
  AND U1064 ( .A(n785), .B(n786), .Z(n12032) );
  NAND U1065 ( .A(sreg[1496]), .B(n12138), .Z(n787) );
  XOR U1066 ( .A(n12138), .B(sreg[1496]), .Z(n788) );
  NANDN U1067 ( .A(n12139), .B(n788), .Z(n789) );
  NAND U1068 ( .A(n787), .B(n789), .Z(n12141) );
  NAND U1069 ( .A(sreg[1500]), .B(n12227), .Z(n790) );
  XOR U1070 ( .A(n12227), .B(sreg[1500]), .Z(n791) );
  NANDN U1071 ( .A(n12228), .B(n791), .Z(n792) );
  NAND U1072 ( .A(n790), .B(n792), .Z(n12245) );
  NAND U1073 ( .A(sreg[1504]), .B(n12306), .Z(n793) );
  XOR U1074 ( .A(n12306), .B(sreg[1504]), .Z(n794) );
  NANDN U1075 ( .A(n12307), .B(n794), .Z(n795) );
  NAND U1076 ( .A(n793), .B(n795), .Z(n12309) );
  NAND U1077 ( .A(n12377), .B(n12376), .Z(n796) );
  XOR U1078 ( .A(n12376), .B(n12377), .Z(n797) );
  NAND U1079 ( .A(n797), .B(sreg[1508]), .Z(n798) );
  NAND U1080 ( .A(n796), .B(n798), .Z(n12415) );
  NAND U1081 ( .A(n12465), .B(n12464), .Z(n799) );
  XOR U1082 ( .A(n12464), .B(n12465), .Z(n800) );
  NAND U1083 ( .A(n800), .B(sreg[1512]), .Z(n801) );
  NAND U1084 ( .A(n799), .B(n801), .Z(n12503) );
  NAND U1085 ( .A(n12707), .B(sreg[1522]), .Z(n802) );
  XOR U1086 ( .A(sreg[1522]), .B(n12707), .Z(n803) );
  NANDN U1087 ( .A(n12706), .B(n803), .Z(n804) );
  NAND U1088 ( .A(n802), .B(n804), .Z(n12728) );
  XOR U1089 ( .A(sreg[1530]), .B(n12866), .Z(n805) );
  NANDN U1090 ( .A(n12867), .B(n805), .Z(n806) );
  NAND U1091 ( .A(sreg[1530]), .B(n12866), .Z(n807) );
  AND U1092 ( .A(n806), .B(n807), .Z(n12906) );
  XOR U1093 ( .A(n12978), .B(sreg[1535]), .Z(n808) );
  NAND U1094 ( .A(n808), .B(n12977), .Z(n809) );
  NAND U1095 ( .A(n12978), .B(sreg[1535]), .Z(n810) );
  AND U1096 ( .A(n809), .B(n810), .Z(n13013) );
  NAND U1097 ( .A(n13126), .B(n13125), .Z(n811) );
  XOR U1098 ( .A(n13125), .B(n13126), .Z(n812) );
  NAND U1099 ( .A(n812), .B(sreg[1541]), .Z(n813) );
  NAND U1100 ( .A(n811), .B(n813), .Z(n13129) );
  XOR U1101 ( .A(sreg[1545]), .B(n13195), .Z(n814) );
  NANDN U1102 ( .A(n13196), .B(n814), .Z(n815) );
  NAND U1103 ( .A(sreg[1545]), .B(n13195), .Z(n816) );
  AND U1104 ( .A(n815), .B(n816), .Z(n13235) );
  NAND U1105 ( .A(sreg[1550]), .B(n13324), .Z(n817) );
  XOR U1106 ( .A(n13324), .B(sreg[1550]), .Z(n818) );
  NANDN U1107 ( .A(n13325), .B(n818), .Z(n819) );
  NAND U1108 ( .A(n817), .B(n819), .Z(n13345) );
  NAND U1109 ( .A(n13393), .B(sreg[1554]), .Z(n820) );
  XOR U1110 ( .A(sreg[1554]), .B(n13393), .Z(n821) );
  NANDN U1111 ( .A(n13392), .B(n821), .Z(n822) );
  NAND U1112 ( .A(n820), .B(n822), .Z(n13431) );
  NAND U1113 ( .A(sreg[1560]), .B(n13542), .Z(n823) );
  XOR U1114 ( .A(n13542), .B(sreg[1560]), .Z(n824) );
  NANDN U1115 ( .A(n13543), .B(n824), .Z(n825) );
  NAND U1116 ( .A(n823), .B(n825), .Z(n13545) );
  NAND U1117 ( .A(sreg[1574]), .B(n13856), .Z(n826) );
  XOR U1118 ( .A(n13856), .B(sreg[1574]), .Z(n827) );
  NANDN U1119 ( .A(n13857), .B(n827), .Z(n828) );
  NAND U1120 ( .A(n826), .B(n828), .Z(n13859) );
  NAND U1121 ( .A(sreg[1581]), .B(n14013), .Z(n829) );
  XOR U1122 ( .A(n14013), .B(sreg[1581]), .Z(n830) );
  NANDN U1123 ( .A(n14014), .B(n830), .Z(n831) );
  NAND U1124 ( .A(n829), .B(n831), .Z(n14016) );
  NAND U1125 ( .A(n14098), .B(n14097), .Z(n832) );
  XOR U1126 ( .A(n14097), .B(n14098), .Z(n833) );
  NANDN U1127 ( .A(sreg[1585]), .B(n833), .Z(n834) );
  NAND U1128 ( .A(n832), .B(n834), .Z(n14100) );
  XOR U1129 ( .A(n14166), .B(sreg[1589]), .Z(n835) );
  NAND U1130 ( .A(n835), .B(n14165), .Z(n836) );
  NAND U1131 ( .A(n14166), .B(sreg[1589]), .Z(n837) );
  AND U1132 ( .A(n836), .B(n837), .Z(n14205) );
  XOR U1133 ( .A(sreg[1593]), .B(n14253), .Z(n838) );
  NANDN U1134 ( .A(n14254), .B(n838), .Z(n839) );
  NAND U1135 ( .A(sreg[1593]), .B(n14253), .Z(n840) );
  AND U1136 ( .A(n839), .B(n840), .Z(n14293) );
  NAND U1137 ( .A(n14365), .B(sreg[1598]), .Z(n841) );
  XOR U1138 ( .A(sreg[1598]), .B(n14365), .Z(n842) );
  NANDN U1139 ( .A(n14364), .B(n842), .Z(n843) );
  NAND U1140 ( .A(n841), .B(n843), .Z(n14403) );
  NAND U1141 ( .A(n14451), .B(n14450), .Z(n844) );
  XOR U1142 ( .A(n14450), .B(n14451), .Z(n845) );
  NAND U1143 ( .A(n845), .B(sreg[1602]), .Z(n846) );
  NAND U1144 ( .A(n844), .B(n846), .Z(n14489) );
  NAND U1145 ( .A(n14582), .B(sreg[1608]), .Z(n847) );
  XOR U1146 ( .A(sreg[1608]), .B(n14582), .Z(n848) );
  NANDN U1147 ( .A(n14583), .B(n848), .Z(n849) );
  NAND U1148 ( .A(n847), .B(n849), .Z(n14603) );
  XOR U1149 ( .A(n14715), .B(sreg[1614]), .Z(n850) );
  NAND U1150 ( .A(n850), .B(n14714), .Z(n851) );
  NAND U1151 ( .A(n14715), .B(sreg[1614]), .Z(n852) );
  AND U1152 ( .A(n851), .B(n852), .Z(n14736) );
  XOR U1153 ( .A(sreg[1618]), .B(n14802), .Z(n853) );
  NANDN U1154 ( .A(n14803), .B(n853), .Z(n854) );
  NAND U1155 ( .A(sreg[1618]), .B(n14802), .Z(n855) );
  AND U1156 ( .A(n854), .B(n855), .Z(n14823) );
  XOR U1157 ( .A(sreg[1622]), .B(n14888), .Z(n856) );
  NANDN U1158 ( .A(n14889), .B(n856), .Z(n857) );
  NAND U1159 ( .A(sreg[1622]), .B(n14888), .Z(n858) );
  AND U1160 ( .A(n857), .B(n858), .Z(n14928) );
  NAND U1161 ( .A(n14975), .B(n14974), .Z(n859) );
  XOR U1162 ( .A(n14974), .B(n14975), .Z(n860) );
  NAND U1163 ( .A(n860), .B(sreg[1626]), .Z(n861) );
  NAND U1164 ( .A(n859), .B(n861), .Z(n15013) );
  NAND U1165 ( .A(sreg[1630]), .B(n15080), .Z(n862) );
  XOR U1166 ( .A(n15080), .B(sreg[1630]), .Z(n863) );
  NANDN U1167 ( .A(n15081), .B(n863), .Z(n864) );
  NAND U1168 ( .A(n862), .B(n864), .Z(n15101) );
  NAND U1169 ( .A(n15149), .B(sreg[1634]), .Z(n865) );
  XOR U1170 ( .A(sreg[1634]), .B(n15149), .Z(n866) );
  NANDN U1171 ( .A(n15148), .B(n866), .Z(n867) );
  NAND U1172 ( .A(n865), .B(n867), .Z(n15187) );
  NAND U1173 ( .A(sreg[1642]), .B(n15346), .Z(n868) );
  XOR U1174 ( .A(n15346), .B(sreg[1642]), .Z(n869) );
  NANDN U1175 ( .A(n15347), .B(n869), .Z(n870) );
  NAND U1176 ( .A(n868), .B(n870), .Z(n15349) );
  NAND U1177 ( .A(n15433), .B(sreg[1646]), .Z(n871) );
  XOR U1178 ( .A(sreg[1646]), .B(n15433), .Z(n872) );
  NAND U1179 ( .A(n872), .B(n15432), .Z(n873) );
  NAND U1180 ( .A(n871), .B(n873), .Z(n15435) );
  NAND U1181 ( .A(n15501), .B(n15500), .Z(n874) );
  XOR U1182 ( .A(n15500), .B(n15501), .Z(n875) );
  NAND U1183 ( .A(n875), .B(sreg[1650]), .Z(n876) );
  NAND U1184 ( .A(n874), .B(n876), .Z(n15539) );
  XOR U1185 ( .A(n15672), .B(n15671), .Z(n877) );
  NANDN U1186 ( .A(sreg[1657]), .B(n877), .Z(n878) );
  NAND U1187 ( .A(n15672), .B(n15671), .Z(n879) );
  AND U1188 ( .A(n878), .B(n879), .Z(n15674) );
  XOR U1189 ( .A(sreg[1661]), .B(n15741), .Z(n880) );
  NANDN U1190 ( .A(n15742), .B(n880), .Z(n881) );
  NAND U1191 ( .A(sreg[1661]), .B(n15741), .Z(n882) );
  AND U1192 ( .A(n881), .B(n882), .Z(n15781) );
  XOR U1193 ( .A(n15853), .B(sreg[1666]), .Z(n883) );
  NAND U1194 ( .A(n883), .B(n15852), .Z(n884) );
  NAND U1195 ( .A(n15853), .B(sreg[1666]), .Z(n885) );
  AND U1196 ( .A(n884), .B(n885), .Z(n15892) );
  XOR U1197 ( .A(sreg[1671]), .B(n15963), .Z(n886) );
  NANDN U1198 ( .A(n15964), .B(n886), .Z(n887) );
  NAND U1199 ( .A(sreg[1671]), .B(n15963), .Z(n888) );
  AND U1200 ( .A(n887), .B(n888), .Z(n16003) );
  NAND U1201 ( .A(n16090), .B(n16089), .Z(n889) );
  XOR U1202 ( .A(n16089), .B(n16090), .Z(n890) );
  NANDN U1203 ( .A(sreg[1676]), .B(n890), .Z(n891) );
  NAND U1204 ( .A(n889), .B(n891), .Z(n16107) );
  XOR U1205 ( .A(sreg[1680]), .B(n16155), .Z(n892) );
  NANDN U1206 ( .A(n16156), .B(n892), .Z(n893) );
  NAND U1207 ( .A(sreg[1680]), .B(n16155), .Z(n894) );
  AND U1208 ( .A(n893), .B(n894), .Z(n16190) );
  NAND U1209 ( .A(n16299), .B(n16298), .Z(n895) );
  XOR U1210 ( .A(n16298), .B(n16299), .Z(n896) );
  NAND U1211 ( .A(n896), .B(sreg[1686]), .Z(n897) );
  NAND U1212 ( .A(n895), .B(n897), .Z(n16301) );
  NAND U1213 ( .A(sreg[1690]), .B(n16386), .Z(n898) );
  XOR U1214 ( .A(n16386), .B(sreg[1690]), .Z(n899) );
  NANDN U1215 ( .A(n16387), .B(n899), .Z(n900) );
  NAND U1216 ( .A(n898), .B(n900), .Z(n16389) );
  NAND U1217 ( .A(n16457), .B(n16456), .Z(n901) );
  XOR U1218 ( .A(n16456), .B(n16457), .Z(n902) );
  NAND U1219 ( .A(n902), .B(sreg[1694]), .Z(n903) );
  NAND U1220 ( .A(n901), .B(n903), .Z(n16495) );
  NAND U1221 ( .A(n16545), .B(n16544), .Z(n904) );
  XOR U1222 ( .A(n16544), .B(n16545), .Z(n905) );
  NAND U1223 ( .A(n905), .B(sreg[1698]), .Z(n906) );
  NAND U1224 ( .A(n904), .B(n906), .Z(n16583) );
  NAND U1225 ( .A(n16654), .B(n16653), .Z(n907) );
  XOR U1226 ( .A(n16653), .B(n16654), .Z(n908) );
  NAND U1227 ( .A(n908), .B(sreg[1703]), .Z(n909) );
  NAND U1228 ( .A(n907), .B(n909), .Z(n16692) );
  NAND U1229 ( .A(n16802), .B(sreg[1709]), .Z(n910) );
  XOR U1230 ( .A(sreg[1709]), .B(n16802), .Z(n911) );
  NAND U1231 ( .A(n911), .B(n16801), .Z(n912) );
  NAND U1232 ( .A(n910), .B(n912), .Z(n16822) );
  NAND U1233 ( .A(sreg[1713]), .B(n16883), .Z(n913) );
  XOR U1234 ( .A(n16883), .B(sreg[1713]), .Z(n914) );
  NANDN U1235 ( .A(n16884), .B(n914), .Z(n915) );
  NAND U1236 ( .A(n913), .B(n915), .Z(n16886) );
  NAND U1237 ( .A(sreg[1718]), .B(n16992), .Z(n916) );
  XOR U1238 ( .A(n16992), .B(sreg[1718]), .Z(n917) );
  NANDN U1239 ( .A(n16993), .B(n917), .Z(n918) );
  NAND U1240 ( .A(n916), .B(n918), .Z(n17013) );
  NAND U1241 ( .A(sreg[1722]), .B(n17078), .Z(n919) );
  XOR U1242 ( .A(n17078), .B(sreg[1722]), .Z(n920) );
  NANDN U1243 ( .A(n17079), .B(n920), .Z(n921) );
  NAND U1244 ( .A(n919), .B(n921), .Z(n17081) );
  NAND U1245 ( .A(n17172), .B(n17171), .Z(n922) );
  XOR U1246 ( .A(n17171), .B(n17172), .Z(n923) );
  NAND U1247 ( .A(n923), .B(sreg[1727]), .Z(n924) );
  NAND U1248 ( .A(n922), .B(n924), .Z(n17193) );
  XOR U1249 ( .A(sreg[1732]), .B(n17278), .Z(n925) );
  NANDN U1250 ( .A(n17279), .B(n925), .Z(n926) );
  NAND U1251 ( .A(sreg[1732]), .B(n17278), .Z(n927) );
  AND U1252 ( .A(n926), .B(n927), .Z(n17318) );
  XOR U1253 ( .A(n17383), .B(n17382), .Z(n928) );
  NANDN U1254 ( .A(sreg[1736]), .B(n928), .Z(n929) );
  NAND U1255 ( .A(n17383), .B(n17382), .Z(n930) );
  AND U1256 ( .A(n929), .B(n930), .Z(n17403) );
  XOR U1257 ( .A(sreg[1740]), .B(n17450), .Z(n931) );
  NANDN U1258 ( .A(n17451), .B(n931), .Z(n932) );
  NAND U1259 ( .A(sreg[1740]), .B(n17450), .Z(n933) );
  AND U1260 ( .A(n932), .B(n933), .Z(n17491) );
  XOR U1261 ( .A(sreg[1752]), .B(n17718), .Z(n934) );
  NANDN U1262 ( .A(n17719), .B(n934), .Z(n935) );
  NAND U1263 ( .A(sreg[1752]), .B(n17718), .Z(n936) );
  AND U1264 ( .A(n935), .B(n936), .Z(n17758) );
  NAND U1265 ( .A(n17966), .B(sreg[1763]), .Z(n937) );
  XOR U1266 ( .A(sreg[1763]), .B(n17966), .Z(n938) );
  NANDN U1267 ( .A(n17965), .B(n938), .Z(n939) );
  NAND U1268 ( .A(n937), .B(n939), .Z(n18004) );
  NAND U1269 ( .A(sreg[1768]), .B(n18092), .Z(n940) );
  XOR U1270 ( .A(n18092), .B(sreg[1768]), .Z(n941) );
  NANDN U1271 ( .A(n18093), .B(n941), .Z(n942) );
  NAND U1272 ( .A(n940), .B(n942), .Z(n18095) );
  XOR U1273 ( .A(sreg[1772]), .B(n18162), .Z(n943) );
  NANDN U1274 ( .A(n18163), .B(n943), .Z(n944) );
  NAND U1275 ( .A(sreg[1772]), .B(n18162), .Z(n945) );
  AND U1276 ( .A(n944), .B(n945), .Z(n18202) );
  XOR U1277 ( .A(sreg[1776]), .B(n18250), .Z(n946) );
  NANDN U1278 ( .A(n18251), .B(n946), .Z(n947) );
  NAND U1279 ( .A(sreg[1776]), .B(n18250), .Z(n948) );
  AND U1280 ( .A(n947), .B(n948), .Z(n18290) );
  NAND U1281 ( .A(n18448), .B(n18447), .Z(n949) );
  XOR U1282 ( .A(n18447), .B(n18448), .Z(n950) );
  NAND U1283 ( .A(n950), .B(sreg[1785]), .Z(n951) );
  NAND U1284 ( .A(n949), .B(n951), .Z(n18486) );
  XOR U1285 ( .A(sreg[1792]), .B(n18599), .Z(n952) );
  NANDN U1286 ( .A(n18600), .B(n952), .Z(n953) );
  NAND U1287 ( .A(sreg[1792]), .B(n18599), .Z(n954) );
  AND U1288 ( .A(n953), .B(n954), .Z(n18616) );
  NAND U1289 ( .A(n18750), .B(n18749), .Z(n955) );
  XOR U1290 ( .A(n18749), .B(n18750), .Z(n956) );
  NAND U1291 ( .A(n956), .B(sreg[1799]), .Z(n957) );
  NAND U1292 ( .A(n955), .B(n957), .Z(n18771) );
  NAND U1293 ( .A(n18838), .B(sreg[1803]), .Z(n958) );
  XOR U1294 ( .A(sreg[1803]), .B(n18838), .Z(n959) );
  NANDN U1295 ( .A(n18837), .B(n959), .Z(n960) );
  NAND U1296 ( .A(n958), .B(n960), .Z(n18876) );
  XOR U1297 ( .A(n19032), .B(n19031), .Z(n961) );
  NANDN U1298 ( .A(sreg[1811]), .B(n961), .Z(n962) );
  NAND U1299 ( .A(n19032), .B(n19031), .Z(n963) );
  AND U1300 ( .A(n962), .B(n963), .Z(n19034) );
  NAND U1301 ( .A(n19167), .B(n19166), .Z(n964) );
  XOR U1302 ( .A(n19166), .B(n19167), .Z(n965) );
  NAND U1303 ( .A(n965), .B(sreg[1818]), .Z(n966) );
  NAND U1304 ( .A(n964), .B(n966), .Z(n19205) );
  XOR U1305 ( .A(n19274), .B(sreg[1823]), .Z(n967) );
  NAND U1306 ( .A(n967), .B(n19273), .Z(n968) );
  NAND U1307 ( .A(n19274), .B(sreg[1823]), .Z(n969) );
  AND U1308 ( .A(n968), .B(n969), .Z(n19310) );
  NAND U1309 ( .A(n19418), .B(sreg[1829]), .Z(n970) );
  XOR U1310 ( .A(sreg[1829]), .B(n19418), .Z(n971) );
  NAND U1311 ( .A(n971), .B(n19417), .Z(n972) );
  NAND U1312 ( .A(n970), .B(n972), .Z(n19420) );
  XOR U1313 ( .A(n19525), .B(n19524), .Z(n973) );
  NANDN U1314 ( .A(sreg[1834]), .B(n973), .Z(n974) );
  NAND U1315 ( .A(n19525), .B(n19524), .Z(n975) );
  AND U1316 ( .A(n974), .B(n975), .Z(n19527) );
  XOR U1317 ( .A(sreg[1838]), .B(n19592), .Z(n976) );
  NANDN U1318 ( .A(n19593), .B(n976), .Z(n977) );
  NAND U1319 ( .A(sreg[1838]), .B(n19592), .Z(n978) );
  AND U1320 ( .A(n977), .B(n978), .Z(n19632) );
  NAND U1321 ( .A(n19746), .B(n19745), .Z(n979) );
  XOR U1322 ( .A(n19745), .B(n19746), .Z(n980) );
  NAND U1323 ( .A(n980), .B(sreg[1845]), .Z(n981) );
  NAND U1324 ( .A(n979), .B(n981), .Z(n19766) );
  XOR U1325 ( .A(sreg[1850]), .B(n19854), .Z(n982) );
  NANDN U1326 ( .A(n19855), .B(n982), .Z(n983) );
  NAND U1327 ( .A(sreg[1850]), .B(n19854), .Z(n984) );
  AND U1328 ( .A(n983), .B(n984), .Z(n19894) );
  XOR U1329 ( .A(n20028), .B(n20027), .Z(n985) );
  NANDN U1330 ( .A(sreg[1857]), .B(n985), .Z(n986) );
  NAND U1331 ( .A(n20028), .B(n20027), .Z(n987) );
  AND U1332 ( .A(n986), .B(n987), .Z(n20030) );
  NAND U1333 ( .A(n20098), .B(n20097), .Z(n988) );
  XOR U1334 ( .A(n20097), .B(n20098), .Z(n989) );
  NAND U1335 ( .A(n989), .B(sreg[1861]), .Z(n990) );
  NAND U1336 ( .A(n988), .B(n990), .Z(n20136) );
  XOR U1337 ( .A(n20186), .B(sreg[1865]), .Z(n991) );
  NAND U1338 ( .A(n991), .B(n20185), .Z(n992) );
  NAND U1339 ( .A(n20186), .B(sreg[1865]), .Z(n993) );
  AND U1340 ( .A(n992), .B(n993), .Z(n20224) );
  NAND U1341 ( .A(n20294), .B(sreg[1870]), .Z(n994) );
  XOR U1342 ( .A(sreg[1870]), .B(n20294), .Z(n995) );
  NANDN U1343 ( .A(n20295), .B(n995), .Z(n996) );
  NAND U1344 ( .A(n994), .B(n996), .Z(n20333) );
  NAND U1345 ( .A(n20406), .B(n20405), .Z(n997) );
  XOR U1346 ( .A(n20405), .B(n20406), .Z(n998) );
  NAND U1347 ( .A(n998), .B(sreg[1875]), .Z(n999) );
  NAND U1348 ( .A(n997), .B(n999), .Z(n20444) );
  NAND U1349 ( .A(n20493), .B(sreg[1879]), .Z(n1000) );
  XOR U1350 ( .A(sreg[1879]), .B(n20493), .Z(n1001) );
  NANDN U1351 ( .A(n20494), .B(n1001), .Z(n1002) );
  NAND U1352 ( .A(n1000), .B(n1002), .Z(n20532) );
  XOR U1353 ( .A(sreg[1884]), .B(n20600), .Z(n1003) );
  NANDN U1354 ( .A(n20601), .B(n1003), .Z(n1004) );
  NAND U1355 ( .A(sreg[1884]), .B(n20600), .Z(n1005) );
  AND U1356 ( .A(n1004), .B(n1005), .Z(n20638) );
  NAND U1357 ( .A(n20685), .B(sreg[1888]), .Z(n1006) );
  XOR U1358 ( .A(sreg[1888]), .B(n20685), .Z(n1007) );
  NANDN U1359 ( .A(n20686), .B(n1007), .Z(n1008) );
  NAND U1360 ( .A(n1006), .B(n1008), .Z(n20719) );
  NAND U1361 ( .A(n20831), .B(n20830), .Z(n1009) );
  XOR U1362 ( .A(n20830), .B(n20831), .Z(n1010) );
  NAND U1363 ( .A(n1010), .B(sreg[1894]), .Z(n1011) );
  NAND U1364 ( .A(n1009), .B(n1011), .Z(n20833) );
  XOR U1365 ( .A(sreg[1898]), .B(n20898), .Z(n1012) );
  NANDN U1366 ( .A(n20899), .B(n1012), .Z(n1013) );
  NAND U1367 ( .A(sreg[1898]), .B(n20898), .Z(n1014) );
  AND U1368 ( .A(n1013), .B(n1014), .Z(n20938) );
  XOR U1369 ( .A(sreg[1902]), .B(n20986), .Z(n1015) );
  NANDN U1370 ( .A(n20987), .B(n1015), .Z(n1016) );
  NAND U1371 ( .A(sreg[1902]), .B(n20986), .Z(n1017) );
  AND U1372 ( .A(n1016), .B(n1017), .Z(n21026) );
  NAND U1373 ( .A(sreg[1908]), .B(n21136), .Z(n1018) );
  XOR U1374 ( .A(n21136), .B(sreg[1908]), .Z(n1019) );
  NANDN U1375 ( .A(n21137), .B(n1019), .Z(n1020) );
  NAND U1376 ( .A(n1018), .B(n1020), .Z(n21139) );
  NAND U1377 ( .A(n21205), .B(n21204), .Z(n1021) );
  XOR U1378 ( .A(n21204), .B(n21205), .Z(n1022) );
  NAND U1379 ( .A(n1022), .B(sreg[1912]), .Z(n1023) );
  NAND U1380 ( .A(n1021), .B(n1023), .Z(n21225) );
  XOR U1381 ( .A(sreg[1916]), .B(n21290), .Z(n1024) );
  NANDN U1382 ( .A(n21291), .B(n1024), .Z(n1025) );
  NAND U1383 ( .A(sreg[1916]), .B(n21290), .Z(n1026) );
  AND U1384 ( .A(n1025), .B(n1026), .Z(n21330) );
  NAND U1385 ( .A(sreg[1921]), .B(n21419), .Z(n1027) );
  XOR U1386 ( .A(n21419), .B(sreg[1921]), .Z(n1028) );
  NANDN U1387 ( .A(n21420), .B(n1028), .Z(n1029) );
  NAND U1388 ( .A(n1027), .B(n1029), .Z(n21440) );
  NAND U1389 ( .A(n21506), .B(sreg[1925]), .Z(n1030) );
  XOR U1390 ( .A(sreg[1925]), .B(n21506), .Z(n1031) );
  NANDN U1391 ( .A(n21505), .B(n1031), .Z(n1032) );
  NAND U1392 ( .A(n1030), .B(n1032), .Z(n21526) );
  NAND U1393 ( .A(n21571), .B(sreg[1929]), .Z(n1033) );
  XOR U1394 ( .A(sreg[1929]), .B(n21571), .Z(n1034) );
  NANDN U1395 ( .A(n21572), .B(n1034), .Z(n1035) );
  NAND U1396 ( .A(n1033), .B(n1035), .Z(n21610) );
  XOR U1397 ( .A(sreg[1939]), .B(n21793), .Z(n1036) );
  NANDN U1398 ( .A(n21794), .B(n1036), .Z(n1037) );
  NAND U1399 ( .A(sreg[1939]), .B(n21793), .Z(n1038) );
  AND U1400 ( .A(n1037), .B(n1038), .Z(n21832) );
  NAND U1401 ( .A(n21882), .B(n21881), .Z(n1039) );
  XOR U1402 ( .A(n21881), .B(n21882), .Z(n1040) );
  NAND U1403 ( .A(n1040), .B(sreg[1943]), .Z(n1041) );
  NAND U1404 ( .A(n1039), .B(n1041), .Z(n21903) );
  NAND U1405 ( .A(n22033), .B(sreg[1949]), .Z(n1042) );
  XOR U1406 ( .A(sreg[1949]), .B(n22033), .Z(n1043) );
  NANDN U1407 ( .A(n22032), .B(n1043), .Z(n1044) );
  NAND U1408 ( .A(n1042), .B(n1044), .Z(n22035) );
  XOR U1409 ( .A(n22101), .B(n22100), .Z(n1045) );
  NANDN U1410 ( .A(sreg[1953]), .B(n1045), .Z(n1046) );
  NAND U1411 ( .A(n22101), .B(n22100), .Z(n1047) );
  AND U1412 ( .A(n1046), .B(n1047), .Z(n22134) );
  NAND U1413 ( .A(sreg[1961]), .B(n22291), .Z(n1048) );
  XOR U1414 ( .A(n22291), .B(sreg[1961]), .Z(n1049) );
  NANDN U1415 ( .A(n22292), .B(n1049), .Z(n1050) );
  NAND U1416 ( .A(n1048), .B(n1050), .Z(n22294) );
  NAND U1417 ( .A(n22475), .B(sreg[1970]), .Z(n1051) );
  XOR U1418 ( .A(sreg[1970]), .B(n22475), .Z(n1052) );
  NAND U1419 ( .A(n1052), .B(n22474), .Z(n1053) );
  NAND U1420 ( .A(n1051), .B(n1053), .Z(n22513) );
  XOR U1421 ( .A(sreg[1975]), .B(n22585), .Z(n1054) );
  NANDN U1422 ( .A(n22586), .B(n1054), .Z(n1055) );
  NAND U1423 ( .A(sreg[1975]), .B(n22585), .Z(n1056) );
  AND U1424 ( .A(n1055), .B(n1056), .Z(n22624) );
  XOR U1425 ( .A(sreg[1980]), .B(n22696), .Z(n1057) );
  NANDN U1426 ( .A(n22697), .B(n1057), .Z(n1058) );
  NAND U1427 ( .A(sreg[1980]), .B(n22696), .Z(n1059) );
  AND U1428 ( .A(n1058), .B(n1059), .Z(n22736) );
  NAND U1429 ( .A(n22785), .B(sreg[1984]), .Z(n1060) );
  XOR U1430 ( .A(sreg[1984]), .B(n22785), .Z(n1061) );
  NANDN U1431 ( .A(n22784), .B(n1061), .Z(n1062) );
  NAND U1432 ( .A(n1060), .B(n1062), .Z(n22823) );
  NAND U1433 ( .A(n22958), .B(sreg[1992]), .Z(n1063) );
  XOR U1434 ( .A(sreg[1992]), .B(n22958), .Z(n1064) );
  NANDN U1435 ( .A(n22959), .B(n1064), .Z(n1065) );
  NAND U1436 ( .A(n1063), .B(n1065), .Z(n22979) );
  NAND U1437 ( .A(sreg[1997]), .B(n23085), .Z(n1066) );
  XOR U1438 ( .A(n23085), .B(sreg[1997]), .Z(n1067) );
  NANDN U1439 ( .A(n23086), .B(n1067), .Z(n1068) );
  NAND U1440 ( .A(n1066), .B(n1068), .Z(n23088) );
  NAND U1441 ( .A(n23170), .B(n23169), .Z(n1069) );
  XOR U1442 ( .A(n23169), .B(n23170), .Z(n1070) );
  NANDN U1443 ( .A(sreg[2001]), .B(n1070), .Z(n1071) );
  NAND U1444 ( .A(n1069), .B(n1071), .Z(n23172) );
  NAND U1445 ( .A(n23238), .B(n23237), .Z(n1072) );
  XOR U1446 ( .A(n23237), .B(n23238), .Z(n1073) );
  NAND U1447 ( .A(n1073), .B(sreg[2005]), .Z(n1074) );
  NAND U1448 ( .A(n1072), .B(n1074), .Z(n23276) );
  XOR U1449 ( .A(sreg[2010]), .B(n23348), .Z(n1075) );
  NANDN U1450 ( .A(n23349), .B(n1075), .Z(n1076) );
  NAND U1451 ( .A(sreg[2010]), .B(n23348), .Z(n1077) );
  AND U1452 ( .A(n1076), .B(n1077), .Z(n23388) );
  NAND U1453 ( .A(n23437), .B(n23436), .Z(n1078) );
  XOR U1454 ( .A(n23436), .B(n23437), .Z(n1079) );
  NAND U1455 ( .A(n1079), .B(sreg[2014]), .Z(n1080) );
  NAND U1456 ( .A(n1078), .B(n1080), .Z(n23475) );
  NAND U1457 ( .A(n23525), .B(n23524), .Z(n1081) );
  XOR U1458 ( .A(n23524), .B(n23525), .Z(n1082) );
  NAND U1459 ( .A(n1082), .B(sreg[2018]), .Z(n1083) );
  NAND U1460 ( .A(n1081), .B(n1083), .Z(n23563) );
  XOR U1461 ( .A(sreg[2022]), .B(n23610), .Z(n1084) );
  NANDN U1462 ( .A(n23611), .B(n1084), .Z(n1085) );
  NAND U1463 ( .A(sreg[2022]), .B(n23610), .Z(n1086) );
  AND U1464 ( .A(n1085), .B(n1086), .Z(n23650) );
  XOR U1465 ( .A(sreg[2026]), .B(n23696), .Z(n1087) );
  NANDN U1466 ( .A(n23697), .B(n1087), .Z(n1088) );
  NAND U1467 ( .A(sreg[2026]), .B(n23696), .Z(n1089) );
  AND U1468 ( .A(n1088), .B(n1089), .Z(n23736) );
  NAND U1469 ( .A(n23808), .B(sreg[2031]), .Z(n1090) );
  XOR U1470 ( .A(sreg[2031]), .B(n23808), .Z(n1091) );
  NANDN U1471 ( .A(n23807), .B(n1091), .Z(n1092) );
  NAND U1472 ( .A(n1090), .B(n1092), .Z(n23846) );
  NAND U1473 ( .A(n23965), .B(n23964), .Z(n1093) );
  XOR U1474 ( .A(n23964), .B(n23965), .Z(n1094) );
  NAND U1475 ( .A(n1094), .B(sreg[2038]), .Z(n1095) );
  NAND U1476 ( .A(n1093), .B(n1095), .Z(n23985) );
  NAND U1477 ( .A(b[2]), .B(a[2]), .Z(n1846) );
  XOR U1478 ( .A(n1867), .B(n1868), .Z(n1869) );
  NANDN U1479 ( .A(n11483), .B(n11482), .Z(n1096) );
  NANDN U1480 ( .A(n11484), .B(n11485), .Z(n1097) );
  NAND U1481 ( .A(n1096), .B(n1097), .Z(n11487) );
  NANDN U1482 ( .A(n11601), .B(n11600), .Z(n1098) );
  NANDN U1483 ( .A(n11602), .B(n11603), .Z(n1099) );
  NAND U1484 ( .A(n1098), .B(n1099), .Z(n11622) );
  NANDN U1485 ( .A(n3939), .B(n3938), .Z(n1100) );
  NANDN U1486 ( .A(n3940), .B(n3941), .Z(n1101) );
  NAND U1487 ( .A(n1100), .B(n1101), .Z(n3943) );
  NANDN U1488 ( .A(n6644), .B(n6643), .Z(n1102) );
  NANDN U1489 ( .A(n6645), .B(n6646), .Z(n1103) );
  NAND U1490 ( .A(n1102), .B(n1103), .Z(n6648) );
  NAND U1491 ( .A(n9509), .B(n9508), .Z(n1104) );
  XOR U1492 ( .A(n9508), .B(n9509), .Z(n1105) );
  NAND U1493 ( .A(n1105), .B(n9507), .Z(n1106) );
  NAND U1494 ( .A(n1104), .B(n1106), .Z(n9522) );
  NAND U1495 ( .A(n9999), .B(n9997), .Z(n1107) );
  XOR U1496 ( .A(n9997), .B(n9999), .Z(n1108) );
  NANDN U1497 ( .A(n9998), .B(n1108), .Z(n1109) );
  NAND U1498 ( .A(n1107), .B(n1109), .Z(n10020) );
  XOR U1499 ( .A(n10125), .B(n10124), .Z(n1110) );
  NANDN U1500 ( .A(n10123), .B(n1110), .Z(n1111) );
  NAND U1501 ( .A(n10125), .B(n10124), .Z(n1112) );
  AND U1502 ( .A(n1111), .B(n1112), .Z(n10146) );
  NAND U1503 ( .A(n11410), .B(n11408), .Z(n1113) );
  XOR U1504 ( .A(n11408), .B(n11410), .Z(n1114) );
  NANDN U1505 ( .A(n11409), .B(n1114), .Z(n1115) );
  NAND U1506 ( .A(n1113), .B(n1115), .Z(n11426) );
  NANDN U1507 ( .A(n16043), .B(n16042), .Z(n1116) );
  NANDN U1508 ( .A(n16044), .B(n16045), .Z(n1117) );
  NAND U1509 ( .A(n1116), .B(n1117), .Z(n16059) );
  NAND U1510 ( .A(n18602), .B(n18601), .Z(n1118) );
  XOR U1511 ( .A(n18601), .B(n18602), .Z(n1119) );
  NANDN U1512 ( .A(n18603), .B(n1119), .Z(n1120) );
  NAND U1513 ( .A(n1118), .B(n1120), .Z(n18634) );
  NANDN U1514 ( .A(n20573), .B(n20572), .Z(n1121) );
  NANDN U1515 ( .A(n20574), .B(n20575), .Z(n1122) );
  NAND U1516 ( .A(n1121), .B(n1122), .Z(n20577) );
  NAND U1517 ( .A(n21684), .B(n21682), .Z(n1123) );
  XOR U1518 ( .A(n21682), .B(n21684), .Z(n1124) );
  NANDN U1519 ( .A(n21683), .B(n1124), .Z(n1125) );
  NAND U1520 ( .A(n1123), .B(n1125), .Z(n21705) );
  NAND U1521 ( .A(n22104), .B(n22103), .Z(n1126) );
  XOR U1522 ( .A(n22103), .B(n22104), .Z(n1127) );
  NAND U1523 ( .A(n1127), .B(n22102), .Z(n1128) );
  NAND U1524 ( .A(n1126), .B(n1128), .Z(n22117) );
  NANDN U1525 ( .A(n24086), .B(n24087), .Z(n1129) );
  NANDN U1526 ( .A(n24085), .B(n24084), .Z(n1130) );
  AND U1527 ( .A(n1129), .B(n1130), .Z(n24090) );
  NAND U1528 ( .A(sreg[1022]), .B(n1814), .Z(n1131) );
  XOR U1529 ( .A(n1814), .B(sreg[1022]), .Z(n1132) );
  NANDN U1530 ( .A(n1815), .B(n1132), .Z(n1133) );
  NAND U1531 ( .A(n1131), .B(n1133), .Z(n1832) );
  NAND U1532 ( .A(n3237), .B(n3236), .Z(n1134) );
  XOR U1533 ( .A(n3236), .B(n3237), .Z(n1135) );
  NANDN U1534 ( .A(n3238), .B(n1135), .Z(n1136) );
  NAND U1535 ( .A(n1134), .B(n1136), .Z(n3257) );
  NAND U1536 ( .A(n5708), .B(n5707), .Z(n1137) );
  XOR U1537 ( .A(n5707), .B(n5708), .Z(n1138) );
  NANDN U1538 ( .A(n5709), .B(n1138), .Z(n1139) );
  NAND U1539 ( .A(n1137), .B(n1139), .Z(n5730) );
  XOR U1540 ( .A(n6573), .B(n6572), .Z(n1140) );
  NANDN U1541 ( .A(n6571), .B(n1140), .Z(n1141) );
  NAND U1542 ( .A(n6573), .B(n6572), .Z(n1142) );
  AND U1543 ( .A(n1141), .B(n1142), .Z(n6592) );
  XOR U1544 ( .A(n7025), .B(n7024), .Z(n1143) );
  NANDN U1545 ( .A(n7023), .B(n1143), .Z(n1144) );
  NAND U1546 ( .A(n7025), .B(n7024), .Z(n1145) );
  AND U1547 ( .A(n1144), .B(n1145), .Z(n7049) );
  NAND U1548 ( .A(n7779), .B(n7778), .Z(n1146) );
  XOR U1549 ( .A(n7778), .B(n7779), .Z(n1147) );
  NANDN U1550 ( .A(n7780), .B(n1147), .Z(n1148) );
  NAND U1551 ( .A(n1146), .B(n1148), .Z(n7799) );
  NAND U1552 ( .A(n8483), .B(n8482), .Z(n1149) );
  XOR U1553 ( .A(n8482), .B(n8483), .Z(n1150) );
  NAND U1554 ( .A(n1150), .B(n8481), .Z(n1151) );
  NAND U1555 ( .A(n1149), .B(n1151), .Z(n8502) );
  NAND U1556 ( .A(n9871), .B(n9869), .Z(n1152) );
  XOR U1557 ( .A(n9869), .B(n9871), .Z(n1153) );
  NANDN U1558 ( .A(n9870), .B(n1153), .Z(n1154) );
  NAND U1559 ( .A(n1152), .B(n1154), .Z(n9895) );
  NAND U1560 ( .A(n11536), .B(n11534), .Z(n1155) );
  XOR U1561 ( .A(n11534), .B(n11536), .Z(n1156) );
  NANDN U1562 ( .A(n11535), .B(n1156), .Z(n1157) );
  NAND U1563 ( .A(n1155), .B(n1157), .Z(n11555) );
  NAND U1564 ( .A(n19254), .B(n19252), .Z(n1158) );
  XOR U1565 ( .A(n19252), .B(n19254), .Z(n1159) );
  NANDN U1566 ( .A(n19253), .B(n1159), .Z(n1160) );
  NAND U1567 ( .A(n1158), .B(n1160), .Z(n19278) );
  NANDN U1568 ( .A(n24055), .B(n24056), .Z(n1161) );
  NANDN U1569 ( .A(n24053), .B(n24054), .Z(n1162) );
  NAND U1570 ( .A(n1161), .B(n1162), .Z(n24075) );
  NANDN U1571 ( .A(n24097), .B(n24096), .Z(n1163) );
  NANDN U1572 ( .A(n24098), .B(n24099), .Z(n1164) );
  NAND U1573 ( .A(n1163), .B(n1164), .Z(n24102) );
  XOR U1574 ( .A(sreg[1027]), .B(n1903), .Z(n1165) );
  NANDN U1575 ( .A(n1904), .B(n1165), .Z(n1166) );
  NAND U1576 ( .A(sreg[1027]), .B(n1903), .Z(n1167) );
  AND U1577 ( .A(n1166), .B(n1167), .Z(n1943) );
  NAND U1578 ( .A(n1992), .B(n1991), .Z(n1168) );
  XOR U1579 ( .A(n1991), .B(n1992), .Z(n1169) );
  NAND U1580 ( .A(n1169), .B(sreg[1031]), .Z(n1170) );
  NAND U1581 ( .A(n1168), .B(n1170), .Z(n2030) );
  XOR U1582 ( .A(sreg[1036]), .B(n2102), .Z(n1171) );
  NANDN U1583 ( .A(n2103), .B(n1171), .Z(n1172) );
  NAND U1584 ( .A(sreg[1036]), .B(n2102), .Z(n1173) );
  AND U1585 ( .A(n1172), .B(n1173), .Z(n2142) );
  XOR U1586 ( .A(sreg[1040]), .B(n2190), .Z(n1174) );
  NANDN U1587 ( .A(n2191), .B(n1174), .Z(n1175) );
  NAND U1588 ( .A(sreg[1040]), .B(n2190), .Z(n1176) );
  AND U1589 ( .A(n1175), .B(n1176), .Z(n2229) );
  XOR U1590 ( .A(sreg[1045]), .B(n2301), .Z(n1177) );
  NANDN U1591 ( .A(n2302), .B(n1177), .Z(n1178) );
  NAND U1592 ( .A(sreg[1045]), .B(n2301), .Z(n1179) );
  AND U1593 ( .A(n1178), .B(n1179), .Z(n2341) );
  XOR U1594 ( .A(sreg[1049]), .B(n2387), .Z(n1180) );
  NANDN U1595 ( .A(n2388), .B(n1180), .Z(n1181) );
  NAND U1596 ( .A(sreg[1049]), .B(n2387), .Z(n1182) );
  AND U1597 ( .A(n1181), .B(n1182), .Z(n2426) );
  XOR U1598 ( .A(n2513), .B(sreg[1054]), .Z(n1183) );
  NAND U1599 ( .A(n1183), .B(n2512), .Z(n1184) );
  NAND U1600 ( .A(n2513), .B(sreg[1054]), .Z(n1185) );
  AND U1601 ( .A(n1184), .B(n1185), .Z(n2535) );
  NAND U1602 ( .A(n2577), .B(sreg[1058]), .Z(n1186) );
  XOR U1603 ( .A(sreg[1058]), .B(n2577), .Z(n1187) );
  NANDN U1604 ( .A(n2576), .B(n1187), .Z(n1188) );
  NAND U1605 ( .A(n1186), .B(n1188), .Z(n2597) );
  NAND U1606 ( .A(sreg[1062]), .B(n2682), .Z(n1189) );
  XOR U1607 ( .A(n2682), .B(sreg[1062]), .Z(n1190) );
  NANDN U1608 ( .A(n2683), .B(n1190), .Z(n1191) );
  NAND U1609 ( .A(n1189), .B(n1191), .Z(n2685) );
  NAND U1610 ( .A(n2753), .B(sreg[1066]), .Z(n1192) );
  XOR U1611 ( .A(sreg[1066]), .B(n2753), .Z(n1193) );
  NANDN U1612 ( .A(n2752), .B(n1193), .Z(n1194) );
  NAND U1613 ( .A(n1192), .B(n1194), .Z(n2791) );
  NAND U1614 ( .A(n2887), .B(n2886), .Z(n1195) );
  XOR U1615 ( .A(n2886), .B(n2887), .Z(n1196) );
  NANDN U1616 ( .A(sreg[1072]), .B(n1196), .Z(n1197) );
  NAND U1617 ( .A(n1195), .B(n1197), .Z(n2926) );
  NAND U1618 ( .A(sreg[1078]), .B(n3038), .Z(n1198) );
  XOR U1619 ( .A(n3038), .B(sreg[1078]), .Z(n1199) );
  NANDN U1620 ( .A(n3039), .B(n1199), .Z(n1200) );
  NAND U1621 ( .A(n1198), .B(n1200), .Z(n3041) );
  XOR U1622 ( .A(sreg[1082]), .B(n3106), .Z(n1201) );
  NANDN U1623 ( .A(n3107), .B(n1201), .Z(n1202) );
  NAND U1624 ( .A(sreg[1082]), .B(n3106), .Z(n1203) );
  AND U1625 ( .A(n1202), .B(n1203), .Z(n3146) );
  NAND U1626 ( .A(n3192), .B(sreg[1086]), .Z(n1204) );
  XOR U1627 ( .A(sreg[1086]), .B(n3192), .Z(n1205) );
  NANDN U1628 ( .A(n3193), .B(n1205), .Z(n1206) );
  NAND U1629 ( .A(n1204), .B(n1206), .Z(n3232) );
  NAND U1630 ( .A(sreg[1092]), .B(n3338), .Z(n1207) );
  XOR U1631 ( .A(n3338), .B(sreg[1092]), .Z(n1208) );
  NANDN U1632 ( .A(n3339), .B(n1208), .Z(n1209) );
  NAND U1633 ( .A(n1207), .B(n1209), .Z(n3341) );
  NAND U1634 ( .A(n3407), .B(n3406), .Z(n1210) );
  XOR U1635 ( .A(n3406), .B(n3407), .Z(n1211) );
  NANDN U1636 ( .A(sreg[1096]), .B(n1211), .Z(n1212) );
  NAND U1637 ( .A(n1210), .B(n1212), .Z(n3428) );
  NAND U1638 ( .A(sreg[1100]), .B(n3510), .Z(n1213) );
  XOR U1639 ( .A(n3510), .B(sreg[1100]), .Z(n1214) );
  NANDN U1640 ( .A(n3511), .B(n1214), .Z(n1215) );
  NAND U1641 ( .A(n1213), .B(n1215), .Z(n3531) );
  NAND U1642 ( .A(n3579), .B(sreg[1104]), .Z(n1216) );
  XOR U1643 ( .A(sreg[1104]), .B(n3579), .Z(n1217) );
  NANDN U1644 ( .A(n3578), .B(n1217), .Z(n1218) );
  NAND U1645 ( .A(n1216), .B(n1218), .Z(n3617) );
  NAND U1646 ( .A(n3685), .B(sreg[1109]), .Z(n1219) );
  XOR U1647 ( .A(sreg[1109]), .B(n3685), .Z(n1220) );
  NANDN U1648 ( .A(n3686), .B(n1220), .Z(n1221) );
  NAND U1649 ( .A(n1219), .B(n1221), .Z(n3724) );
  XOR U1650 ( .A(n3797), .B(n3796), .Z(n1222) );
  NANDN U1651 ( .A(sreg[1114]), .B(n1222), .Z(n1223) );
  NAND U1652 ( .A(n3797), .B(n3796), .Z(n1224) );
  AND U1653 ( .A(n1223), .B(n1224), .Z(n3835) );
  XOR U1654 ( .A(sreg[1120]), .B(n3927), .Z(n1225) );
  NANDN U1655 ( .A(n3928), .B(n1225), .Z(n1226) );
  NAND U1656 ( .A(sreg[1120]), .B(n3927), .Z(n1227) );
  AND U1657 ( .A(n1226), .B(n1227), .Z(n3962) );
  XOR U1658 ( .A(sreg[1125]), .B(n4033), .Z(n1228) );
  NANDN U1659 ( .A(n4034), .B(n1228), .Z(n1229) );
  NAND U1660 ( .A(sreg[1125]), .B(n4033), .Z(n1230) );
  AND U1661 ( .A(n1229), .B(n1230), .Z(n4073) );
  NAND U1662 ( .A(n4143), .B(n4142), .Z(n1231) );
  XOR U1663 ( .A(n4142), .B(n4143), .Z(n1232) );
  NANDN U1664 ( .A(sreg[1130]), .B(n1232), .Z(n1233) );
  NAND U1665 ( .A(n1231), .B(n1233), .Z(n4182) );
  NAND U1666 ( .A(n4341), .B(sreg[1138]), .Z(n1234) );
  XOR U1667 ( .A(sreg[1138]), .B(n4341), .Z(n1235) );
  NAND U1668 ( .A(n1235), .B(n4340), .Z(n1236) );
  NAND U1669 ( .A(n1234), .B(n1236), .Z(n4361) );
  NAND U1670 ( .A(n4425), .B(n4424), .Z(n1237) );
  XOR U1671 ( .A(n4424), .B(n4425), .Z(n1238) );
  NAND U1672 ( .A(n1238), .B(sreg[1142]), .Z(n1239) );
  NAND U1673 ( .A(n1237), .B(n1239), .Z(n4427) );
  XOR U1674 ( .A(sreg[1146]), .B(n4492), .Z(n1240) );
  NANDN U1675 ( .A(n4493), .B(n1240), .Z(n1241) );
  NAND U1676 ( .A(sreg[1146]), .B(n4492), .Z(n1242) );
  AND U1677 ( .A(n1241), .B(n1242), .Z(n4532) );
  XOR U1678 ( .A(sreg[1150]), .B(n4582), .Z(n1243) );
  NANDN U1679 ( .A(n4583), .B(n1243), .Z(n1244) );
  NAND U1680 ( .A(sreg[1150]), .B(n4582), .Z(n1245) );
  AND U1681 ( .A(n1244), .B(n1245), .Z(n4622) );
  NAND U1682 ( .A(n4740), .B(n4739), .Z(n1246) );
  XOR U1683 ( .A(n4739), .B(n4740), .Z(n1247) );
  NAND U1684 ( .A(n1247), .B(sreg[1157]), .Z(n1248) );
  NAND U1685 ( .A(n1246), .B(n1248), .Z(n4760) );
  XOR U1686 ( .A(n4851), .B(n4850), .Z(n1249) );
  NANDN U1687 ( .A(sreg[1162]), .B(n1249), .Z(n1250) );
  NAND U1688 ( .A(n4851), .B(n4850), .Z(n1251) );
  AND U1689 ( .A(n1250), .B(n1251), .Z(n4889) );
  NAND U1690 ( .A(n4962), .B(n4961), .Z(n1252) );
  XOR U1691 ( .A(n4961), .B(n4962), .Z(n1253) );
  NAND U1692 ( .A(n1253), .B(sreg[1167]), .Z(n1254) );
  NAND U1693 ( .A(n1252), .B(n1254), .Z(n5000) );
  NAND U1694 ( .A(n5091), .B(sreg[1172]), .Z(n1255) );
  XOR U1695 ( .A(sreg[1172]), .B(n5091), .Z(n1256) );
  NANDN U1696 ( .A(n5090), .B(n1256), .Z(n1257) );
  NAND U1697 ( .A(n1255), .B(n1257), .Z(n5093) );
  NAND U1698 ( .A(sreg[1176]), .B(n5178), .Z(n1258) );
  XOR U1699 ( .A(n5178), .B(sreg[1176]), .Z(n1259) );
  NANDN U1700 ( .A(n5179), .B(n1259), .Z(n1260) );
  NAND U1701 ( .A(n1258), .B(n1260), .Z(n5181) );
  XOR U1702 ( .A(sreg[1180]), .B(n5248), .Z(n1261) );
  NANDN U1703 ( .A(n5249), .B(n1261), .Z(n1262) );
  NAND U1704 ( .A(sreg[1180]), .B(n5248), .Z(n1263) );
  AND U1705 ( .A(n1262), .B(n1263), .Z(n5288) );
  NAND U1706 ( .A(n5378), .B(n5377), .Z(n1264) );
  XOR U1707 ( .A(n5377), .B(n5378), .Z(n1265) );
  NAND U1708 ( .A(n1265), .B(sreg[1185]), .Z(n1266) );
  NAND U1709 ( .A(n1264), .B(n1266), .Z(n5380) );
  NAND U1710 ( .A(n5448), .B(sreg[1189]), .Z(n1267) );
  XOR U1711 ( .A(sreg[1189]), .B(n5448), .Z(n1268) );
  NANDN U1712 ( .A(n5447), .B(n1268), .Z(n1269) );
  NAND U1713 ( .A(n1267), .B(n1269), .Z(n5486) );
  XOR U1714 ( .A(n5621), .B(n5620), .Z(n1270) );
  NANDN U1715 ( .A(sreg[1196]), .B(n1270), .Z(n1271) );
  NAND U1716 ( .A(n5621), .B(n5620), .Z(n1272) );
  AND U1717 ( .A(n1271), .B(n1272), .Z(n5642) );
  XOR U1718 ( .A(sreg[1200]), .B(n5686), .Z(n1273) );
  NANDN U1719 ( .A(n5687), .B(n1273), .Z(n1274) );
  NAND U1720 ( .A(sreg[1200]), .B(n5686), .Z(n1275) );
  AND U1721 ( .A(n1274), .B(n1275), .Z(n5722) );
  NAND U1722 ( .A(n5771), .B(n5770), .Z(n1276) );
  XOR U1723 ( .A(n5770), .B(n5771), .Z(n1277) );
  NAND U1724 ( .A(n1277), .B(sreg[1204]), .Z(n1278) );
  NAND U1725 ( .A(n1276), .B(n1278), .Z(n5809) );
  XOR U1726 ( .A(sreg[1211]), .B(n5927), .Z(n1279) );
  NANDN U1727 ( .A(n5928), .B(n1279), .Z(n1280) );
  NAND U1728 ( .A(sreg[1211]), .B(n5927), .Z(n1281) );
  AND U1729 ( .A(n1280), .B(n1281), .Z(n5967) );
  NAND U1730 ( .A(n6035), .B(n6034), .Z(n1282) );
  XOR U1731 ( .A(n6034), .B(n6035), .Z(n1283) );
  NAND U1732 ( .A(n1283), .B(sreg[1216]), .Z(n1284) );
  NAND U1733 ( .A(n1282), .B(n1284), .Z(n6073) );
  XOR U1734 ( .A(n6123), .B(n6122), .Z(n1285) );
  NANDN U1735 ( .A(sreg[1220]), .B(n1285), .Z(n1286) );
  NAND U1736 ( .A(n6123), .B(n6122), .Z(n1287) );
  AND U1737 ( .A(n1286), .B(n1287), .Z(n6161) );
  XOR U1738 ( .A(n6229), .B(sreg[1224]), .Z(n1288) );
  NANDN U1739 ( .A(n6228), .B(n1288), .Z(n1289) );
  NAND U1740 ( .A(n6229), .B(sreg[1224]), .Z(n1290) );
  AND U1741 ( .A(n1289), .B(n1290), .Z(n6231) );
  XOR U1742 ( .A(sreg[1228]), .B(n6300), .Z(n1291) );
  NANDN U1743 ( .A(n6301), .B(n1291), .Z(n1292) );
  NAND U1744 ( .A(sreg[1228]), .B(n6300), .Z(n1293) );
  AND U1745 ( .A(n1292), .B(n1293), .Z(n6340) );
  XOR U1746 ( .A(n6430), .B(n6429), .Z(n1294) );
  NAND U1747 ( .A(n1294), .B(sreg[1233]), .Z(n1295) );
  NAND U1748 ( .A(n6430), .B(n6429), .Z(n1296) );
  AND U1749 ( .A(n1295), .B(n1296), .Z(n6432) );
  NAND U1750 ( .A(n6500), .B(sreg[1237]), .Z(n1297) );
  XOR U1751 ( .A(sreg[1237]), .B(n6500), .Z(n1298) );
  NANDN U1752 ( .A(n6499), .B(n1298), .Z(n1299) );
  NAND U1753 ( .A(n1297), .B(n1299), .Z(n6538) );
  NAND U1754 ( .A(n6632), .B(sreg[1243]), .Z(n1300) );
  XOR U1755 ( .A(sreg[1243]), .B(n6632), .Z(n1301) );
  NANDN U1756 ( .A(n6633), .B(n1301), .Z(n1302) );
  NAND U1757 ( .A(n1300), .B(n1302), .Z(n6666) );
  NAND U1758 ( .A(sreg[1248]), .B(n6754), .Z(n1303) );
  XOR U1759 ( .A(n6754), .B(sreg[1248]), .Z(n1304) );
  NANDN U1760 ( .A(n6755), .B(n1304), .Z(n1305) );
  NAND U1761 ( .A(n1303), .B(n1305), .Z(n6775) );
  XOR U1762 ( .A(sreg[1252]), .B(n6822), .Z(n1306) );
  NANDN U1763 ( .A(n6823), .B(n1306), .Z(n1307) );
  NAND U1764 ( .A(sreg[1252]), .B(n6822), .Z(n1308) );
  AND U1765 ( .A(n1307), .B(n1308), .Z(n6862) );
  NAND U1766 ( .A(n6980), .B(n6979), .Z(n1309) );
  XOR U1767 ( .A(n6979), .B(n6980), .Z(n1310) );
  NAND U1768 ( .A(n1310), .B(sreg[1259]), .Z(n1311) );
  NAND U1769 ( .A(n1309), .B(n1311), .Z(n7019) );
  XOR U1770 ( .A(n7123), .B(sreg[1265]), .Z(n1312) );
  NANDN U1771 ( .A(n7124), .B(n1312), .Z(n1313) );
  NAND U1772 ( .A(n7123), .B(sreg[1265]), .Z(n1314) );
  AND U1773 ( .A(n1313), .B(n1314), .Z(n7144) );
  NAND U1774 ( .A(n7190), .B(n7189), .Z(n1315) );
  XOR U1775 ( .A(n7189), .B(n7190), .Z(n1316) );
  NAND U1776 ( .A(n1316), .B(sreg[1269]), .Z(n1317) );
  NAND U1777 ( .A(n1315), .B(n1317), .Z(n7228) );
  XOR U1778 ( .A(sreg[1273]), .B(n7277), .Z(n1318) );
  NANDN U1779 ( .A(n7278), .B(n1318), .Z(n1319) );
  NAND U1780 ( .A(sreg[1273]), .B(n7277), .Z(n1320) );
  AND U1781 ( .A(n1319), .B(n1320), .Z(n7317) );
  NAND U1782 ( .A(n7412), .B(n7411), .Z(n1321) );
  XOR U1783 ( .A(n7411), .B(n7412), .Z(n1322) );
  NAND U1784 ( .A(n1322), .B(sreg[1279]), .Z(n1323) );
  NAND U1785 ( .A(n1321), .B(n1323), .Z(n7451) );
  NAND U1786 ( .A(sreg[1283]), .B(n7515), .Z(n1324) );
  XOR U1787 ( .A(n7515), .B(sreg[1283]), .Z(n1325) );
  NANDN U1788 ( .A(n7516), .B(n1325), .Z(n1326) );
  NAND U1789 ( .A(n1324), .B(n1326), .Z(n7536) );
  XOR U1790 ( .A(n7602), .B(sreg[1287]), .Z(n1327) );
  NANDN U1791 ( .A(n7601), .B(n1327), .Z(n1328) );
  NAND U1792 ( .A(n7602), .B(sreg[1287]), .Z(n1329) );
  AND U1793 ( .A(n1328), .B(n1329), .Z(n7604) );
  XOR U1794 ( .A(n7688), .B(n7687), .Z(n1330) );
  NANDN U1795 ( .A(sreg[1291]), .B(n1330), .Z(n1331) );
  NAND U1796 ( .A(n7688), .B(n7687), .Z(n1332) );
  AND U1797 ( .A(n1331), .B(n1332), .Z(n7690) );
  NAND U1798 ( .A(n7758), .B(sreg[1295]), .Z(n1333) );
  XOR U1799 ( .A(sreg[1295]), .B(n7758), .Z(n1334) );
  NANDN U1800 ( .A(n7757), .B(n1334), .Z(n1335) );
  NAND U1801 ( .A(n1333), .B(n1335), .Z(n7792) );
  NAND U1802 ( .A(n7863), .B(sreg[1300]), .Z(n1336) );
  XOR U1803 ( .A(sreg[1300]), .B(n7863), .Z(n1337) );
  NANDN U1804 ( .A(n7862), .B(n1337), .Z(n1338) );
  NAND U1805 ( .A(n1336), .B(n1338), .Z(n7901) );
  NAND U1806 ( .A(n7972), .B(n7971), .Z(n1339) );
  XOR U1807 ( .A(n7971), .B(n7972), .Z(n1340) );
  NAND U1808 ( .A(n1340), .B(sreg[1305]), .Z(n1341) );
  NAND U1809 ( .A(n1339), .B(n1341), .Z(n8010) );
  XOR U1810 ( .A(n8080), .B(sreg[1310]), .Z(n1342) );
  NANDN U1811 ( .A(n8079), .B(n1342), .Z(n1343) );
  NAND U1812 ( .A(n8080), .B(sreg[1310]), .Z(n1344) );
  AND U1813 ( .A(n1343), .B(n1344), .Z(n8098) );
  NAND U1814 ( .A(n8179), .B(sreg[1314]), .Z(n1345) );
  XOR U1815 ( .A(sreg[1314]), .B(n8179), .Z(n1346) );
  NAND U1816 ( .A(n1346), .B(n8178), .Z(n1347) );
  NAND U1817 ( .A(n1345), .B(n1347), .Z(n8199) );
  NAND U1818 ( .A(n8245), .B(n8244), .Z(n1348) );
  XOR U1819 ( .A(n8244), .B(n8245), .Z(n1349) );
  NAND U1820 ( .A(n1349), .B(sreg[1318]), .Z(n1350) );
  NAND U1821 ( .A(n1348), .B(n1350), .Z(n8283) );
  XOR U1822 ( .A(n8354), .B(sreg[1323]), .Z(n1351) );
  NAND U1823 ( .A(n1351), .B(n8353), .Z(n1352) );
  NAND U1824 ( .A(n8354), .B(sreg[1323]), .Z(n1353) );
  AND U1825 ( .A(n1352), .B(n1353), .Z(n8374) );
  NAND U1826 ( .A(n8437), .B(sreg[1327]), .Z(n1354) );
  XOR U1827 ( .A(sreg[1327]), .B(n8437), .Z(n1355) );
  NANDN U1828 ( .A(n8438), .B(n1355), .Z(n1356) );
  NAND U1829 ( .A(n1354), .B(n1356), .Z(n8477) );
  NAND U1830 ( .A(n8582), .B(sreg[1333]), .Z(n1357) );
  XOR U1831 ( .A(sreg[1333]), .B(n8582), .Z(n1358) );
  NAND U1832 ( .A(n1358), .B(n8581), .Z(n1359) );
  NAND U1833 ( .A(n1357), .B(n1359), .Z(n8602) );
  NAND U1834 ( .A(n8648), .B(n8647), .Z(n1360) );
  XOR U1835 ( .A(n8647), .B(n8648), .Z(n1361) );
  NAND U1836 ( .A(n1361), .B(sreg[1337]), .Z(n1362) );
  NAND U1837 ( .A(n1360), .B(n1362), .Z(n8686) );
  XOR U1838 ( .A(sreg[1342]), .B(n8758), .Z(n1363) );
  NANDN U1839 ( .A(n8759), .B(n1363), .Z(n1364) );
  NAND U1840 ( .A(sreg[1342]), .B(n8758), .Z(n1365) );
  AND U1841 ( .A(n1364), .B(n1365), .Z(n8798) );
  XOR U1842 ( .A(n8891), .B(n8890), .Z(n1366) );
  NANDN U1843 ( .A(sreg[1348]), .B(n1366), .Z(n1367) );
  NAND U1844 ( .A(n8891), .B(n8890), .Z(n1368) );
  AND U1845 ( .A(n1367), .B(n1368), .Z(n8929) );
  XOR U1846 ( .A(sreg[1355]), .B(n9047), .Z(n1369) );
  NANDN U1847 ( .A(n9048), .B(n1369), .Z(n1370) );
  NAND U1848 ( .A(sreg[1355]), .B(n9047), .Z(n1371) );
  AND U1849 ( .A(n1370), .B(n1371), .Z(n9087) );
  XOR U1850 ( .A(sreg[1360]), .B(n9156), .Z(n1372) );
  NANDN U1851 ( .A(n9157), .B(n1372), .Z(n1373) );
  NAND U1852 ( .A(sreg[1360]), .B(n9156), .Z(n1374) );
  AND U1853 ( .A(n1373), .B(n1374), .Z(n9196) );
  NAND U1854 ( .A(n9243), .B(n9242), .Z(n1375) );
  XOR U1855 ( .A(n9242), .B(n9243), .Z(n1376) );
  NANDN U1856 ( .A(sreg[1364]), .B(n1376), .Z(n1377) );
  NAND U1857 ( .A(n1375), .B(n1377), .Z(n9282) );
  XOR U1858 ( .A(sreg[1370]), .B(n9374), .Z(n1378) );
  NANDN U1859 ( .A(n9375), .B(n1378), .Z(n1379) );
  NAND U1860 ( .A(sreg[1370]), .B(n9374), .Z(n1380) );
  AND U1861 ( .A(n1379), .B(n1380), .Z(n9414) );
  NAND U1862 ( .A(n9503), .B(sreg[1375]), .Z(n1381) );
  XOR U1863 ( .A(sreg[1375]), .B(n9503), .Z(n1382) );
  NAND U1864 ( .A(n1382), .B(n9502), .Z(n1383) );
  NAND U1865 ( .A(n1381), .B(n1383), .Z(n9505) );
  XOR U1866 ( .A(n9584), .B(n9583), .Z(n1384) );
  NAND U1867 ( .A(n1384), .B(sreg[1379]), .Z(n1385) );
  NAND U1868 ( .A(n9584), .B(n9583), .Z(n1386) );
  AND U1869 ( .A(n1385), .B(n1386), .Z(n9604) );
  NAND U1870 ( .A(n9650), .B(n9649), .Z(n1387) );
  XOR U1871 ( .A(n9649), .B(n9650), .Z(n1388) );
  NANDN U1872 ( .A(sreg[1383]), .B(n1388), .Z(n1389) );
  NAND U1873 ( .A(n1387), .B(n1389), .Z(n9689) );
  NAND U1874 ( .A(sreg[1388]), .B(n9779), .Z(n1390) );
  XOR U1875 ( .A(n9779), .B(sreg[1388]), .Z(n1391) );
  NANDN U1876 ( .A(n9778), .B(n1391), .Z(n1392) );
  NAND U1877 ( .A(n1390), .B(n1392), .Z(n9781) );
  XOR U1878 ( .A(sreg[1392]), .B(n9848), .Z(n1393) );
  NANDN U1879 ( .A(n9849), .B(n1393), .Z(n1394) );
  NAND U1880 ( .A(sreg[1392]), .B(n9848), .Z(n1395) );
  AND U1881 ( .A(n1394), .B(n1395), .Z(n9886) );
  XOR U1882 ( .A(n9954), .B(n9953), .Z(n1396) );
  NANDN U1883 ( .A(sreg[1397]), .B(n1396), .Z(n1397) );
  NAND U1884 ( .A(n9954), .B(n9953), .Z(n1398) );
  AND U1885 ( .A(n1397), .B(n1398), .Z(n9993) );
  XOR U1886 ( .A(sreg[1403]), .B(n10079), .Z(n1399) );
  NANDN U1887 ( .A(n10080), .B(n1399), .Z(n1400) );
  NAND U1888 ( .A(sreg[1403]), .B(n10079), .Z(n1401) );
  AND U1889 ( .A(n1400), .B(n1401), .Z(n10120) );
  NAND U1890 ( .A(n10231), .B(n10230), .Z(n1402) );
  XOR U1891 ( .A(n10230), .B(n10231), .Z(n1403) );
  NAND U1892 ( .A(n1403), .B(sreg[1410]), .Z(n1404) );
  NAND U1893 ( .A(n1402), .B(n1404), .Z(n10269) );
  NAND U1894 ( .A(n10365), .B(n10364), .Z(n1405) );
  XOR U1895 ( .A(n10364), .B(n10365), .Z(n1406) );
  NAND U1896 ( .A(n1406), .B(sreg[1416]), .Z(n1407) );
  NAND U1897 ( .A(n1405), .B(n1407), .Z(n10403) );
  XOR U1898 ( .A(sreg[1420]), .B(n10454), .Z(n1408) );
  NANDN U1899 ( .A(n10455), .B(n1408), .Z(n1409) );
  NAND U1900 ( .A(sreg[1420]), .B(n10454), .Z(n1410) );
  AND U1901 ( .A(n1409), .B(n1410), .Z(n10494) );
  XOR U1902 ( .A(sreg[1424]), .B(n10542), .Z(n1411) );
  NANDN U1903 ( .A(n10543), .B(n1411), .Z(n1412) );
  NAND U1904 ( .A(sreg[1424]), .B(n10542), .Z(n1413) );
  AND U1905 ( .A(n1412), .B(n1413), .Z(n10582) );
  NAND U1906 ( .A(n10652), .B(sreg[1429]), .Z(n1414) );
  XOR U1907 ( .A(sreg[1429]), .B(n10652), .Z(n1415) );
  NANDN U1908 ( .A(n10651), .B(n1415), .Z(n1416) );
  NAND U1909 ( .A(n1414), .B(n1416), .Z(n10690) );
  XOR U1910 ( .A(n10763), .B(n10762), .Z(n1417) );
  NANDN U1911 ( .A(sreg[1434]), .B(n1417), .Z(n1418) );
  NAND U1912 ( .A(n10763), .B(n10762), .Z(n1419) );
  AND U1913 ( .A(n1418), .B(n1419), .Z(n10801) );
  XOR U1914 ( .A(sreg[1439]), .B(n10873), .Z(n1420) );
  NANDN U1915 ( .A(n10874), .B(n1420), .Z(n1421) );
  NAND U1916 ( .A(sreg[1439]), .B(n10873), .Z(n1422) );
  AND U1917 ( .A(n1421), .B(n1422), .Z(n10913) );
  XOR U1918 ( .A(n11008), .B(sreg[1445]), .Z(n1423) );
  NAND U1919 ( .A(n1423), .B(n11007), .Z(n1424) );
  NAND U1920 ( .A(n11008), .B(sreg[1445]), .Z(n1425) );
  AND U1921 ( .A(n1424), .B(n1425), .Z(n11047) );
  XOR U1922 ( .A(sreg[1450]), .B(n11118), .Z(n1426) );
  NANDN U1923 ( .A(n11119), .B(n1426), .Z(n1427) );
  NAND U1924 ( .A(sreg[1450]), .B(n11118), .Z(n1428) );
  AND U1925 ( .A(n1427), .B(n1428), .Z(n11158) );
  XOR U1926 ( .A(sreg[1455]), .B(n11229), .Z(n1429) );
  NANDN U1927 ( .A(n11230), .B(n1429), .Z(n1430) );
  NAND U1928 ( .A(sreg[1455]), .B(n11229), .Z(n1431) );
  AND U1929 ( .A(n1430), .B(n1431), .Z(n11269) );
  XOR U1930 ( .A(sreg[1461]), .B(n11361), .Z(n1432) );
  NANDN U1931 ( .A(n11362), .B(n1432), .Z(n1433) );
  NAND U1932 ( .A(sreg[1461]), .B(n11361), .Z(n1434) );
  AND U1933 ( .A(n1433), .B(n1434), .Z(n11383) );
  XOR U1934 ( .A(sreg[1466]), .B(n11471), .Z(n1435) );
  NANDN U1935 ( .A(n11472), .B(n1435), .Z(n1436) );
  NAND U1936 ( .A(sreg[1466]), .B(n11471), .Z(n1437) );
  AND U1937 ( .A(n1436), .B(n1437), .Z(n11506) );
  XOR U1938 ( .A(sreg[1472]), .B(n11595), .Z(n1438) );
  NANDN U1939 ( .A(n11596), .B(n1438), .Z(n1439) );
  NAND U1940 ( .A(sreg[1472]), .B(n11595), .Z(n1440) );
  AND U1941 ( .A(n1439), .B(n1440), .Z(n11630) );
  NAND U1942 ( .A(n11702), .B(sreg[1477]), .Z(n1441) );
  XOR U1943 ( .A(sreg[1477]), .B(n11702), .Z(n1442) );
  NANDN U1944 ( .A(n11701), .B(n1442), .Z(n1443) );
  NAND U1945 ( .A(n1441), .B(n1443), .Z(n11723) );
  NAND U1946 ( .A(sreg[1488]), .B(n11966), .Z(n1444) );
  XOR U1947 ( .A(n11966), .B(sreg[1488]), .Z(n1445) );
  NANDN U1948 ( .A(n11967), .B(n1445), .Z(n1446) );
  NAND U1949 ( .A(n1444), .B(n1446), .Z(n11987) );
  XOR U1950 ( .A(sreg[1492]), .B(n12032), .Z(n1447) );
  NANDN U1951 ( .A(n12033), .B(n1447), .Z(n1448) );
  NAND U1952 ( .A(sreg[1492]), .B(n12032), .Z(n1449) );
  AND U1953 ( .A(n1448), .B(n1449), .Z(n12072) );
  NAND U1954 ( .A(n12142), .B(n12141), .Z(n1450) );
  XOR U1955 ( .A(n12141), .B(n12142), .Z(n1451) );
  NAND U1956 ( .A(n1451), .B(sreg[1497]), .Z(n1452) );
  NAND U1957 ( .A(n1450), .B(n1452), .Z(n12163) );
  XOR U1958 ( .A(n12246), .B(n12245), .Z(n1453) );
  NAND U1959 ( .A(n1453), .B(sreg[1501]), .Z(n1454) );
  NAND U1960 ( .A(n12246), .B(n12245), .Z(n1455) );
  AND U1961 ( .A(n1454), .B(n1455), .Z(n12248) );
  XOR U1962 ( .A(sreg[1505]), .B(n12309), .Z(n1456) );
  NANDN U1963 ( .A(n12310), .B(n1456), .Z(n1457) );
  NAND U1964 ( .A(sreg[1505]), .B(n12309), .Z(n1458) );
  AND U1965 ( .A(n1457), .B(n1458), .Z(n12349) );
  NAND U1966 ( .A(sreg[1511]), .B(n12461), .Z(n1459) );
  XOR U1967 ( .A(n12461), .B(sreg[1511]), .Z(n1460) );
  NANDN U1968 ( .A(n12462), .B(n1460), .Z(n1461) );
  NAND U1969 ( .A(n1459), .B(n1461), .Z(n12464) );
  NAND U1970 ( .A(n12532), .B(sreg[1515]), .Z(n1462) );
  XOR U1971 ( .A(sreg[1515]), .B(n12532), .Z(n1463) );
  NANDN U1972 ( .A(n12531), .B(n1463), .Z(n1464) );
  NAND U1973 ( .A(n1462), .B(n1464), .Z(n12570) );
  NAND U1974 ( .A(n12645), .B(sreg[1520]), .Z(n1465) );
  XOR U1975 ( .A(sreg[1520]), .B(n12645), .Z(n1466) );
  NANDN U1976 ( .A(n12644), .B(n1466), .Z(n1467) );
  NAND U1977 ( .A(n1465), .B(n1467), .Z(n12683) );
  XOR U1978 ( .A(sreg[1524]), .B(n12732), .Z(n1468) );
  NANDN U1979 ( .A(n12733), .B(n1468), .Z(n1469) );
  NAND U1980 ( .A(sreg[1524]), .B(n12732), .Z(n1470) );
  AND U1981 ( .A(n1469), .B(n1470), .Z(n12772) );
  NAND U1982 ( .A(n12823), .B(sreg[1528]), .Z(n1471) );
  XOR U1983 ( .A(sreg[1528]), .B(n12823), .Z(n1472) );
  NANDN U1984 ( .A(n12822), .B(n1472), .Z(n1473) );
  NAND U1985 ( .A(n1471), .B(n1473), .Z(n12843) );
  XOR U1986 ( .A(n12911), .B(sreg[1532]), .Z(n1474) );
  NAND U1987 ( .A(n1474), .B(n12910), .Z(n1475) );
  NAND U1988 ( .A(n12911), .B(sreg[1532]), .Z(n1476) );
  AND U1989 ( .A(n1475), .B(n1476), .Z(n12950) );
  XOR U1990 ( .A(n13041), .B(sreg[1538]), .Z(n1477) );
  NAND U1991 ( .A(n1477), .B(n13040), .Z(n1478) );
  NAND U1992 ( .A(n13041), .B(sreg[1538]), .Z(n1479) );
  AND U1993 ( .A(n1478), .B(n1479), .Z(n13080) );
  XOR U1994 ( .A(n13129), .B(sreg[1542]), .Z(n1480) );
  NANDN U1995 ( .A(n13128), .B(n1480), .Z(n1481) );
  NAND U1996 ( .A(n13129), .B(sreg[1542]), .Z(n1482) );
  AND U1997 ( .A(n1481), .B(n1482), .Z(n13168) );
  XOR U1998 ( .A(sreg[1547]), .B(n13239), .Z(n1483) );
  NANDN U1999 ( .A(n13240), .B(n1483), .Z(n1484) );
  NAND U2000 ( .A(sreg[1547]), .B(n13239), .Z(n1485) );
  AND U2001 ( .A(n1484), .B(n1485), .Z(n13279) );
  NAND U2002 ( .A(n13349), .B(n13348), .Z(n1486) );
  XOR U2003 ( .A(n13348), .B(n13349), .Z(n1487) );
  NAND U2004 ( .A(n1487), .B(sreg[1552]), .Z(n1488) );
  NAND U2005 ( .A(n1486), .B(n1488), .Z(n13387) );
  XOR U2006 ( .A(n13437), .B(n13436), .Z(n1489) );
  NANDN U2007 ( .A(sreg[1556]), .B(n1489), .Z(n1490) );
  NAND U2008 ( .A(n13437), .B(n13436), .Z(n1491) );
  AND U2009 ( .A(n1490), .B(n1491), .Z(n13475) );
  XOR U2010 ( .A(sreg[1561]), .B(n13545), .Z(n1492) );
  NANDN U2011 ( .A(n13546), .B(n1492), .Z(n1493) );
  NAND U2012 ( .A(sreg[1561]), .B(n13545), .Z(n1494) );
  AND U2013 ( .A(n1493), .B(n1494), .Z(n13585) );
  NAND U2014 ( .A(n13682), .B(n13681), .Z(n1495) );
  XOR U2015 ( .A(n13681), .B(n13682), .Z(n1496) );
  NAND U2016 ( .A(n1496), .B(sreg[1567]), .Z(n1497) );
  NAND U2017 ( .A(n1495), .B(n1497), .Z(n13720) );
  XOR U2018 ( .A(sreg[1575]), .B(n13859), .Z(n1498) );
  NANDN U2019 ( .A(n13860), .B(n1498), .Z(n1499) );
  NAND U2020 ( .A(sreg[1575]), .B(n13859), .Z(n1500) );
  AND U2021 ( .A(n1499), .B(n1500), .Z(n13899) );
  XOR U2022 ( .A(n14017), .B(sreg[1582]), .Z(n1501) );
  NAND U2023 ( .A(n1501), .B(n14016), .Z(n1502) );
  NAND U2024 ( .A(n14017), .B(sreg[1582]), .Z(n1503) );
  AND U2025 ( .A(n1502), .B(n1503), .Z(n14057) );
  XOR U2026 ( .A(n14101), .B(sreg[1586]), .Z(n1504) );
  NANDN U2027 ( .A(n14100), .B(n1504), .Z(n1505) );
  NAND U2028 ( .A(n14101), .B(sreg[1586]), .Z(n1506) );
  AND U2029 ( .A(n1505), .B(n1506), .Z(n14122) );
  NAND U2030 ( .A(n14210), .B(sreg[1591]), .Z(n1507) );
  XOR U2031 ( .A(sreg[1591]), .B(n14210), .Z(n1508) );
  NANDN U2032 ( .A(n14209), .B(n1508), .Z(n1509) );
  NAND U2033 ( .A(n1507), .B(n1509), .Z(n14248) );
  NAND U2034 ( .A(n14298), .B(sreg[1595]), .Z(n1510) );
  XOR U2035 ( .A(sreg[1595]), .B(n14298), .Z(n1511) );
  NANDN U2036 ( .A(n14297), .B(n1511), .Z(n1512) );
  NAND U2037 ( .A(n1510), .B(n1512), .Z(n14336) );
  NAND U2038 ( .A(sreg[1600]), .B(n14426), .Z(n1513) );
  XOR U2039 ( .A(n14426), .B(sreg[1600]), .Z(n1514) );
  NANDN U2040 ( .A(n14427), .B(n1514), .Z(n1515) );
  NAND U2041 ( .A(n1513), .B(n1515), .Z(n14447) );
  XOR U2042 ( .A(sreg[1604]), .B(n14494), .Z(n1516) );
  NANDN U2043 ( .A(n14495), .B(n1516), .Z(n1517) );
  NAND U2044 ( .A(sreg[1604]), .B(n14494), .Z(n1518) );
  AND U2045 ( .A(n1517), .B(n1518), .Z(n14534) );
  XOR U2046 ( .A(sreg[1610]), .B(n14626), .Z(n1519) );
  NANDN U2047 ( .A(n14627), .B(n1519), .Z(n1520) );
  NAND U2048 ( .A(sreg[1610]), .B(n14626), .Z(n1521) );
  AND U2049 ( .A(n1520), .B(n1521), .Z(n14666) );
  XOR U2050 ( .A(sreg[1616]), .B(n14758), .Z(n1522) );
  NANDN U2051 ( .A(n14759), .B(n1522), .Z(n1523) );
  NAND U2052 ( .A(sreg[1616]), .B(n14758), .Z(n1524) );
  AND U2053 ( .A(n1523), .B(n1524), .Z(n14798) );
  XOR U2054 ( .A(n14865), .B(n14864), .Z(n1525) );
  NAND U2055 ( .A(n1525), .B(sreg[1620]), .Z(n1526) );
  NAND U2056 ( .A(n14865), .B(n14864), .Z(n1527) );
  AND U2057 ( .A(n1526), .B(n1527), .Z(n14885) );
  NAND U2058 ( .A(sreg[1624]), .B(n14950), .Z(n1528) );
  XOR U2059 ( .A(n14950), .B(sreg[1624]), .Z(n1529) );
  NANDN U2060 ( .A(n14951), .B(n1529), .Z(n1530) );
  NAND U2061 ( .A(n1528), .B(n1530), .Z(n14971) );
  XOR U2062 ( .A(sreg[1628]), .B(n15018), .Z(n1531) );
  NANDN U2063 ( .A(n15019), .B(n1531), .Z(n1532) );
  NAND U2064 ( .A(sreg[1628]), .B(n15018), .Z(n1533) );
  AND U2065 ( .A(n1532), .B(n1533), .Z(n15058) );
  NAND U2066 ( .A(n15105), .B(n15104), .Z(n1534) );
  XOR U2067 ( .A(n15104), .B(n15105), .Z(n1535) );
  NAND U2068 ( .A(n1535), .B(sreg[1632]), .Z(n1536) );
  NAND U2069 ( .A(n1534), .B(n1536), .Z(n15143) );
  XOR U2070 ( .A(n15193), .B(n15192), .Z(n1537) );
  NANDN U2071 ( .A(sreg[1636]), .B(n1537), .Z(n1538) );
  NAND U2072 ( .A(n15193), .B(n15192), .Z(n1539) );
  AND U2073 ( .A(n1538), .B(n1539), .Z(n15231) );
  NAND U2074 ( .A(n15412), .B(n15411), .Z(n1540) );
  XOR U2075 ( .A(n15411), .B(n15412), .Z(n1541) );
  NAND U2076 ( .A(n1541), .B(sreg[1645]), .Z(n1542) );
  NAND U2077 ( .A(n1540), .B(n1542), .Z(n15433) );
  NAND U2078 ( .A(sreg[1649]), .B(n15497), .Z(n1543) );
  XOR U2079 ( .A(n15497), .B(sreg[1649]), .Z(n1544) );
  NANDN U2080 ( .A(n15498), .B(n1544), .Z(n1545) );
  NAND U2081 ( .A(n1543), .B(n1545), .Z(n15500) );
  XOR U2082 ( .A(sreg[1653]), .B(n15567), .Z(n1546) );
  NANDN U2083 ( .A(n15568), .B(n1546), .Z(n1547) );
  NAND U2084 ( .A(sreg[1653]), .B(n15567), .Z(n1548) );
  AND U2085 ( .A(n1547), .B(n1548), .Z(n15607) );
  XOR U2086 ( .A(sreg[1658]), .B(n15674), .Z(n1549) );
  NANDN U2087 ( .A(n15675), .B(n1549), .Z(n1550) );
  NAND U2088 ( .A(sreg[1658]), .B(n15674), .Z(n1551) );
  AND U2089 ( .A(n1550), .B(n1551), .Z(n15714) );
  XOR U2090 ( .A(n15786), .B(sreg[1663]), .Z(n1552) );
  NAND U2091 ( .A(n1552), .B(n15785), .Z(n1553) );
  NAND U2092 ( .A(n15786), .B(sreg[1663]), .Z(n1554) );
  AND U2093 ( .A(n1553), .B(n1554), .Z(n15825) );
  XOR U2094 ( .A(n15920), .B(sreg[1669]), .Z(n1555) );
  NAND U2095 ( .A(n1555), .B(n15919), .Z(n1556) );
  NAND U2096 ( .A(n15920), .B(sreg[1669]), .Z(n1557) );
  AND U2097 ( .A(n1556), .B(n1557), .Z(n15941) );
  XOR U2098 ( .A(n16032), .B(n16031), .Z(n1558) );
  NANDN U2099 ( .A(sreg[1674]), .B(n1558), .Z(n1559) );
  NAND U2100 ( .A(n16032), .B(n16031), .Z(n1560) );
  AND U2101 ( .A(n1559), .B(n1560), .Z(n16065) );
  NAND U2102 ( .A(n16110), .B(sreg[1678]), .Z(n1561) );
  XOR U2103 ( .A(sreg[1678]), .B(n16110), .Z(n1562) );
  NANDN U2104 ( .A(n16111), .B(n1562), .Z(n1563) );
  NAND U2105 ( .A(n1561), .B(n1563), .Z(n16151) );
  XOR U2106 ( .A(n16195), .B(sreg[1682]), .Z(n1564) );
  NAND U2107 ( .A(n1564), .B(n16194), .Z(n1565) );
  NAND U2108 ( .A(n16195), .B(sreg[1682]), .Z(n1566) );
  AND U2109 ( .A(n1565), .B(n1566), .Z(n16216) );
  NAND U2110 ( .A(n16302), .B(n16301), .Z(n1567) );
  XOR U2111 ( .A(n16301), .B(n16302), .Z(n1568) );
  NAND U2112 ( .A(n1568), .B(sreg[1687]), .Z(n1569) );
  NAND U2113 ( .A(n1567), .B(n1569), .Z(n16340) );
  XOR U2114 ( .A(sreg[1691]), .B(n16389), .Z(n1570) );
  NANDN U2115 ( .A(n16390), .B(n1570), .Z(n1571) );
  NAND U2116 ( .A(sreg[1691]), .B(n16389), .Z(n1572) );
  AND U2117 ( .A(n1571), .B(n1572), .Z(n16429) );
  NAND U2118 ( .A(sreg[1697]), .B(n16541), .Z(n1573) );
  XOR U2119 ( .A(n16541), .B(sreg[1697]), .Z(n1574) );
  NANDN U2120 ( .A(n16542), .B(n1574), .Z(n1575) );
  NAND U2121 ( .A(n1573), .B(n1575), .Z(n16544) );
  NAND U2122 ( .A(sreg[1701]), .B(n16629), .Z(n1576) );
  XOR U2123 ( .A(n16629), .B(sreg[1701]), .Z(n1577) );
  NANDN U2124 ( .A(n16630), .B(n1577), .Z(n1578) );
  NAND U2125 ( .A(n1576), .B(n1578), .Z(n16650) );
  XOR U2126 ( .A(sreg[1705]), .B(n16697), .Z(n1579) );
  NANDN U2127 ( .A(n16698), .B(n1579), .Z(n1580) );
  NAND U2128 ( .A(sreg[1705]), .B(n16697), .Z(n1581) );
  AND U2129 ( .A(n1580), .B(n1581), .Z(n16737) );
  XOR U2130 ( .A(n16822), .B(sreg[1710]), .Z(n1582) );
  NANDN U2131 ( .A(n16823), .B(n1582), .Z(n1583) );
  NAND U2132 ( .A(n16822), .B(sreg[1710]), .Z(n1584) );
  AND U2133 ( .A(n1583), .B(n1584), .Z(n16825) );
  XOR U2134 ( .A(sreg[1714]), .B(n16886), .Z(n1585) );
  NANDN U2135 ( .A(n16887), .B(n1585), .Z(n1586) );
  NAND U2136 ( .A(sreg[1714]), .B(n16886), .Z(n1587) );
  AND U2137 ( .A(n1586), .B(n1587), .Z(n16926) );
  XOR U2138 ( .A(n17014), .B(n17013), .Z(n1588) );
  NAND U2139 ( .A(n1588), .B(sreg[1719]), .Z(n1589) );
  NAND U2140 ( .A(n17014), .B(n17013), .Z(n1590) );
  AND U2141 ( .A(n1589), .B(n1590), .Z(n17016) );
  XOR U2142 ( .A(sreg[1723]), .B(n17081), .Z(n1591) );
  NANDN U2143 ( .A(n17082), .B(n1591), .Z(n1592) );
  NAND U2144 ( .A(sreg[1723]), .B(n17081), .Z(n1593) );
  AND U2145 ( .A(n1592), .B(n1593), .Z(n17121) );
  XOR U2146 ( .A(n17255), .B(n17254), .Z(n1594) );
  NANDN U2147 ( .A(sreg[1730]), .B(n1594), .Z(n1595) );
  NAND U2148 ( .A(n17255), .B(n17254), .Z(n1596) );
  AND U2149 ( .A(n1595), .B(n1596), .Z(n17275) );
  NAND U2150 ( .A(sreg[1734]), .B(n17340), .Z(n1597) );
  XOR U2151 ( .A(n17340), .B(sreg[1734]), .Z(n1598) );
  NANDN U2152 ( .A(n17341), .B(n1598), .Z(n1599) );
  NAND U2153 ( .A(n1597), .B(n1599), .Z(n17361) );
  XOR U2154 ( .A(sreg[1738]), .B(n17406), .Z(n1600) );
  NANDN U2155 ( .A(n17407), .B(n1600), .Z(n1601) );
  NAND U2156 ( .A(sreg[1738]), .B(n17406), .Z(n1602) );
  AND U2157 ( .A(n1601), .B(n1602), .Z(n17446) );
  NAND U2158 ( .A(n17496), .B(sreg[1742]), .Z(n1603) );
  XOR U2159 ( .A(sreg[1742]), .B(n17496), .Z(n1604) );
  NANDN U2160 ( .A(n17495), .B(n1604), .Z(n1605) );
  NAND U2161 ( .A(n1603), .B(n1605), .Z(n17531) );
  XOR U2162 ( .A(sreg[1749]), .B(n17651), .Z(n1606) );
  NANDN U2163 ( .A(n17652), .B(n1606), .Z(n1607) );
  NAND U2164 ( .A(sreg[1749]), .B(n17651), .Z(n1608) );
  AND U2165 ( .A(n1607), .B(n1608), .Z(n17673) );
  XOR U2166 ( .A(sreg[1755]), .B(n17785), .Z(n1609) );
  NANDN U2167 ( .A(n17786), .B(n1609), .Z(n1610) );
  NAND U2168 ( .A(sreg[1755]), .B(n17785), .Z(n1611) );
  AND U2169 ( .A(n1610), .B(n1611), .Z(n17825) );
  XOR U2170 ( .A(sreg[1760]), .B(n17898), .Z(n1612) );
  NANDN U2171 ( .A(n17899), .B(n1612), .Z(n1613) );
  NAND U2172 ( .A(sreg[1760]), .B(n17898), .Z(n1614) );
  AND U2173 ( .A(n1613), .B(n1614), .Z(n17938) );
  XOR U2174 ( .A(n18028), .B(n18027), .Z(n1615) );
  NANDN U2175 ( .A(sreg[1765]), .B(n1615), .Z(n1616) );
  NAND U2176 ( .A(n18028), .B(n18027), .Z(n1617) );
  AND U2177 ( .A(n1616), .B(n1617), .Z(n18031) );
  XOR U2178 ( .A(sreg[1769]), .B(n18095), .Z(n1618) );
  NANDN U2179 ( .A(n18096), .B(n1618), .Z(n1619) );
  NAND U2180 ( .A(sreg[1769]), .B(n18095), .Z(n1620) );
  AND U2181 ( .A(n1619), .B(n1620), .Z(n18135) );
  NAND U2182 ( .A(n18207), .B(sreg[1774]), .Z(n1621) );
  XOR U2183 ( .A(sreg[1774]), .B(n18207), .Z(n1622) );
  NANDN U2184 ( .A(n18206), .B(n1622), .Z(n1623) );
  NAND U2185 ( .A(n1621), .B(n1623), .Z(n18245) );
  XOR U2186 ( .A(n18295), .B(sreg[1778]), .Z(n1624) );
  NAND U2187 ( .A(n1624), .B(n18294), .Z(n1625) );
  NAND U2188 ( .A(n18295), .B(sreg[1778]), .Z(n1626) );
  AND U2189 ( .A(n1625), .B(n1626), .Z(n18334) );
  NAND U2190 ( .A(sreg[1783]), .B(n18423), .Z(n1627) );
  XOR U2191 ( .A(n18423), .B(sreg[1783]), .Z(n1628) );
  NANDN U2192 ( .A(n18424), .B(n1628), .Z(n1629) );
  NAND U2193 ( .A(n1627), .B(n1629), .Z(n18444) );
  XOR U2194 ( .A(n18492), .B(n18491), .Z(n1630) );
  NANDN U2195 ( .A(sreg[1787]), .B(n1630), .Z(n1631) );
  NAND U2196 ( .A(n18492), .B(n18491), .Z(n1632) );
  AND U2197 ( .A(n1631), .B(n1632), .Z(n18531) );
  NAND U2198 ( .A(n18597), .B(sreg[1791]), .Z(n1633) );
  XOR U2199 ( .A(sreg[1791]), .B(n18597), .Z(n1634) );
  NAND U2200 ( .A(n1634), .B(n18596), .Z(n1635) );
  NAND U2201 ( .A(n1633), .B(n1635), .Z(n18599) );
  XOR U2202 ( .A(sreg[1795]), .B(n18661), .Z(n1636) );
  NANDN U2203 ( .A(n18662), .B(n1636), .Z(n1637) );
  NAND U2204 ( .A(sreg[1795]), .B(n18661), .Z(n1638) );
  AND U2205 ( .A(n1637), .B(n1638), .Z(n18701) );
  NAND U2206 ( .A(n18794), .B(n18793), .Z(n1639) );
  XOR U2207 ( .A(n18793), .B(n18794), .Z(n1640) );
  NAND U2208 ( .A(n1640), .B(sreg[1801]), .Z(n1641) );
  NAND U2209 ( .A(n1639), .B(n1641), .Z(n18832) );
  XOR U2210 ( .A(sreg[1806]), .B(n18904), .Z(n1642) );
  NANDN U2211 ( .A(n18905), .B(n1642), .Z(n1643) );
  NAND U2212 ( .A(sreg[1806]), .B(n18904), .Z(n1644) );
  AND U2213 ( .A(n1643), .B(n1644), .Z(n18944) );
  NAND U2214 ( .A(n19035), .B(n19034), .Z(n1645) );
  XOR U2215 ( .A(n19034), .B(n19035), .Z(n1646) );
  NAND U2216 ( .A(n1646), .B(sreg[1812]), .Z(n1647) );
  NAND U2217 ( .A(n1645), .B(n1647), .Z(n19073) );
  XOR U2218 ( .A(sreg[1816]), .B(n19122), .Z(n1648) );
  NANDN U2219 ( .A(n19123), .B(n1648), .Z(n1649) );
  NAND U2220 ( .A(sreg[1816]), .B(n19122), .Z(n1650) );
  AND U2221 ( .A(n1649), .B(n1650), .Z(n19143) );
  NAND U2222 ( .A(n19235), .B(n19234), .Z(n1651) );
  XOR U2223 ( .A(n19234), .B(n19235), .Z(n1652) );
  NAND U2224 ( .A(n1652), .B(sreg[1821]), .Z(n1653) );
  NAND U2225 ( .A(n1651), .B(n1653), .Z(n19268) );
  XOR U2226 ( .A(sreg[1826]), .B(n19332), .Z(n1654) );
  NANDN U2227 ( .A(n19333), .B(n1654), .Z(n1655) );
  NAND U2228 ( .A(sreg[1826]), .B(n19332), .Z(n1656) );
  AND U2229 ( .A(n1655), .B(n1656), .Z(n19354) );
  NAND U2230 ( .A(n19421), .B(n19420), .Z(n1657) );
  XOR U2231 ( .A(n19420), .B(n19421), .Z(n1658) );
  NAND U2232 ( .A(n1658), .B(sreg[1830]), .Z(n1659) );
  NAND U2233 ( .A(n1657), .B(n1659), .Z(n19459) );
  XOR U2234 ( .A(sreg[1835]), .B(n19527), .Z(n1660) );
  NANDN U2235 ( .A(n19528), .B(n1660), .Z(n1661) );
  NAND U2236 ( .A(sreg[1835]), .B(n19527), .Z(n1662) );
  AND U2237 ( .A(n1661), .B(n1662), .Z(n19567) );
  XOR U2238 ( .A(sreg[1840]), .B(n19636), .Z(n1663) );
  NANDN U2239 ( .A(n19637), .B(n1663), .Z(n1664) );
  NAND U2240 ( .A(sreg[1840]), .B(n19636), .Z(n1665) );
  AND U2241 ( .A(n1664), .B(n1665), .Z(n19676) );
  NAND U2242 ( .A(sreg[1844]), .B(n19742), .Z(n1666) );
  XOR U2243 ( .A(n19742), .B(sreg[1844]), .Z(n1667) );
  NANDN U2244 ( .A(n19743), .B(n1667), .Z(n1668) );
  NAND U2245 ( .A(n1666), .B(n1668), .Z(n19745) );
  NAND U2246 ( .A(n19811), .B(n19810), .Z(n1669) );
  XOR U2247 ( .A(n19810), .B(n19811), .Z(n1670) );
  NAND U2248 ( .A(n1670), .B(sreg[1848]), .Z(n1671) );
  NAND U2249 ( .A(n1669), .B(n1671), .Z(n19831) );
  XOR U2250 ( .A(sreg[1853]), .B(n19921), .Z(n1672) );
  NANDN U2251 ( .A(n19922), .B(n1672), .Z(n1673) );
  NAND U2252 ( .A(sreg[1853]), .B(n19921), .Z(n1674) );
  AND U2253 ( .A(n1673), .B(n1674), .Z(n19961) );
  NAND U2254 ( .A(n20031), .B(n20030), .Z(n1675) );
  XOR U2255 ( .A(n20030), .B(n20031), .Z(n1676) );
  NAND U2256 ( .A(n1676), .B(sreg[1858]), .Z(n1677) );
  NAND U2257 ( .A(n1675), .B(n1677), .Z(n20069) );
  XOR U2258 ( .A(sreg[1863]), .B(n20141), .Z(n1678) );
  NANDN U2259 ( .A(n20142), .B(n1678), .Z(n1679) );
  NAND U2260 ( .A(sreg[1863]), .B(n20141), .Z(n1680) );
  AND U2261 ( .A(n1679), .B(n1680), .Z(n20180) );
  NAND U2262 ( .A(n20229), .B(sreg[1867]), .Z(n1681) );
  XOR U2263 ( .A(sreg[1867]), .B(n20229), .Z(n1682) );
  NANDN U2264 ( .A(n20230), .B(n1682), .Z(n1683) );
  NAND U2265 ( .A(n1681), .B(n1683), .Z(n20268) );
  XOR U2266 ( .A(sreg[1872]), .B(n20338), .Z(n1684) );
  NANDN U2267 ( .A(n20339), .B(n1684), .Z(n1685) );
  NAND U2268 ( .A(sreg[1872]), .B(n20338), .Z(n1686) );
  AND U2269 ( .A(n1685), .B(n1686), .Z(n20378) );
  NAND U2270 ( .A(n20491), .B(n20490), .Z(n1687) );
  XOR U2271 ( .A(n20490), .B(n20491), .Z(n1688) );
  NAND U2272 ( .A(n1688), .B(sreg[1878]), .Z(n1689) );
  NAND U2273 ( .A(n1687), .B(n1689), .Z(n20493) );
  XOR U2274 ( .A(sreg[1882]), .B(n20561), .Z(n1690) );
  NANDN U2275 ( .A(n20562), .B(n1690), .Z(n1691) );
  NAND U2276 ( .A(sreg[1882]), .B(n20561), .Z(n1692) );
  AND U2277 ( .A(n1691), .B(n1692), .Z(n20596) );
  NAND U2278 ( .A(n20661), .B(sreg[1886]), .Z(n1693) );
  XOR U2279 ( .A(sreg[1886]), .B(n20661), .Z(n1694) );
  NAND U2280 ( .A(n1694), .B(n20660), .Z(n1695) );
  NAND U2281 ( .A(n1693), .B(n1695), .Z(n20682) );
  XOR U2282 ( .A(n20725), .B(sreg[1890]), .Z(n1696) );
  NAND U2283 ( .A(n1696), .B(n20724), .Z(n1697) );
  NAND U2284 ( .A(n20725), .B(sreg[1890]), .Z(n1698) );
  AND U2285 ( .A(n1697), .B(n1698), .Z(n20763) );
  NAND U2286 ( .A(n20834), .B(n20833), .Z(n1699) );
  XOR U2287 ( .A(n20833), .B(n20834), .Z(n1700) );
  NAND U2288 ( .A(n1700), .B(sreg[1895]), .Z(n1701) );
  NAND U2289 ( .A(n1699), .B(n1701), .Z(n20872) );
  XOR U2290 ( .A(sreg[1900]), .B(n20942), .Z(n1702) );
  NANDN U2291 ( .A(n20943), .B(n1702), .Z(n1703) );
  NAND U2292 ( .A(sreg[1900]), .B(n20942), .Z(n1704) );
  AND U2293 ( .A(n1703), .B(n1704), .Z(n20982) );
  NAND U2294 ( .A(n21072), .B(n21071), .Z(n1705) );
  XOR U2295 ( .A(n21071), .B(n21072), .Z(n1706) );
  NAND U2296 ( .A(n1706), .B(sreg[1905]), .Z(n1707) );
  NAND U2297 ( .A(n1705), .B(n1707), .Z(n21074) );
  NAND U2298 ( .A(n21140), .B(n21139), .Z(n1708) );
  XOR U2299 ( .A(n21139), .B(n21140), .Z(n1709) );
  NAND U2300 ( .A(n1709), .B(sreg[1909]), .Z(n1710) );
  NAND U2301 ( .A(n1708), .B(n1710), .Z(n21178) );
  NAND U2302 ( .A(sreg[1914]), .B(n21266), .Z(n1711) );
  XOR U2303 ( .A(n21266), .B(sreg[1914]), .Z(n1712) );
  NANDN U2304 ( .A(n21267), .B(n1712), .Z(n1713) );
  NAND U2305 ( .A(n1711), .B(n1713), .Z(n21287) );
  XOR U2306 ( .A(sreg[1918]), .B(n21334), .Z(n1714) );
  NANDN U2307 ( .A(n21335), .B(n1714), .Z(n1715) );
  NAND U2308 ( .A(sreg[1918]), .B(n21334), .Z(n1716) );
  AND U2309 ( .A(n1715), .B(n1716), .Z(n21374) );
  XOR U2310 ( .A(sreg[1923]), .B(n21443), .Z(n1717) );
  NANDN U2311 ( .A(n21444), .B(n1717), .Z(n1718) );
  NAND U2312 ( .A(sreg[1923]), .B(n21443), .Z(n1719) );
  AND U2313 ( .A(n1718), .B(n1719), .Z(n21483) );
  XOR U2314 ( .A(n21569), .B(n21568), .Z(n1720) );
  NANDN U2315 ( .A(sreg[1928]), .B(n1720), .Z(n1721) );
  NAND U2316 ( .A(n21569), .B(n21568), .Z(n1722) );
  AND U2317 ( .A(n1721), .B(n1722), .Z(n21571) );
  XOR U2318 ( .A(sreg[1932]), .B(n21638), .Z(n1723) );
  NANDN U2319 ( .A(n21639), .B(n1723), .Z(n1724) );
  NAND U2320 ( .A(sreg[1932]), .B(n21638), .Z(n1725) );
  AND U2321 ( .A(n1724), .B(n1725), .Z(n21679) );
  XOR U2322 ( .A(n21750), .B(sreg[1937]), .Z(n1726) );
  NAND U2323 ( .A(n1726), .B(n21749), .Z(n1727) );
  NAND U2324 ( .A(n21750), .B(sreg[1937]), .Z(n1728) );
  AND U2325 ( .A(n1727), .B(n1728), .Z(n21789) );
  XOR U2326 ( .A(n21838), .B(sreg[1941]), .Z(n1729) );
  NAND U2327 ( .A(n1729), .B(n21837), .Z(n1730) );
  NAND U2328 ( .A(n21838), .B(sreg[1941]), .Z(n1731) );
  AND U2329 ( .A(n1730), .B(n1731), .Z(n21858) );
  NAND U2330 ( .A(sreg[1946]), .B(n21966), .Z(n1732) );
  XOR U2331 ( .A(n21966), .B(sreg[1946]), .Z(n1733) );
  NANDN U2332 ( .A(n21967), .B(n1733), .Z(n1734) );
  NAND U2333 ( .A(n1732), .B(n1734), .Z(n21969) );
  NAND U2334 ( .A(n22036), .B(n22035), .Z(n1735) );
  XOR U2335 ( .A(n22035), .B(n22036), .Z(n1736) );
  NAND U2336 ( .A(n1736), .B(sreg[1950]), .Z(n1737) );
  NAND U2337 ( .A(n1735), .B(n1737), .Z(n22071) );
  XOR U2338 ( .A(n22180), .B(sreg[1956]), .Z(n1738) );
  NANDN U2339 ( .A(n22181), .B(n1738), .Z(n1739) );
  NAND U2340 ( .A(n22180), .B(sreg[1956]), .Z(n1740) );
  AND U2341 ( .A(n1739), .B(n1740), .Z(n22201) );
  XOR U2342 ( .A(sreg[1962]), .B(n22294), .Z(n1741) );
  NANDN U2343 ( .A(n22295), .B(n1741), .Z(n1742) );
  NAND U2344 ( .A(sreg[1962]), .B(n22294), .Z(n1743) );
  AND U2345 ( .A(n1742), .B(n1743), .Z(n22315) );
  XOR U2346 ( .A(sreg[1967]), .B(n22407), .Z(n1744) );
  NANDN U2347 ( .A(n22408), .B(n1744), .Z(n1745) );
  NAND U2348 ( .A(sreg[1967]), .B(n22407), .Z(n1746) );
  AND U2349 ( .A(n1745), .B(n1746), .Z(n22447) );
  NAND U2350 ( .A(n22542), .B(n22541), .Z(n1747) );
  XOR U2351 ( .A(n22541), .B(n22542), .Z(n1748) );
  NAND U2352 ( .A(n1748), .B(sreg[1973]), .Z(n1749) );
  NAND U2353 ( .A(n1747), .B(n1749), .Z(n22580) );
  XOR U2354 ( .A(sreg[1977]), .B(n22629), .Z(n1750) );
  NANDN U2355 ( .A(n22630), .B(n1750), .Z(n1751) );
  NAND U2356 ( .A(sreg[1977]), .B(n22629), .Z(n1752) );
  AND U2357 ( .A(n1751), .B(n1752), .Z(n22669) );
  XOR U2358 ( .A(sreg[1982]), .B(n22740), .Z(n1753) );
  NANDN U2359 ( .A(n22741), .B(n1753), .Z(n1754) );
  NAND U2360 ( .A(sreg[1982]), .B(n22740), .Z(n1755) );
  AND U2361 ( .A(n1754), .B(n1755), .Z(n22780) );
  XOR U2362 ( .A(n22829), .B(sreg[1986]), .Z(n1756) );
  NAND U2363 ( .A(n1756), .B(n22828), .Z(n1757) );
  NAND U2364 ( .A(n22829), .B(sreg[1986]), .Z(n1758) );
  AND U2365 ( .A(n1757), .B(n1758), .Z(n22849) );
  NAND U2366 ( .A(n22935), .B(n22934), .Z(n1759) );
  XOR U2367 ( .A(n22934), .B(n22935), .Z(n1760) );
  NAND U2368 ( .A(n1760), .B(sreg[1990]), .Z(n1761) );
  NAND U2369 ( .A(n1759), .B(n1761), .Z(n22955) );
  NAND U2370 ( .A(sreg[1994]), .B(n23020), .Z(n1762) );
  XOR U2371 ( .A(n23020), .B(sreg[1994]), .Z(n1763) );
  NANDN U2372 ( .A(n23021), .B(n1763), .Z(n1764) );
  NAND U2373 ( .A(n1762), .B(n1764), .Z(n23023) );
  XOR U2374 ( .A(n23089), .B(sreg[1998]), .Z(n1765) );
  NAND U2375 ( .A(n1765), .B(n23088), .Z(n1766) );
  NAND U2376 ( .A(n23089), .B(sreg[1998]), .Z(n1767) );
  AND U2377 ( .A(n1766), .B(n1767), .Z(n23129) );
  XOR U2378 ( .A(n23173), .B(sreg[2002]), .Z(n1768) );
  NANDN U2379 ( .A(n23172), .B(n1768), .Z(n1769) );
  NAND U2380 ( .A(n23173), .B(sreg[2002]), .Z(n1770) );
  AND U2381 ( .A(n1769), .B(n1770), .Z(n23194) );
  XOR U2382 ( .A(sreg[2007]), .B(n23281), .Z(n1771) );
  NANDN U2383 ( .A(n23282), .B(n1771), .Z(n1772) );
  NAND U2384 ( .A(sreg[2007]), .B(n23281), .Z(n1773) );
  AND U2385 ( .A(n1772), .B(n1773), .Z(n23321) );
  XOR U2386 ( .A(sreg[2012]), .B(n23392), .Z(n1774) );
  NANDN U2387 ( .A(n23393), .B(n1774), .Z(n1775) );
  NAND U2388 ( .A(sreg[2012]), .B(n23392), .Z(n1776) );
  AND U2389 ( .A(n1775), .B(n1776), .Z(n23413) );
  NAND U2390 ( .A(n23522), .B(n23521), .Z(n1777) );
  XOR U2391 ( .A(n23521), .B(n23522), .Z(n1778) );
  NAND U2392 ( .A(n1778), .B(sreg[2017]), .Z(n1779) );
  NAND U2393 ( .A(n1777), .B(n1779), .Z(n23524) );
  XOR U2394 ( .A(n23608), .B(n23607), .Z(n1780) );
  NANDN U2395 ( .A(sreg[2021]), .B(n1780), .Z(n1781) );
  NAND U2396 ( .A(n23608), .B(n23607), .Z(n1782) );
  AND U2397 ( .A(n1781), .B(n1782), .Z(n23610) );
  NAND U2398 ( .A(sreg[2025]), .B(n23693), .Z(n1783) );
  XOR U2399 ( .A(n23693), .B(sreg[2025]), .Z(n1784) );
  NANDN U2400 ( .A(n23694), .B(n1784), .Z(n1785) );
  NAND U2401 ( .A(n1783), .B(n1785), .Z(n23696) );
  XOR U2402 ( .A(sreg[2029]), .B(n23763), .Z(n1786) );
  NANDN U2403 ( .A(n23764), .B(n1786), .Z(n1787) );
  NAND U2404 ( .A(sreg[2029]), .B(n23763), .Z(n1788) );
  AND U2405 ( .A(n1787), .B(n1788), .Z(n23803) );
  XOR U2406 ( .A(sreg[2034]), .B(n23874), .Z(n1789) );
  NANDN U2407 ( .A(n23875), .B(n1789), .Z(n1790) );
  NAND U2408 ( .A(sreg[2034]), .B(n23874), .Z(n1791) );
  AND U2409 ( .A(n1790), .B(n1791), .Z(n23914) );
  NAND U2410 ( .A(n24032), .B(n24031), .Z(n1792) );
  XOR U2411 ( .A(n24031), .B(n24032), .Z(n1793) );
  NAND U2412 ( .A(n1793), .B(sreg[2041]), .Z(n1794) );
  NAND U2413 ( .A(n1792), .B(n1794), .Z(n24049) );
  IV U2414 ( .A(b[1]), .Z(n1795) );
  IV U2415 ( .A(b[3]), .Z(n1796) );
  NAND U2416 ( .A(b[0]), .B(a[0]), .Z(n1804) );
  XNOR U2417 ( .A(n1804), .B(sreg[1020]), .Z(c[1020]) );
  AND U2418 ( .A(a[1]), .B(b[0]), .Z(n1798) );
  NAND U2419 ( .A(b[1]), .B(a[0]), .Z(n1797) );
  XNOR U2420 ( .A(n1798), .B(n1797), .Z(n1799) );
  XNOR U2421 ( .A(sreg[1021]), .B(n1799), .Z(n1801) );
  NANDN U2422 ( .A(n1804), .B(sreg[1020]), .Z(n1800) );
  XOR U2423 ( .A(n1801), .B(n1800), .Z(c[1021]) );
  NAND U2424 ( .A(n1799), .B(sreg[1021]), .Z(n1803) );
  OR U2425 ( .A(n1801), .B(n1800), .Z(n1802) );
  AND U2426 ( .A(n1803), .B(n1802), .Z(n1815) );
  ANDN U2427 ( .B(a[1]), .A(n1795), .Z(n1826) );
  ANDN U2428 ( .B(n1826), .A(n1804), .Z(n1811) );
  AND U2429 ( .A(b[2]), .B(a[0]), .Z(n1809) );
  NAND U2430 ( .A(b[0]), .B(a[2]), .Z(n1827) );
  XOR U2431 ( .A(n1827), .B(n1826), .Z(n1808) );
  XNOR U2432 ( .A(n1809), .B(n1808), .Z(n1810) );
  XOR U2433 ( .A(n1811), .B(n1810), .Z(n1814) );
  XNOR U2434 ( .A(sreg[1022]), .B(n1814), .Z(n1805) );
  XOR U2435 ( .A(n1815), .B(n1805), .Z(c[1022]) );
  ANDN U2436 ( .B(a[2]), .A(n1843), .Z(n1806) );
  NAND U2437 ( .A(b[1]), .B(n1806), .Z(n1829) );
  NAND U2438 ( .A(b[3]), .B(a[0]), .Z(n1828) );
  XOR U2439 ( .A(n1829), .B(n1828), .Z(n1816) );
  AND U2440 ( .A(a[3]), .B(b[0]), .Z(n1850) );
  NAND U2441 ( .A(b[2]), .B(a[1]), .Z(n1807) );
  XNOR U2442 ( .A(n1850), .B(n1807), .Z(n1817) );
  XNOR U2443 ( .A(n1816), .B(n1817), .Z(n1819) );
  NANDN U2444 ( .A(n1809), .B(n1808), .Z(n1813) );
  NANDN U2445 ( .A(n1811), .B(n1810), .Z(n1812) );
  AND U2446 ( .A(n1813), .B(n1812), .Z(n1818) );
  XNOR U2447 ( .A(n1819), .B(n1818), .Z(n1833) );
  XNOR U2448 ( .A(n1832), .B(sreg[1023]), .Z(n1834) );
  XNOR U2449 ( .A(n1833), .B(n1834), .Z(c[1023]) );
  NAND U2450 ( .A(n1817), .B(n1816), .Z(n1821) );
  NANDN U2451 ( .A(n1819), .B(n1818), .Z(n1820) );
  NAND U2452 ( .A(n1821), .B(n1820), .Z(n1840) );
  AND U2453 ( .A(b[2]), .B(a[3]), .Z(n1870) );
  NAND U2454 ( .A(b[0]), .B(n1870), .Z(n1822) );
  XNOR U2455 ( .A(b[3]), .B(n1822), .Z(n1823) );
  NAND U2456 ( .A(a[1]), .B(n1823), .Z(n1847) );
  XNOR U2457 ( .A(n1846), .B(n1847), .Z(n1852) );
  AND U2458 ( .A(a[4]), .B(b[0]), .Z(n1825) );
  NAND U2459 ( .A(b[1]), .B(a[3]), .Z(n1824) );
  XNOR U2460 ( .A(n1825), .B(n1824), .Z(n1851) );
  XNOR U2461 ( .A(n1852), .B(n1851), .Z(n1837) );
  NANDN U2462 ( .A(n1827), .B(n1826), .Z(n1831) );
  OR U2463 ( .A(n1829), .B(n1828), .Z(n1830) );
  NAND U2464 ( .A(n1831), .B(n1830), .Z(n1838) );
  XOR U2465 ( .A(n1837), .B(n1838), .Z(n1839) );
  XOR U2466 ( .A(n1840), .B(n1839), .Z(n1855) );
  XNOR U2467 ( .A(n1855), .B(sreg[1024]), .Z(n1857) );
  NAND U2468 ( .A(n1832), .B(sreg[1023]), .Z(n1836) );
  NANDN U2469 ( .A(n1834), .B(n1833), .Z(n1835) );
  AND U2470 ( .A(n1836), .B(n1835), .Z(n1856) );
  XOR U2471 ( .A(n1857), .B(n1856), .Z(c[1024]) );
  OR U2472 ( .A(n1838), .B(n1837), .Z(n1842) );
  NANDN U2473 ( .A(n1840), .B(n1839), .Z(n1841) );
  NAND U2474 ( .A(n1842), .B(n1841), .Z(n1864) );
  ANDN U2475 ( .B(a[4]), .A(n1795), .Z(n1867) );
  AND U2476 ( .A(b[3]), .B(a[2]), .Z(n1868) );
  XNOR U2477 ( .A(n1870), .B(n1869), .Z(n1873) );
  NAND U2478 ( .A(b[0]), .B(a[5]), .Z(n1874) );
  XOR U2479 ( .A(n1873), .B(n1874), .Z(n1875) );
  NAND U2480 ( .A(n1870), .B(n1843), .Z(n1845) );
  NAND U2481 ( .A(b[3]), .B(a[1]), .Z(n1844) );
  AND U2482 ( .A(n1845), .B(n1844), .Z(n1849) );
  NANDN U2483 ( .A(n1847), .B(n1846), .Z(n1848) );
  NANDN U2484 ( .A(n1849), .B(n1848), .Z(n1876) );
  XOR U2485 ( .A(n1875), .B(n1876), .Z(n1861) );
  NAND U2486 ( .A(n1867), .B(n1850), .Z(n1854) );
  NANDN U2487 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U2488 ( .A(n1854), .B(n1853), .Z(n1862) );
  XNOR U2489 ( .A(n1861), .B(n1862), .Z(n1863) );
  XNOR U2490 ( .A(n1864), .B(n1863), .Z(n1880) );
  NAND U2491 ( .A(n1855), .B(sreg[1024]), .Z(n1859) );
  OR U2492 ( .A(n1857), .B(n1856), .Z(n1858) );
  AND U2493 ( .A(n1859), .B(n1858), .Z(n1879) );
  XNOR U2494 ( .A(n1879), .B(sreg[1025]), .Z(n1860) );
  XOR U2495 ( .A(n1880), .B(n1860), .Z(c[1025]) );
  NANDN U2496 ( .A(n1862), .B(n1861), .Z(n1866) );
  NAND U2497 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2498 ( .A(n1866), .B(n1865), .Z(n1885) );
  AND U2499 ( .A(b[2]), .B(a[4]), .Z(n1891) );
  AND U2500 ( .A(a[5]), .B(b[1]), .Z(n1889) );
  AND U2501 ( .A(a[3]), .B(b[3]), .Z(n1888) );
  XOR U2502 ( .A(n1889), .B(n1888), .Z(n1890) );
  XOR U2503 ( .A(n1891), .B(n1890), .Z(n1894) );
  NAND U2504 ( .A(b[0]), .B(a[6]), .Z(n1895) );
  XOR U2505 ( .A(n1894), .B(n1895), .Z(n1897) );
  OR U2506 ( .A(n1868), .B(n1867), .Z(n1872) );
  NANDN U2507 ( .A(n1870), .B(n1869), .Z(n1871) );
  NAND U2508 ( .A(n1872), .B(n1871), .Z(n1896) );
  XNOR U2509 ( .A(n1897), .B(n1896), .Z(n1882) );
  OR U2510 ( .A(n1874), .B(n1873), .Z(n1878) );
  NANDN U2511 ( .A(n1876), .B(n1875), .Z(n1877) );
  NAND U2512 ( .A(n1878), .B(n1877), .Z(n1883) );
  XNOR U2513 ( .A(n1882), .B(n1883), .Z(n1884) );
  XOR U2514 ( .A(n1885), .B(n1884), .Z(n1901) );
  XOR U2515 ( .A(sreg[1026]), .B(n1900), .Z(n1881) );
  XOR U2516 ( .A(n1901), .B(n1881), .Z(c[1026]) );
  NANDN U2517 ( .A(n1883), .B(n1882), .Z(n1887) );
  NAND U2518 ( .A(n1885), .B(n1884), .Z(n1886) );
  NAND U2519 ( .A(n1887), .B(n1886), .Z(n1908) );
  AND U2520 ( .A(b[2]), .B(a[5]), .Z(n1914) );
  AND U2521 ( .A(a[6]), .B(b[1]), .Z(n1912) );
  AND U2522 ( .A(a[4]), .B(b[3]), .Z(n1911) );
  XOR U2523 ( .A(n1912), .B(n1911), .Z(n1913) );
  XOR U2524 ( .A(n1914), .B(n1913), .Z(n1917) );
  NAND U2525 ( .A(b[0]), .B(a[7]), .Z(n1918) );
  XOR U2526 ( .A(n1917), .B(n1918), .Z(n1920) );
  OR U2527 ( .A(n1889), .B(n1888), .Z(n1893) );
  NANDN U2528 ( .A(n1891), .B(n1890), .Z(n1892) );
  NAND U2529 ( .A(n1893), .B(n1892), .Z(n1919) );
  XNOR U2530 ( .A(n1920), .B(n1919), .Z(n1905) );
  NANDN U2531 ( .A(n1895), .B(n1894), .Z(n1899) );
  OR U2532 ( .A(n1897), .B(n1896), .Z(n1898) );
  NAND U2533 ( .A(n1899), .B(n1898), .Z(n1906) );
  XNOR U2534 ( .A(n1905), .B(n1906), .Z(n1907) );
  XOR U2535 ( .A(n1908), .B(n1907), .Z(n1904) );
  XNOR U2536 ( .A(sreg[1027]), .B(n1903), .Z(n1902) );
  XOR U2537 ( .A(n1904), .B(n1902), .Z(c[1027]) );
  NANDN U2538 ( .A(n1906), .B(n1905), .Z(n1910) );
  NAND U2539 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U2540 ( .A(n1910), .B(n1909), .Z(n1926) );
  AND U2541 ( .A(b[2]), .B(a[6]), .Z(n1932) );
  AND U2542 ( .A(a[7]), .B(b[1]), .Z(n1930) );
  AND U2543 ( .A(a[5]), .B(b[3]), .Z(n1929) );
  XOR U2544 ( .A(n1930), .B(n1929), .Z(n1931) );
  XOR U2545 ( .A(n1932), .B(n1931), .Z(n1935) );
  NAND U2546 ( .A(b[0]), .B(a[8]), .Z(n1936) );
  XOR U2547 ( .A(n1935), .B(n1936), .Z(n1938) );
  OR U2548 ( .A(n1912), .B(n1911), .Z(n1916) );
  NANDN U2549 ( .A(n1914), .B(n1913), .Z(n1915) );
  NAND U2550 ( .A(n1916), .B(n1915), .Z(n1937) );
  XNOR U2551 ( .A(n1938), .B(n1937), .Z(n1923) );
  NANDN U2552 ( .A(n1918), .B(n1917), .Z(n1922) );
  OR U2553 ( .A(n1920), .B(n1919), .Z(n1921) );
  NAND U2554 ( .A(n1922), .B(n1921), .Z(n1924) );
  XNOR U2555 ( .A(n1923), .B(n1924), .Z(n1925) );
  XNOR U2556 ( .A(n1926), .B(n1925), .Z(n1941) );
  XNOR U2557 ( .A(n1941), .B(sreg[1028]), .Z(n1942) );
  XOR U2558 ( .A(n1943), .B(n1942), .Z(c[1028]) );
  NANDN U2559 ( .A(n1924), .B(n1923), .Z(n1928) );
  NAND U2560 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2561 ( .A(n1928), .B(n1927), .Z(n1949) );
  AND U2562 ( .A(b[2]), .B(a[7]), .Z(n1955) );
  AND U2563 ( .A(a[8]), .B(b[1]), .Z(n1953) );
  AND U2564 ( .A(a[6]), .B(b[3]), .Z(n1952) );
  XOR U2565 ( .A(n1953), .B(n1952), .Z(n1954) );
  XOR U2566 ( .A(n1955), .B(n1954), .Z(n1958) );
  NAND U2567 ( .A(b[0]), .B(a[9]), .Z(n1959) );
  XOR U2568 ( .A(n1958), .B(n1959), .Z(n1961) );
  OR U2569 ( .A(n1930), .B(n1929), .Z(n1934) );
  NANDN U2570 ( .A(n1932), .B(n1931), .Z(n1933) );
  NAND U2571 ( .A(n1934), .B(n1933), .Z(n1960) );
  XNOR U2572 ( .A(n1961), .B(n1960), .Z(n1946) );
  NANDN U2573 ( .A(n1936), .B(n1935), .Z(n1940) );
  OR U2574 ( .A(n1938), .B(n1937), .Z(n1939) );
  NAND U2575 ( .A(n1940), .B(n1939), .Z(n1947) );
  XNOR U2576 ( .A(n1946), .B(n1947), .Z(n1948) );
  XNOR U2577 ( .A(n1949), .B(n1948), .Z(n1964) );
  XNOR U2578 ( .A(n1964), .B(sreg[1029]), .Z(n1966) );
  NAND U2579 ( .A(n1941), .B(sreg[1028]), .Z(n1945) );
  OR U2580 ( .A(n1943), .B(n1942), .Z(n1944) );
  AND U2581 ( .A(n1945), .B(n1944), .Z(n1965) );
  XOR U2582 ( .A(n1966), .B(n1965), .Z(c[1029]) );
  NANDN U2583 ( .A(n1947), .B(n1946), .Z(n1951) );
  NAND U2584 ( .A(n1949), .B(n1948), .Z(n1950) );
  NAND U2585 ( .A(n1951), .B(n1950), .Z(n1973) );
  AND U2586 ( .A(b[2]), .B(a[8]), .Z(n1979) );
  AND U2587 ( .A(a[9]), .B(b[1]), .Z(n1977) );
  AND U2588 ( .A(a[7]), .B(b[3]), .Z(n1976) );
  XOR U2589 ( .A(n1977), .B(n1976), .Z(n1978) );
  XOR U2590 ( .A(n1979), .B(n1978), .Z(n1982) );
  NAND U2591 ( .A(b[0]), .B(a[10]), .Z(n1983) );
  XOR U2592 ( .A(n1982), .B(n1983), .Z(n1985) );
  OR U2593 ( .A(n1953), .B(n1952), .Z(n1957) );
  NANDN U2594 ( .A(n1955), .B(n1954), .Z(n1956) );
  NAND U2595 ( .A(n1957), .B(n1956), .Z(n1984) );
  XNOR U2596 ( .A(n1985), .B(n1984), .Z(n1970) );
  NANDN U2597 ( .A(n1959), .B(n1958), .Z(n1963) );
  OR U2598 ( .A(n1961), .B(n1960), .Z(n1962) );
  NAND U2599 ( .A(n1963), .B(n1962), .Z(n1971) );
  XNOR U2600 ( .A(n1970), .B(n1971), .Z(n1972) );
  XOR U2601 ( .A(n1973), .B(n1972), .Z(n1989) );
  NAND U2602 ( .A(n1964), .B(sreg[1029]), .Z(n1968) );
  OR U2603 ( .A(n1966), .B(n1965), .Z(n1967) );
  NAND U2604 ( .A(n1968), .B(n1967), .Z(n1988) );
  XNOR U2605 ( .A(sreg[1030]), .B(n1988), .Z(n1969) );
  XOR U2606 ( .A(n1989), .B(n1969), .Z(c[1030]) );
  NANDN U2607 ( .A(n1971), .B(n1970), .Z(n1975) );
  NAND U2608 ( .A(n1973), .B(n1972), .Z(n1974) );
  NAND U2609 ( .A(n1975), .B(n1974), .Z(n1996) );
  AND U2610 ( .A(b[2]), .B(a[9]), .Z(n2002) );
  AND U2611 ( .A(a[10]), .B(b[1]), .Z(n2000) );
  AND U2612 ( .A(a[8]), .B(b[3]), .Z(n1999) );
  XOR U2613 ( .A(n2000), .B(n1999), .Z(n2001) );
  XOR U2614 ( .A(n2002), .B(n2001), .Z(n2005) );
  NAND U2615 ( .A(b[0]), .B(a[11]), .Z(n2006) );
  XOR U2616 ( .A(n2005), .B(n2006), .Z(n2008) );
  OR U2617 ( .A(n1977), .B(n1976), .Z(n1981) );
  NANDN U2618 ( .A(n1979), .B(n1978), .Z(n1980) );
  NAND U2619 ( .A(n1981), .B(n1980), .Z(n2007) );
  XNOR U2620 ( .A(n2008), .B(n2007), .Z(n1993) );
  NANDN U2621 ( .A(n1983), .B(n1982), .Z(n1987) );
  OR U2622 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U2623 ( .A(n1987), .B(n1986), .Z(n1994) );
  XNOR U2624 ( .A(n1993), .B(n1994), .Z(n1995) );
  XNOR U2625 ( .A(n1996), .B(n1995), .Z(n1992) );
  XOR U2626 ( .A(n1991), .B(sreg[1031]), .Z(n1990) );
  XOR U2627 ( .A(n1992), .B(n1990), .Z(c[1031]) );
  NANDN U2628 ( .A(n1994), .B(n1993), .Z(n1998) );
  NAND U2629 ( .A(n1996), .B(n1995), .Z(n1997) );
  NAND U2630 ( .A(n1998), .B(n1997), .Z(n2014) );
  AND U2631 ( .A(b[2]), .B(a[10]), .Z(n2020) );
  AND U2632 ( .A(a[11]), .B(b[1]), .Z(n2018) );
  AND U2633 ( .A(a[9]), .B(b[3]), .Z(n2017) );
  XOR U2634 ( .A(n2018), .B(n2017), .Z(n2019) );
  XOR U2635 ( .A(n2020), .B(n2019), .Z(n2023) );
  NAND U2636 ( .A(b[0]), .B(a[12]), .Z(n2024) );
  XOR U2637 ( .A(n2023), .B(n2024), .Z(n2026) );
  OR U2638 ( .A(n2000), .B(n1999), .Z(n2004) );
  NANDN U2639 ( .A(n2002), .B(n2001), .Z(n2003) );
  NAND U2640 ( .A(n2004), .B(n2003), .Z(n2025) );
  XNOR U2641 ( .A(n2026), .B(n2025), .Z(n2011) );
  NANDN U2642 ( .A(n2006), .B(n2005), .Z(n2010) );
  OR U2643 ( .A(n2008), .B(n2007), .Z(n2009) );
  NAND U2644 ( .A(n2010), .B(n2009), .Z(n2012) );
  XNOR U2645 ( .A(n2011), .B(n2012), .Z(n2013) );
  XNOR U2646 ( .A(n2014), .B(n2013), .Z(n2029) );
  XNOR U2647 ( .A(n2029), .B(sreg[1032]), .Z(n2031) );
  XNOR U2648 ( .A(n2030), .B(n2031), .Z(c[1032]) );
  NANDN U2649 ( .A(n2012), .B(n2011), .Z(n2016) );
  NAND U2650 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U2651 ( .A(n2016), .B(n2015), .Z(n2040) );
  AND U2652 ( .A(b[2]), .B(a[11]), .Z(n2046) );
  AND U2653 ( .A(a[12]), .B(b[1]), .Z(n2044) );
  AND U2654 ( .A(a[10]), .B(b[3]), .Z(n2043) );
  XOR U2655 ( .A(n2044), .B(n2043), .Z(n2045) );
  XOR U2656 ( .A(n2046), .B(n2045), .Z(n2049) );
  NAND U2657 ( .A(b[0]), .B(a[13]), .Z(n2050) );
  XOR U2658 ( .A(n2049), .B(n2050), .Z(n2052) );
  OR U2659 ( .A(n2018), .B(n2017), .Z(n2022) );
  NANDN U2660 ( .A(n2020), .B(n2019), .Z(n2021) );
  NAND U2661 ( .A(n2022), .B(n2021), .Z(n2051) );
  XNOR U2662 ( .A(n2052), .B(n2051), .Z(n2037) );
  NANDN U2663 ( .A(n2024), .B(n2023), .Z(n2028) );
  OR U2664 ( .A(n2026), .B(n2025), .Z(n2027) );
  NAND U2665 ( .A(n2028), .B(n2027), .Z(n2038) );
  XNOR U2666 ( .A(n2037), .B(n2038), .Z(n2039) );
  XNOR U2667 ( .A(n2040), .B(n2039), .Z(n2036) );
  NAND U2668 ( .A(n2029), .B(sreg[1032]), .Z(n2033) );
  NANDN U2669 ( .A(n2031), .B(n2030), .Z(n2032) );
  AND U2670 ( .A(n2033), .B(n2032), .Z(n2035) );
  XNOR U2671 ( .A(n2035), .B(sreg[1033]), .Z(n2034) );
  XOR U2672 ( .A(n2036), .B(n2034), .Z(c[1033]) );
  NANDN U2673 ( .A(n2038), .B(n2037), .Z(n2042) );
  NAND U2674 ( .A(n2040), .B(n2039), .Z(n2041) );
  NAND U2675 ( .A(n2042), .B(n2041), .Z(n2058) );
  AND U2676 ( .A(b[2]), .B(a[12]), .Z(n2064) );
  AND U2677 ( .A(a[13]), .B(b[1]), .Z(n2062) );
  AND U2678 ( .A(a[11]), .B(b[3]), .Z(n2061) );
  XOR U2679 ( .A(n2062), .B(n2061), .Z(n2063) );
  XOR U2680 ( .A(n2064), .B(n2063), .Z(n2067) );
  NAND U2681 ( .A(b[0]), .B(a[14]), .Z(n2068) );
  XOR U2682 ( .A(n2067), .B(n2068), .Z(n2070) );
  OR U2683 ( .A(n2044), .B(n2043), .Z(n2048) );
  NANDN U2684 ( .A(n2046), .B(n2045), .Z(n2047) );
  NAND U2685 ( .A(n2048), .B(n2047), .Z(n2069) );
  XNOR U2686 ( .A(n2070), .B(n2069), .Z(n2055) );
  NANDN U2687 ( .A(n2050), .B(n2049), .Z(n2054) );
  OR U2688 ( .A(n2052), .B(n2051), .Z(n2053) );
  NAND U2689 ( .A(n2054), .B(n2053), .Z(n2056) );
  XNOR U2690 ( .A(n2055), .B(n2056), .Z(n2057) );
  XNOR U2691 ( .A(n2058), .B(n2057), .Z(n2073) );
  XNOR U2692 ( .A(n2073), .B(sreg[1034]), .Z(n2075) );
  XNOR U2693 ( .A(n2074), .B(n2075), .Z(c[1034]) );
  NANDN U2694 ( .A(n2056), .B(n2055), .Z(n2060) );
  NAND U2695 ( .A(n2058), .B(n2057), .Z(n2059) );
  NAND U2696 ( .A(n2060), .B(n2059), .Z(n2081) );
  AND U2697 ( .A(b[2]), .B(a[13]), .Z(n2087) );
  AND U2698 ( .A(a[14]), .B(b[1]), .Z(n2085) );
  AND U2699 ( .A(a[12]), .B(b[3]), .Z(n2084) );
  XOR U2700 ( .A(n2085), .B(n2084), .Z(n2086) );
  XOR U2701 ( .A(n2087), .B(n2086), .Z(n2090) );
  NAND U2702 ( .A(b[0]), .B(a[15]), .Z(n2091) );
  XOR U2703 ( .A(n2090), .B(n2091), .Z(n2093) );
  OR U2704 ( .A(n2062), .B(n2061), .Z(n2066) );
  NANDN U2705 ( .A(n2064), .B(n2063), .Z(n2065) );
  NAND U2706 ( .A(n2066), .B(n2065), .Z(n2092) );
  XNOR U2707 ( .A(n2093), .B(n2092), .Z(n2078) );
  NANDN U2708 ( .A(n2068), .B(n2067), .Z(n2072) );
  OR U2709 ( .A(n2070), .B(n2069), .Z(n2071) );
  NAND U2710 ( .A(n2072), .B(n2071), .Z(n2079) );
  XNOR U2711 ( .A(n2078), .B(n2079), .Z(n2080) );
  XNOR U2712 ( .A(n2081), .B(n2080), .Z(n2096) );
  XNOR U2713 ( .A(n2096), .B(sreg[1035]), .Z(n2098) );
  NAND U2714 ( .A(n2073), .B(sreg[1034]), .Z(n2077) );
  NANDN U2715 ( .A(n2075), .B(n2074), .Z(n2076) );
  AND U2716 ( .A(n2077), .B(n2076), .Z(n2097) );
  XOR U2717 ( .A(n2098), .B(n2097), .Z(c[1035]) );
  NANDN U2718 ( .A(n2079), .B(n2078), .Z(n2083) );
  NAND U2719 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U2720 ( .A(n2083), .B(n2082), .Z(n2107) );
  AND U2721 ( .A(b[2]), .B(a[14]), .Z(n2113) );
  AND U2722 ( .A(a[15]), .B(b[1]), .Z(n2111) );
  AND U2723 ( .A(a[13]), .B(b[3]), .Z(n2110) );
  XOR U2724 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U2725 ( .A(n2113), .B(n2112), .Z(n2116) );
  NAND U2726 ( .A(b[0]), .B(a[16]), .Z(n2117) );
  XOR U2727 ( .A(n2116), .B(n2117), .Z(n2119) );
  OR U2728 ( .A(n2085), .B(n2084), .Z(n2089) );
  NANDN U2729 ( .A(n2087), .B(n2086), .Z(n2088) );
  NAND U2730 ( .A(n2089), .B(n2088), .Z(n2118) );
  XNOR U2731 ( .A(n2119), .B(n2118), .Z(n2104) );
  NANDN U2732 ( .A(n2091), .B(n2090), .Z(n2095) );
  OR U2733 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2734 ( .A(n2095), .B(n2094), .Z(n2105) );
  XNOR U2735 ( .A(n2104), .B(n2105), .Z(n2106) );
  XOR U2736 ( .A(n2107), .B(n2106), .Z(n2103) );
  NAND U2737 ( .A(n2096), .B(sreg[1035]), .Z(n2100) );
  OR U2738 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U2739 ( .A(n2100), .B(n2099), .Z(n2102) );
  XNOR U2740 ( .A(sreg[1036]), .B(n2102), .Z(n2101) );
  XOR U2741 ( .A(n2103), .B(n2101), .Z(c[1036]) );
  NANDN U2742 ( .A(n2105), .B(n2104), .Z(n2109) );
  NAND U2743 ( .A(n2107), .B(n2106), .Z(n2108) );
  NAND U2744 ( .A(n2109), .B(n2108), .Z(n2125) );
  AND U2745 ( .A(b[2]), .B(a[15]), .Z(n2131) );
  AND U2746 ( .A(a[16]), .B(b[1]), .Z(n2129) );
  AND U2747 ( .A(a[14]), .B(b[3]), .Z(n2128) );
  XOR U2748 ( .A(n2129), .B(n2128), .Z(n2130) );
  XOR U2749 ( .A(n2131), .B(n2130), .Z(n2134) );
  NAND U2750 ( .A(b[0]), .B(a[17]), .Z(n2135) );
  XOR U2751 ( .A(n2134), .B(n2135), .Z(n2137) );
  OR U2752 ( .A(n2111), .B(n2110), .Z(n2115) );
  NANDN U2753 ( .A(n2113), .B(n2112), .Z(n2114) );
  NAND U2754 ( .A(n2115), .B(n2114), .Z(n2136) );
  XNOR U2755 ( .A(n2137), .B(n2136), .Z(n2122) );
  NANDN U2756 ( .A(n2117), .B(n2116), .Z(n2121) );
  OR U2757 ( .A(n2119), .B(n2118), .Z(n2120) );
  NAND U2758 ( .A(n2121), .B(n2120), .Z(n2123) );
  XNOR U2759 ( .A(n2122), .B(n2123), .Z(n2124) );
  XNOR U2760 ( .A(n2125), .B(n2124), .Z(n2140) );
  XNOR U2761 ( .A(n2140), .B(sreg[1037]), .Z(n2141) );
  XOR U2762 ( .A(n2142), .B(n2141), .Z(c[1037]) );
  NANDN U2763 ( .A(n2123), .B(n2122), .Z(n2127) );
  NAND U2764 ( .A(n2125), .B(n2124), .Z(n2126) );
  NAND U2765 ( .A(n2127), .B(n2126), .Z(n2151) );
  AND U2766 ( .A(b[2]), .B(a[16]), .Z(n2157) );
  AND U2767 ( .A(a[17]), .B(b[1]), .Z(n2155) );
  AND U2768 ( .A(a[15]), .B(b[3]), .Z(n2154) );
  XOR U2769 ( .A(n2155), .B(n2154), .Z(n2156) );
  XOR U2770 ( .A(n2157), .B(n2156), .Z(n2160) );
  NAND U2771 ( .A(b[0]), .B(a[18]), .Z(n2161) );
  XOR U2772 ( .A(n2160), .B(n2161), .Z(n2163) );
  OR U2773 ( .A(n2129), .B(n2128), .Z(n2133) );
  NANDN U2774 ( .A(n2131), .B(n2130), .Z(n2132) );
  NAND U2775 ( .A(n2133), .B(n2132), .Z(n2162) );
  XNOR U2776 ( .A(n2163), .B(n2162), .Z(n2148) );
  NANDN U2777 ( .A(n2135), .B(n2134), .Z(n2139) );
  OR U2778 ( .A(n2137), .B(n2136), .Z(n2138) );
  NAND U2779 ( .A(n2139), .B(n2138), .Z(n2149) );
  XNOR U2780 ( .A(n2148), .B(n2149), .Z(n2150) );
  XOR U2781 ( .A(n2151), .B(n2150), .Z(n2147) );
  NAND U2782 ( .A(n2140), .B(sreg[1037]), .Z(n2144) );
  OR U2783 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U2784 ( .A(n2144), .B(n2143), .Z(n2146) );
  XNOR U2785 ( .A(sreg[1038]), .B(n2146), .Z(n2145) );
  XOR U2786 ( .A(n2147), .B(n2145), .Z(c[1038]) );
  NANDN U2787 ( .A(n2149), .B(n2148), .Z(n2153) );
  NAND U2788 ( .A(n2151), .B(n2150), .Z(n2152) );
  NAND U2789 ( .A(n2153), .B(n2152), .Z(n2169) );
  AND U2790 ( .A(b[2]), .B(a[17]), .Z(n2175) );
  AND U2791 ( .A(a[18]), .B(b[1]), .Z(n2173) );
  AND U2792 ( .A(a[16]), .B(b[3]), .Z(n2172) );
  XOR U2793 ( .A(n2173), .B(n2172), .Z(n2174) );
  XOR U2794 ( .A(n2175), .B(n2174), .Z(n2178) );
  NAND U2795 ( .A(b[0]), .B(a[19]), .Z(n2179) );
  XOR U2796 ( .A(n2178), .B(n2179), .Z(n2181) );
  OR U2797 ( .A(n2155), .B(n2154), .Z(n2159) );
  NANDN U2798 ( .A(n2157), .B(n2156), .Z(n2158) );
  NAND U2799 ( .A(n2159), .B(n2158), .Z(n2180) );
  XNOR U2800 ( .A(n2181), .B(n2180), .Z(n2166) );
  NANDN U2801 ( .A(n2161), .B(n2160), .Z(n2165) );
  OR U2802 ( .A(n2163), .B(n2162), .Z(n2164) );
  NAND U2803 ( .A(n2165), .B(n2164), .Z(n2167) );
  XNOR U2804 ( .A(n2166), .B(n2167), .Z(n2168) );
  XOR U2805 ( .A(n2169), .B(n2168), .Z(n2184) );
  XNOR U2806 ( .A(sreg[1039]), .B(n2184), .Z(n2185) );
  XNOR U2807 ( .A(n2186), .B(n2185), .Z(c[1039]) );
  NANDN U2808 ( .A(n2167), .B(n2166), .Z(n2171) );
  NAND U2809 ( .A(n2169), .B(n2168), .Z(n2170) );
  NAND U2810 ( .A(n2171), .B(n2170), .Z(n2195) );
  AND U2811 ( .A(b[2]), .B(a[18]), .Z(n2201) );
  AND U2812 ( .A(a[19]), .B(b[1]), .Z(n2199) );
  AND U2813 ( .A(a[17]), .B(b[3]), .Z(n2198) );
  XOR U2814 ( .A(n2199), .B(n2198), .Z(n2200) );
  XOR U2815 ( .A(n2201), .B(n2200), .Z(n2204) );
  NAND U2816 ( .A(b[0]), .B(a[20]), .Z(n2205) );
  XOR U2817 ( .A(n2204), .B(n2205), .Z(n2207) );
  OR U2818 ( .A(n2173), .B(n2172), .Z(n2177) );
  NANDN U2819 ( .A(n2175), .B(n2174), .Z(n2176) );
  NAND U2820 ( .A(n2177), .B(n2176), .Z(n2206) );
  XNOR U2821 ( .A(n2207), .B(n2206), .Z(n2192) );
  NANDN U2822 ( .A(n2179), .B(n2178), .Z(n2183) );
  OR U2823 ( .A(n2181), .B(n2180), .Z(n2182) );
  NAND U2824 ( .A(n2183), .B(n2182), .Z(n2193) );
  XNOR U2825 ( .A(n2192), .B(n2193), .Z(n2194) );
  XOR U2826 ( .A(n2195), .B(n2194), .Z(n2191) );
  NANDN U2827 ( .A(sreg[1039]), .B(n2184), .Z(n2188) );
  NAND U2828 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2829 ( .A(n2188), .B(n2187), .Z(n2190) );
  XNOR U2830 ( .A(sreg[1040]), .B(n2190), .Z(n2189) );
  XOR U2831 ( .A(n2191), .B(n2189), .Z(c[1040]) );
  NANDN U2832 ( .A(n2193), .B(n2192), .Z(n2197) );
  NAND U2833 ( .A(n2195), .B(n2194), .Z(n2196) );
  NAND U2834 ( .A(n2197), .B(n2196), .Z(n2213) );
  AND U2835 ( .A(b[2]), .B(a[19]), .Z(n2219) );
  AND U2836 ( .A(a[20]), .B(b[1]), .Z(n2217) );
  AND U2837 ( .A(a[18]), .B(b[3]), .Z(n2216) );
  XOR U2838 ( .A(n2217), .B(n2216), .Z(n2218) );
  XOR U2839 ( .A(n2219), .B(n2218), .Z(n2222) );
  NAND U2840 ( .A(b[0]), .B(a[21]), .Z(n2223) );
  XOR U2841 ( .A(n2222), .B(n2223), .Z(n2225) );
  OR U2842 ( .A(n2199), .B(n2198), .Z(n2203) );
  NANDN U2843 ( .A(n2201), .B(n2200), .Z(n2202) );
  NAND U2844 ( .A(n2203), .B(n2202), .Z(n2224) );
  XNOR U2845 ( .A(n2225), .B(n2224), .Z(n2210) );
  NANDN U2846 ( .A(n2205), .B(n2204), .Z(n2209) );
  OR U2847 ( .A(n2207), .B(n2206), .Z(n2208) );
  NAND U2848 ( .A(n2209), .B(n2208), .Z(n2211) );
  XNOR U2849 ( .A(n2210), .B(n2211), .Z(n2212) );
  XNOR U2850 ( .A(n2213), .B(n2212), .Z(n2228) );
  XOR U2851 ( .A(sreg[1041]), .B(n2228), .Z(n2230) );
  XNOR U2852 ( .A(n2229), .B(n2230), .Z(c[1041]) );
  NANDN U2853 ( .A(n2211), .B(n2210), .Z(n2215) );
  NAND U2854 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U2855 ( .A(n2215), .B(n2214), .Z(n2236) );
  AND U2856 ( .A(b[2]), .B(a[20]), .Z(n2242) );
  AND U2857 ( .A(a[21]), .B(b[1]), .Z(n2240) );
  AND U2858 ( .A(a[19]), .B(b[3]), .Z(n2239) );
  XOR U2859 ( .A(n2240), .B(n2239), .Z(n2241) );
  XOR U2860 ( .A(n2242), .B(n2241), .Z(n2245) );
  NAND U2861 ( .A(b[0]), .B(a[22]), .Z(n2246) );
  XOR U2862 ( .A(n2245), .B(n2246), .Z(n2248) );
  OR U2863 ( .A(n2217), .B(n2216), .Z(n2221) );
  NANDN U2864 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2865 ( .A(n2221), .B(n2220), .Z(n2247) );
  XNOR U2866 ( .A(n2248), .B(n2247), .Z(n2233) );
  NANDN U2867 ( .A(n2223), .B(n2222), .Z(n2227) );
  OR U2868 ( .A(n2225), .B(n2224), .Z(n2226) );
  NAND U2869 ( .A(n2227), .B(n2226), .Z(n2234) );
  XNOR U2870 ( .A(n2233), .B(n2234), .Z(n2235) );
  XNOR U2871 ( .A(n2236), .B(n2235), .Z(n2251) );
  XOR U2872 ( .A(sreg[1042]), .B(n2251), .Z(n2252) );
  OR U2873 ( .A(n2228), .B(sreg[1041]), .Z(n2232) );
  NAND U2874 ( .A(n2230), .B(n2229), .Z(n2231) );
  AND U2875 ( .A(n2232), .B(n2231), .Z(n2253) );
  XOR U2876 ( .A(n2252), .B(n2253), .Z(c[1042]) );
  NANDN U2877 ( .A(n2234), .B(n2233), .Z(n2238) );
  NAND U2878 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2879 ( .A(n2238), .B(n2237), .Z(n2262) );
  AND U2880 ( .A(b[2]), .B(a[21]), .Z(n2268) );
  AND U2881 ( .A(a[22]), .B(b[1]), .Z(n2266) );
  AND U2882 ( .A(a[20]), .B(b[3]), .Z(n2265) );
  XOR U2883 ( .A(n2266), .B(n2265), .Z(n2267) );
  XOR U2884 ( .A(n2268), .B(n2267), .Z(n2271) );
  NAND U2885 ( .A(b[0]), .B(a[23]), .Z(n2272) );
  XOR U2886 ( .A(n2271), .B(n2272), .Z(n2274) );
  OR U2887 ( .A(n2240), .B(n2239), .Z(n2244) );
  NANDN U2888 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U2889 ( .A(n2244), .B(n2243), .Z(n2273) );
  XNOR U2890 ( .A(n2274), .B(n2273), .Z(n2259) );
  NANDN U2891 ( .A(n2246), .B(n2245), .Z(n2250) );
  OR U2892 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U2893 ( .A(n2250), .B(n2249), .Z(n2260) );
  XNOR U2894 ( .A(n2259), .B(n2260), .Z(n2261) );
  XOR U2895 ( .A(n2262), .B(n2261), .Z(n2258) );
  OR U2896 ( .A(n2251), .B(sreg[1042]), .Z(n2255) );
  NANDN U2897 ( .A(n2253), .B(n2252), .Z(n2254) );
  AND U2898 ( .A(n2255), .B(n2254), .Z(n2257) );
  XNOR U2899 ( .A(sreg[1043]), .B(n2257), .Z(n2256) );
  XOR U2900 ( .A(n2258), .B(n2256), .Z(c[1043]) );
  NANDN U2901 ( .A(n2260), .B(n2259), .Z(n2264) );
  NAND U2902 ( .A(n2262), .B(n2261), .Z(n2263) );
  NAND U2903 ( .A(n2264), .B(n2263), .Z(n2280) );
  AND U2904 ( .A(b[2]), .B(a[22]), .Z(n2286) );
  AND U2905 ( .A(a[23]), .B(b[1]), .Z(n2284) );
  AND U2906 ( .A(a[21]), .B(b[3]), .Z(n2283) );
  XOR U2907 ( .A(n2284), .B(n2283), .Z(n2285) );
  XOR U2908 ( .A(n2286), .B(n2285), .Z(n2289) );
  NAND U2909 ( .A(b[0]), .B(a[24]), .Z(n2290) );
  XOR U2910 ( .A(n2289), .B(n2290), .Z(n2292) );
  OR U2911 ( .A(n2266), .B(n2265), .Z(n2270) );
  NANDN U2912 ( .A(n2268), .B(n2267), .Z(n2269) );
  NAND U2913 ( .A(n2270), .B(n2269), .Z(n2291) );
  XNOR U2914 ( .A(n2292), .B(n2291), .Z(n2277) );
  NANDN U2915 ( .A(n2272), .B(n2271), .Z(n2276) );
  OR U2916 ( .A(n2274), .B(n2273), .Z(n2275) );
  NAND U2917 ( .A(n2276), .B(n2275), .Z(n2278) );
  XNOR U2918 ( .A(n2277), .B(n2278), .Z(n2279) );
  XNOR U2919 ( .A(n2280), .B(n2279), .Z(n2295) );
  XOR U2920 ( .A(sreg[1044]), .B(n2295), .Z(n2297) );
  XNOR U2921 ( .A(n2296), .B(n2297), .Z(c[1044]) );
  NANDN U2922 ( .A(n2278), .B(n2277), .Z(n2282) );
  NAND U2923 ( .A(n2280), .B(n2279), .Z(n2281) );
  NAND U2924 ( .A(n2282), .B(n2281), .Z(n2306) );
  AND U2925 ( .A(b[2]), .B(a[23]), .Z(n2312) );
  AND U2926 ( .A(a[24]), .B(b[1]), .Z(n2310) );
  AND U2927 ( .A(a[22]), .B(b[3]), .Z(n2309) );
  XOR U2928 ( .A(n2310), .B(n2309), .Z(n2311) );
  XOR U2929 ( .A(n2312), .B(n2311), .Z(n2315) );
  NAND U2930 ( .A(b[0]), .B(a[25]), .Z(n2316) );
  XOR U2931 ( .A(n2315), .B(n2316), .Z(n2318) );
  OR U2932 ( .A(n2284), .B(n2283), .Z(n2288) );
  NANDN U2933 ( .A(n2286), .B(n2285), .Z(n2287) );
  NAND U2934 ( .A(n2288), .B(n2287), .Z(n2317) );
  XNOR U2935 ( .A(n2318), .B(n2317), .Z(n2303) );
  NANDN U2936 ( .A(n2290), .B(n2289), .Z(n2294) );
  OR U2937 ( .A(n2292), .B(n2291), .Z(n2293) );
  NAND U2938 ( .A(n2294), .B(n2293), .Z(n2304) );
  XNOR U2939 ( .A(n2303), .B(n2304), .Z(n2305) );
  XOR U2940 ( .A(n2306), .B(n2305), .Z(n2302) );
  OR U2941 ( .A(n2295), .B(sreg[1044]), .Z(n2299) );
  NAND U2942 ( .A(n2297), .B(n2296), .Z(n2298) );
  AND U2943 ( .A(n2299), .B(n2298), .Z(n2301) );
  XNOR U2944 ( .A(sreg[1045]), .B(n2301), .Z(n2300) );
  XOR U2945 ( .A(n2302), .B(n2300), .Z(c[1045]) );
  NANDN U2946 ( .A(n2304), .B(n2303), .Z(n2308) );
  NAND U2947 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U2948 ( .A(n2308), .B(n2307), .Z(n2324) );
  AND U2949 ( .A(b[2]), .B(a[24]), .Z(n2330) );
  AND U2950 ( .A(a[25]), .B(b[1]), .Z(n2328) );
  AND U2951 ( .A(a[23]), .B(b[3]), .Z(n2327) );
  XOR U2952 ( .A(n2328), .B(n2327), .Z(n2329) );
  XOR U2953 ( .A(n2330), .B(n2329), .Z(n2333) );
  NAND U2954 ( .A(b[0]), .B(a[26]), .Z(n2334) );
  XOR U2955 ( .A(n2333), .B(n2334), .Z(n2336) );
  OR U2956 ( .A(n2310), .B(n2309), .Z(n2314) );
  NANDN U2957 ( .A(n2312), .B(n2311), .Z(n2313) );
  NAND U2958 ( .A(n2314), .B(n2313), .Z(n2335) );
  XNOR U2959 ( .A(n2336), .B(n2335), .Z(n2321) );
  NANDN U2960 ( .A(n2316), .B(n2315), .Z(n2320) );
  OR U2961 ( .A(n2318), .B(n2317), .Z(n2319) );
  NAND U2962 ( .A(n2320), .B(n2319), .Z(n2322) );
  XNOR U2963 ( .A(n2321), .B(n2322), .Z(n2323) );
  XNOR U2964 ( .A(n2324), .B(n2323), .Z(n2339) );
  XNOR U2965 ( .A(n2339), .B(sreg[1046]), .Z(n2340) );
  XOR U2966 ( .A(n2341), .B(n2340), .Z(c[1046]) );
  NANDN U2967 ( .A(n2322), .B(n2321), .Z(n2326) );
  NAND U2968 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U2969 ( .A(n2326), .B(n2325), .Z(n2348) );
  AND U2970 ( .A(b[2]), .B(a[25]), .Z(n2354) );
  AND U2971 ( .A(a[26]), .B(b[1]), .Z(n2352) );
  AND U2972 ( .A(a[24]), .B(b[3]), .Z(n2351) );
  XOR U2973 ( .A(n2352), .B(n2351), .Z(n2353) );
  XOR U2974 ( .A(n2354), .B(n2353), .Z(n2357) );
  NAND U2975 ( .A(b[0]), .B(a[27]), .Z(n2358) );
  XOR U2976 ( .A(n2357), .B(n2358), .Z(n2360) );
  OR U2977 ( .A(n2328), .B(n2327), .Z(n2332) );
  NANDN U2978 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U2979 ( .A(n2332), .B(n2331), .Z(n2359) );
  XNOR U2980 ( .A(n2360), .B(n2359), .Z(n2345) );
  NANDN U2981 ( .A(n2334), .B(n2333), .Z(n2338) );
  OR U2982 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U2983 ( .A(n2338), .B(n2337), .Z(n2346) );
  XNOR U2984 ( .A(n2345), .B(n2346), .Z(n2347) );
  XOR U2985 ( .A(n2348), .B(n2347), .Z(n2364) );
  NAND U2986 ( .A(n2339), .B(sreg[1046]), .Z(n2343) );
  OR U2987 ( .A(n2341), .B(n2340), .Z(n2342) );
  NAND U2988 ( .A(n2343), .B(n2342), .Z(n2363) );
  XNOR U2989 ( .A(sreg[1047]), .B(n2363), .Z(n2344) );
  XOR U2990 ( .A(n2364), .B(n2344), .Z(c[1047]) );
  NANDN U2991 ( .A(n2346), .B(n2345), .Z(n2350) );
  NAND U2992 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U2993 ( .A(n2350), .B(n2349), .Z(n2369) );
  AND U2994 ( .A(b[2]), .B(a[26]), .Z(n2375) );
  AND U2995 ( .A(a[27]), .B(b[1]), .Z(n2373) );
  AND U2996 ( .A(a[25]), .B(b[3]), .Z(n2372) );
  XOR U2997 ( .A(n2373), .B(n2372), .Z(n2374) );
  XOR U2998 ( .A(n2375), .B(n2374), .Z(n2378) );
  NAND U2999 ( .A(b[0]), .B(a[28]), .Z(n2379) );
  XOR U3000 ( .A(n2378), .B(n2379), .Z(n2381) );
  OR U3001 ( .A(n2352), .B(n2351), .Z(n2356) );
  NANDN U3002 ( .A(n2354), .B(n2353), .Z(n2355) );
  NAND U3003 ( .A(n2356), .B(n2355), .Z(n2380) );
  XNOR U3004 ( .A(n2381), .B(n2380), .Z(n2366) );
  NANDN U3005 ( .A(n2358), .B(n2357), .Z(n2362) );
  OR U3006 ( .A(n2360), .B(n2359), .Z(n2361) );
  NAND U3007 ( .A(n2362), .B(n2361), .Z(n2367) );
  XNOR U3008 ( .A(n2366), .B(n2367), .Z(n2368) );
  XOR U3009 ( .A(n2369), .B(n2368), .Z(n2385) );
  XNOR U3010 ( .A(sreg[1048]), .B(n2384), .Z(n2365) );
  XOR U3011 ( .A(n2385), .B(n2365), .Z(c[1048]) );
  NANDN U3012 ( .A(n2367), .B(n2366), .Z(n2371) );
  NAND U3013 ( .A(n2369), .B(n2368), .Z(n2370) );
  NAND U3014 ( .A(n2371), .B(n2370), .Z(n2392) );
  AND U3015 ( .A(b[2]), .B(a[27]), .Z(n2398) );
  AND U3016 ( .A(a[28]), .B(b[1]), .Z(n2396) );
  AND U3017 ( .A(a[26]), .B(b[3]), .Z(n2395) );
  XOR U3018 ( .A(n2396), .B(n2395), .Z(n2397) );
  XOR U3019 ( .A(n2398), .B(n2397), .Z(n2401) );
  NAND U3020 ( .A(b[0]), .B(a[29]), .Z(n2402) );
  XOR U3021 ( .A(n2401), .B(n2402), .Z(n2404) );
  OR U3022 ( .A(n2373), .B(n2372), .Z(n2377) );
  NANDN U3023 ( .A(n2375), .B(n2374), .Z(n2376) );
  NAND U3024 ( .A(n2377), .B(n2376), .Z(n2403) );
  XNOR U3025 ( .A(n2404), .B(n2403), .Z(n2389) );
  NANDN U3026 ( .A(n2379), .B(n2378), .Z(n2383) );
  OR U3027 ( .A(n2381), .B(n2380), .Z(n2382) );
  NAND U3028 ( .A(n2383), .B(n2382), .Z(n2390) );
  XNOR U3029 ( .A(n2389), .B(n2390), .Z(n2391) );
  XOR U3030 ( .A(n2392), .B(n2391), .Z(n2388) );
  XNOR U3031 ( .A(sreg[1049]), .B(n2387), .Z(n2386) );
  XOR U3032 ( .A(n2388), .B(n2386), .Z(c[1049]) );
  NANDN U3033 ( .A(n2390), .B(n2389), .Z(n2394) );
  NAND U3034 ( .A(n2392), .B(n2391), .Z(n2393) );
  NAND U3035 ( .A(n2394), .B(n2393), .Z(n2410) );
  AND U3036 ( .A(b[2]), .B(a[28]), .Z(n2416) );
  AND U3037 ( .A(a[29]), .B(b[1]), .Z(n2414) );
  AND U3038 ( .A(a[27]), .B(b[3]), .Z(n2413) );
  XOR U3039 ( .A(n2414), .B(n2413), .Z(n2415) );
  XOR U3040 ( .A(n2416), .B(n2415), .Z(n2419) );
  NAND U3041 ( .A(b[0]), .B(a[30]), .Z(n2420) );
  XOR U3042 ( .A(n2419), .B(n2420), .Z(n2422) );
  OR U3043 ( .A(n2396), .B(n2395), .Z(n2400) );
  NANDN U3044 ( .A(n2398), .B(n2397), .Z(n2399) );
  NAND U3045 ( .A(n2400), .B(n2399), .Z(n2421) );
  XNOR U3046 ( .A(n2422), .B(n2421), .Z(n2407) );
  NANDN U3047 ( .A(n2402), .B(n2401), .Z(n2406) );
  OR U3048 ( .A(n2404), .B(n2403), .Z(n2405) );
  NAND U3049 ( .A(n2406), .B(n2405), .Z(n2408) );
  XNOR U3050 ( .A(n2407), .B(n2408), .Z(n2409) );
  XNOR U3051 ( .A(n2410), .B(n2409), .Z(n2425) );
  XOR U3052 ( .A(sreg[1050]), .B(n2425), .Z(n2427) );
  XNOR U3053 ( .A(n2426), .B(n2427), .Z(c[1050]) );
  NANDN U3054 ( .A(n2408), .B(n2407), .Z(n2412) );
  NAND U3055 ( .A(n2410), .B(n2409), .Z(n2411) );
  NAND U3056 ( .A(n2412), .B(n2411), .Z(n2436) );
  AND U3057 ( .A(b[2]), .B(a[29]), .Z(n2442) );
  AND U3058 ( .A(a[30]), .B(b[1]), .Z(n2440) );
  AND U3059 ( .A(a[28]), .B(b[3]), .Z(n2439) );
  XOR U3060 ( .A(n2440), .B(n2439), .Z(n2441) );
  XOR U3061 ( .A(n2442), .B(n2441), .Z(n2445) );
  NAND U3062 ( .A(b[0]), .B(a[31]), .Z(n2446) );
  XOR U3063 ( .A(n2445), .B(n2446), .Z(n2448) );
  OR U3064 ( .A(n2414), .B(n2413), .Z(n2418) );
  NANDN U3065 ( .A(n2416), .B(n2415), .Z(n2417) );
  NAND U3066 ( .A(n2418), .B(n2417), .Z(n2447) );
  XNOR U3067 ( .A(n2448), .B(n2447), .Z(n2433) );
  NANDN U3068 ( .A(n2420), .B(n2419), .Z(n2424) );
  OR U3069 ( .A(n2422), .B(n2421), .Z(n2423) );
  NAND U3070 ( .A(n2424), .B(n2423), .Z(n2434) );
  XNOR U3071 ( .A(n2433), .B(n2434), .Z(n2435) );
  XOR U3072 ( .A(n2436), .B(n2435), .Z(n2432) );
  OR U3073 ( .A(n2425), .B(sreg[1050]), .Z(n2429) );
  NAND U3074 ( .A(n2427), .B(n2426), .Z(n2428) );
  AND U3075 ( .A(n2429), .B(n2428), .Z(n2431) );
  XNOR U3076 ( .A(sreg[1051]), .B(n2431), .Z(n2430) );
  XOR U3077 ( .A(n2432), .B(n2430), .Z(c[1051]) );
  NANDN U3078 ( .A(n2434), .B(n2433), .Z(n2438) );
  NAND U3079 ( .A(n2436), .B(n2435), .Z(n2437) );
  NAND U3080 ( .A(n2438), .B(n2437), .Z(n2454) );
  AND U3081 ( .A(b[2]), .B(a[30]), .Z(n2466) );
  AND U3082 ( .A(a[31]), .B(b[1]), .Z(n2464) );
  AND U3083 ( .A(a[29]), .B(b[3]), .Z(n2463) );
  XOR U3084 ( .A(n2464), .B(n2463), .Z(n2465) );
  XOR U3085 ( .A(n2466), .B(n2465), .Z(n2457) );
  NAND U3086 ( .A(b[0]), .B(a[32]), .Z(n2458) );
  XOR U3087 ( .A(n2457), .B(n2458), .Z(n2460) );
  OR U3088 ( .A(n2440), .B(n2439), .Z(n2444) );
  NANDN U3089 ( .A(n2442), .B(n2441), .Z(n2443) );
  NAND U3090 ( .A(n2444), .B(n2443), .Z(n2459) );
  XNOR U3091 ( .A(n2460), .B(n2459), .Z(n2451) );
  NANDN U3092 ( .A(n2446), .B(n2445), .Z(n2450) );
  OR U3093 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U3094 ( .A(n2450), .B(n2449), .Z(n2452) );
  XNOR U3095 ( .A(n2451), .B(n2452), .Z(n2453) );
  XNOR U3096 ( .A(n2454), .B(n2453), .Z(n2470) );
  XOR U3097 ( .A(sreg[1052]), .B(n2470), .Z(n2472) );
  XNOR U3098 ( .A(n2471), .B(n2472), .Z(c[1052]) );
  NANDN U3099 ( .A(n2452), .B(n2451), .Z(n2456) );
  NAND U3100 ( .A(n2454), .B(n2453), .Z(n2455) );
  AND U3101 ( .A(n2456), .B(n2455), .Z(n2478) );
  NANDN U3102 ( .A(n2458), .B(n2457), .Z(n2462) );
  OR U3103 ( .A(n2460), .B(n2459), .Z(n2461) );
  AND U3104 ( .A(n2462), .B(n2461), .Z(n2477) );
  AND U3105 ( .A(b[2]), .B(a[31]), .Z(n2482) );
  AND U3106 ( .A(a[32]), .B(b[1]), .Z(n2480) );
  AND U3107 ( .A(a[30]), .B(b[3]), .Z(n2479) );
  XOR U3108 ( .A(n2480), .B(n2479), .Z(n2481) );
  XOR U3109 ( .A(n2482), .B(n2481), .Z(n2485) );
  NAND U3110 ( .A(b[0]), .B(a[33]), .Z(n2486) );
  XOR U3111 ( .A(n2485), .B(n2486), .Z(n2488) );
  OR U3112 ( .A(n2464), .B(n2463), .Z(n2468) );
  NANDN U3113 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U3114 ( .A(n2468), .B(n2467), .Z(n2487) );
  XOR U3115 ( .A(n2488), .B(n2487), .Z(n2476) );
  XNOR U3116 ( .A(n2477), .B(n2476), .Z(n2469) );
  XOR U3117 ( .A(n2478), .B(n2469), .Z(n2492) );
  OR U3118 ( .A(n2470), .B(sreg[1052]), .Z(n2474) );
  NAND U3119 ( .A(n2472), .B(n2471), .Z(n2473) );
  AND U3120 ( .A(n2474), .B(n2473), .Z(n2491) );
  XNOR U3121 ( .A(sreg[1053]), .B(n2491), .Z(n2475) );
  XNOR U3122 ( .A(n2492), .B(n2475), .Z(c[1053]) );
  AND U3123 ( .A(b[2]), .B(a[32]), .Z(n2503) );
  AND U3124 ( .A(a[33]), .B(b[1]), .Z(n2501) );
  AND U3125 ( .A(a[31]), .B(b[3]), .Z(n2500) );
  XOR U3126 ( .A(n2501), .B(n2500), .Z(n2502) );
  XOR U3127 ( .A(n2503), .B(n2502), .Z(n2506) );
  NAND U3128 ( .A(b[0]), .B(a[34]), .Z(n2507) );
  XOR U3129 ( .A(n2506), .B(n2507), .Z(n2509) );
  OR U3130 ( .A(n2480), .B(n2479), .Z(n2484) );
  NANDN U3131 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U3132 ( .A(n2484), .B(n2483), .Z(n2508) );
  XNOR U3133 ( .A(n2509), .B(n2508), .Z(n2494) );
  NANDN U3134 ( .A(n2486), .B(n2485), .Z(n2490) );
  OR U3135 ( .A(n2488), .B(n2487), .Z(n2489) );
  NAND U3136 ( .A(n2490), .B(n2489), .Z(n2495) );
  XNOR U3137 ( .A(n2494), .B(n2495), .Z(n2496) );
  XOR U3138 ( .A(n2497), .B(n2496), .Z(n2513) );
  XNOR U3139 ( .A(sreg[1054]), .B(n2512), .Z(n2493) );
  XNOR U3140 ( .A(n2513), .B(n2493), .Z(c[1054]) );
  NANDN U3141 ( .A(n2495), .B(n2494), .Z(n2499) );
  NANDN U3142 ( .A(n2497), .B(n2496), .Z(n2498) );
  NAND U3143 ( .A(n2499), .B(n2498), .Z(n2518) );
  AND U3144 ( .A(b[2]), .B(a[33]), .Z(n2524) );
  AND U3145 ( .A(a[34]), .B(b[1]), .Z(n2522) );
  AND U3146 ( .A(a[32]), .B(b[3]), .Z(n2521) );
  XOR U3147 ( .A(n2522), .B(n2521), .Z(n2523) );
  XOR U3148 ( .A(n2524), .B(n2523), .Z(n2527) );
  NAND U3149 ( .A(b[0]), .B(a[35]), .Z(n2528) );
  XOR U3150 ( .A(n2527), .B(n2528), .Z(n2530) );
  OR U3151 ( .A(n2501), .B(n2500), .Z(n2505) );
  NANDN U3152 ( .A(n2503), .B(n2502), .Z(n2504) );
  NAND U3153 ( .A(n2505), .B(n2504), .Z(n2529) );
  XNOR U3154 ( .A(n2530), .B(n2529), .Z(n2515) );
  NANDN U3155 ( .A(n2507), .B(n2506), .Z(n2511) );
  OR U3156 ( .A(n2509), .B(n2508), .Z(n2510) );
  NAND U3157 ( .A(n2511), .B(n2510), .Z(n2516) );
  XNOR U3158 ( .A(n2515), .B(n2516), .Z(n2517) );
  XNOR U3159 ( .A(n2518), .B(n2517), .Z(n2534) );
  XOR U3160 ( .A(sreg[1055]), .B(n2535), .Z(n2514) );
  XNOR U3161 ( .A(n2534), .B(n2514), .Z(c[1055]) );
  NANDN U3162 ( .A(n2516), .B(n2515), .Z(n2520) );
  NAND U3163 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U3164 ( .A(n2520), .B(n2519), .Z(n2541) );
  AND U3165 ( .A(b[2]), .B(a[34]), .Z(n2549) );
  AND U3166 ( .A(a[35]), .B(b[1]), .Z(n2547) );
  AND U3167 ( .A(a[33]), .B(b[3]), .Z(n2546) );
  XOR U3168 ( .A(n2547), .B(n2546), .Z(n2548) );
  XOR U3169 ( .A(n2549), .B(n2548), .Z(n2542) );
  NAND U3170 ( .A(b[0]), .B(a[36]), .Z(n2543) );
  XOR U3171 ( .A(n2542), .B(n2543), .Z(n2544) );
  OR U3172 ( .A(n2522), .B(n2521), .Z(n2526) );
  NANDN U3173 ( .A(n2524), .B(n2523), .Z(n2525) );
  AND U3174 ( .A(n2526), .B(n2525), .Z(n2545) );
  XOR U3175 ( .A(n2544), .B(n2545), .Z(n2539) );
  NANDN U3176 ( .A(n2528), .B(n2527), .Z(n2532) );
  OR U3177 ( .A(n2530), .B(n2529), .Z(n2531) );
  AND U3178 ( .A(n2532), .B(n2531), .Z(n2540) );
  XOR U3179 ( .A(n2539), .B(n2540), .Z(n2533) );
  XOR U3180 ( .A(n2541), .B(n2533), .Z(n2538) );
  XOR U3181 ( .A(n2537), .B(sreg[1056]), .Z(n2536) );
  XNOR U3182 ( .A(n2538), .B(n2536), .Z(c[1056]) );
  AND U3183 ( .A(b[2]), .B(a[35]), .Z(n2555) );
  AND U3184 ( .A(a[36]), .B(b[1]), .Z(n2553) );
  AND U3185 ( .A(a[34]), .B(b[3]), .Z(n2552) );
  XOR U3186 ( .A(n2553), .B(n2552), .Z(n2554) );
  XOR U3187 ( .A(n2555), .B(n2554), .Z(n2558) );
  NAND U3188 ( .A(b[0]), .B(a[37]), .Z(n2559) );
  XNOR U3189 ( .A(n2558), .B(n2559), .Z(n2560) );
  OR U3190 ( .A(n2547), .B(n2546), .Z(n2551) );
  NANDN U3191 ( .A(n2549), .B(n2548), .Z(n2550) );
  AND U3192 ( .A(n2551), .B(n2550), .Z(n2561) );
  XNOR U3193 ( .A(n2560), .B(n2561), .Z(n2565) );
  XNOR U3194 ( .A(n2564), .B(n2565), .Z(n2566) );
  XNOR U3195 ( .A(n2567), .B(n2566), .Z(n2570) );
  XNOR U3196 ( .A(sreg[1057]), .B(n2570), .Z(n2572) );
  XNOR U3197 ( .A(n2571), .B(n2572), .Z(c[1057]) );
  AND U3198 ( .A(b[2]), .B(a[36]), .Z(n2587) );
  AND U3199 ( .A(a[37]), .B(b[1]), .Z(n2585) );
  AND U3200 ( .A(a[35]), .B(b[3]), .Z(n2584) );
  XOR U3201 ( .A(n2585), .B(n2584), .Z(n2586) );
  XOR U3202 ( .A(n2587), .B(n2586), .Z(n2590) );
  NAND U3203 ( .A(b[0]), .B(a[38]), .Z(n2591) );
  XOR U3204 ( .A(n2590), .B(n2591), .Z(n2593) );
  OR U3205 ( .A(n2553), .B(n2552), .Z(n2557) );
  NANDN U3206 ( .A(n2555), .B(n2554), .Z(n2556) );
  NAND U3207 ( .A(n2557), .B(n2556), .Z(n2592) );
  XNOR U3208 ( .A(n2593), .B(n2592), .Z(n2578) );
  NANDN U3209 ( .A(n2559), .B(n2558), .Z(n2563) );
  NAND U3210 ( .A(n2561), .B(n2560), .Z(n2562) );
  NAND U3211 ( .A(n2563), .B(n2562), .Z(n2579) );
  XNOR U3212 ( .A(n2578), .B(n2579), .Z(n2580) );
  NANDN U3213 ( .A(n2565), .B(n2564), .Z(n2569) );
  NANDN U3214 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U3215 ( .A(n2569), .B(n2568), .Z(n2581) );
  XNOR U3216 ( .A(n2580), .B(n2581), .Z(n2577) );
  NAND U3217 ( .A(sreg[1057]), .B(n2570), .Z(n2574) );
  NANDN U3218 ( .A(n2572), .B(n2571), .Z(n2573) );
  AND U3219 ( .A(n2574), .B(n2573), .Z(n2576) );
  XNOR U3220 ( .A(n2576), .B(sreg[1058]), .Z(n2575) );
  XOR U3221 ( .A(n2577), .B(n2575), .Z(c[1058]) );
  NANDN U3222 ( .A(n2579), .B(n2578), .Z(n2583) );
  NAND U3223 ( .A(n2581), .B(n2580), .Z(n2582) );
  NAND U3224 ( .A(n2583), .B(n2582), .Z(n2616) );
  AND U3225 ( .A(b[2]), .B(a[37]), .Z(n2610) );
  AND U3226 ( .A(a[38]), .B(b[1]), .Z(n2608) );
  AND U3227 ( .A(a[36]), .B(b[3]), .Z(n2607) );
  XOR U3228 ( .A(n2608), .B(n2607), .Z(n2609) );
  XOR U3229 ( .A(n2610), .B(n2609), .Z(n2601) );
  NAND U3230 ( .A(b[0]), .B(a[39]), .Z(n2602) );
  XOR U3231 ( .A(n2601), .B(n2602), .Z(n2604) );
  OR U3232 ( .A(n2585), .B(n2584), .Z(n2589) );
  NANDN U3233 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U3234 ( .A(n2589), .B(n2588), .Z(n2603) );
  XNOR U3235 ( .A(n2604), .B(n2603), .Z(n2613) );
  NANDN U3236 ( .A(n2591), .B(n2590), .Z(n2595) );
  OR U3237 ( .A(n2593), .B(n2592), .Z(n2594) );
  NAND U3238 ( .A(n2595), .B(n2594), .Z(n2614) );
  XNOR U3239 ( .A(n2613), .B(n2614), .Z(n2615) );
  XNOR U3240 ( .A(n2616), .B(n2615), .Z(n2596) );
  XNOR U3241 ( .A(n2596), .B(sreg[1059]), .Z(n2598) );
  XNOR U3242 ( .A(n2597), .B(n2598), .Z(c[1059]) );
  NAND U3243 ( .A(n2596), .B(sreg[1059]), .Z(n2600) );
  NANDN U3244 ( .A(n2598), .B(n2597), .Z(n2599) );
  NAND U3245 ( .A(n2600), .B(n2599), .Z(n2620) );
  NANDN U3246 ( .A(n2602), .B(n2601), .Z(n2606) );
  OR U3247 ( .A(n2604), .B(n2603), .Z(n2605) );
  NAND U3248 ( .A(n2606), .B(n2605), .Z(n2634) );
  AND U3249 ( .A(b[2]), .B(a[38]), .Z(n2625) );
  AND U3250 ( .A(a[39]), .B(b[1]), .Z(n2623) );
  AND U3251 ( .A(a[37]), .B(b[3]), .Z(n2622) );
  XOR U3252 ( .A(n2623), .B(n2622), .Z(n2624) );
  XOR U3253 ( .A(n2625), .B(n2624), .Z(n2628) );
  NAND U3254 ( .A(b[0]), .B(a[40]), .Z(n2629) );
  XNOR U3255 ( .A(n2628), .B(n2629), .Z(n2630) );
  OR U3256 ( .A(n2608), .B(n2607), .Z(n2612) );
  NANDN U3257 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U3258 ( .A(n2612), .B(n2611), .Z(n2631) );
  XNOR U3259 ( .A(n2630), .B(n2631), .Z(n2635) );
  XNOR U3260 ( .A(n2634), .B(n2635), .Z(n2636) );
  NANDN U3261 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U3262 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U3263 ( .A(n2618), .B(n2617), .Z(n2637) );
  XNOR U3264 ( .A(n2636), .B(n2637), .Z(n2621) );
  XOR U3265 ( .A(sreg[1060]), .B(n2621), .Z(n2619) );
  XNOR U3266 ( .A(n2620), .B(n2619), .Z(c[1060]) );
  AND U3267 ( .A(b[2]), .B(a[39]), .Z(n2649) );
  AND U3268 ( .A(a[40]), .B(b[1]), .Z(n2647) );
  AND U3269 ( .A(a[38]), .B(b[3]), .Z(n2646) );
  XOR U3270 ( .A(n2647), .B(n2646), .Z(n2648) );
  XOR U3271 ( .A(n2649), .B(n2648), .Z(n2652) );
  NAND U3272 ( .A(b[0]), .B(a[41]), .Z(n2653) );
  XOR U3273 ( .A(n2652), .B(n2653), .Z(n2655) );
  OR U3274 ( .A(n2623), .B(n2622), .Z(n2627) );
  NANDN U3275 ( .A(n2625), .B(n2624), .Z(n2626) );
  NAND U3276 ( .A(n2627), .B(n2626), .Z(n2654) );
  XNOR U3277 ( .A(n2655), .B(n2654), .Z(n2640) );
  NANDN U3278 ( .A(n2629), .B(n2628), .Z(n2633) );
  NAND U3279 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U3280 ( .A(n2633), .B(n2632), .Z(n2641) );
  XNOR U3281 ( .A(n2640), .B(n2641), .Z(n2642) );
  NANDN U3282 ( .A(n2635), .B(n2634), .Z(n2639) );
  NAND U3283 ( .A(n2637), .B(n2636), .Z(n2638) );
  NAND U3284 ( .A(n2639), .B(n2638), .Z(n2643) );
  XOR U3285 ( .A(n2642), .B(n2643), .Z(n2658) );
  XNOR U3286 ( .A(n2658), .B(sreg[1061]), .Z(n2659) );
  XOR U3287 ( .A(n2660), .B(n2659), .Z(c[1061]) );
  NANDN U3288 ( .A(n2641), .B(n2640), .Z(n2645) );
  NANDN U3289 ( .A(n2643), .B(n2642), .Z(n2644) );
  NAND U3290 ( .A(n2645), .B(n2644), .Z(n2667) );
  AND U3291 ( .A(b[2]), .B(a[40]), .Z(n2673) );
  AND U3292 ( .A(a[41]), .B(b[1]), .Z(n2671) );
  AND U3293 ( .A(a[39]), .B(b[3]), .Z(n2670) );
  XOR U3294 ( .A(n2671), .B(n2670), .Z(n2672) );
  XOR U3295 ( .A(n2673), .B(n2672), .Z(n2676) );
  NAND U3296 ( .A(b[0]), .B(a[42]), .Z(n2677) );
  XOR U3297 ( .A(n2676), .B(n2677), .Z(n2679) );
  OR U3298 ( .A(n2647), .B(n2646), .Z(n2651) );
  NANDN U3299 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U3300 ( .A(n2651), .B(n2650), .Z(n2678) );
  XNOR U3301 ( .A(n2679), .B(n2678), .Z(n2664) );
  NANDN U3302 ( .A(n2653), .B(n2652), .Z(n2657) );
  OR U3303 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U3304 ( .A(n2657), .B(n2656), .Z(n2665) );
  XNOR U3305 ( .A(n2664), .B(n2665), .Z(n2666) );
  XOR U3306 ( .A(n2667), .B(n2666), .Z(n2683) );
  NAND U3307 ( .A(n2658), .B(sreg[1061]), .Z(n2662) );
  OR U3308 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U3309 ( .A(n2662), .B(n2661), .Z(n2682) );
  XNOR U3310 ( .A(sreg[1062]), .B(n2682), .Z(n2663) );
  XOR U3311 ( .A(n2683), .B(n2663), .Z(c[1062]) );
  NANDN U3312 ( .A(n2665), .B(n2664), .Z(n2669) );
  NAND U3313 ( .A(n2667), .B(n2666), .Z(n2668) );
  NAND U3314 ( .A(n2669), .B(n2668), .Z(n2690) );
  AND U3315 ( .A(b[2]), .B(a[41]), .Z(n2696) );
  AND U3316 ( .A(a[42]), .B(b[1]), .Z(n2694) );
  AND U3317 ( .A(a[40]), .B(b[3]), .Z(n2693) );
  XOR U3318 ( .A(n2694), .B(n2693), .Z(n2695) );
  XOR U3319 ( .A(n2696), .B(n2695), .Z(n2699) );
  NAND U3320 ( .A(b[0]), .B(a[43]), .Z(n2700) );
  XOR U3321 ( .A(n2699), .B(n2700), .Z(n2702) );
  OR U3322 ( .A(n2671), .B(n2670), .Z(n2675) );
  NANDN U3323 ( .A(n2673), .B(n2672), .Z(n2674) );
  NAND U3324 ( .A(n2675), .B(n2674), .Z(n2701) );
  XNOR U3325 ( .A(n2702), .B(n2701), .Z(n2687) );
  NANDN U3326 ( .A(n2677), .B(n2676), .Z(n2681) );
  OR U3327 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U3328 ( .A(n2681), .B(n2680), .Z(n2688) );
  XNOR U3329 ( .A(n2687), .B(n2688), .Z(n2689) );
  XNOR U3330 ( .A(n2690), .B(n2689), .Z(n2686) );
  XOR U3331 ( .A(n2685), .B(sreg[1063]), .Z(n2684) );
  XOR U3332 ( .A(n2686), .B(n2684), .Z(c[1063]) );
  NANDN U3333 ( .A(n2688), .B(n2687), .Z(n2692) );
  NAND U3334 ( .A(n2690), .B(n2689), .Z(n2691) );
  NAND U3335 ( .A(n2692), .B(n2691), .Z(n2708) );
  AND U3336 ( .A(b[2]), .B(a[42]), .Z(n2714) );
  AND U3337 ( .A(a[43]), .B(b[1]), .Z(n2712) );
  AND U3338 ( .A(a[41]), .B(b[3]), .Z(n2711) );
  XOR U3339 ( .A(n2712), .B(n2711), .Z(n2713) );
  XOR U3340 ( .A(n2714), .B(n2713), .Z(n2717) );
  NAND U3341 ( .A(b[0]), .B(a[44]), .Z(n2718) );
  XOR U3342 ( .A(n2717), .B(n2718), .Z(n2720) );
  OR U3343 ( .A(n2694), .B(n2693), .Z(n2698) );
  NANDN U3344 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U3345 ( .A(n2698), .B(n2697), .Z(n2719) );
  XNOR U3346 ( .A(n2720), .B(n2719), .Z(n2705) );
  NANDN U3347 ( .A(n2700), .B(n2699), .Z(n2704) );
  OR U3348 ( .A(n2702), .B(n2701), .Z(n2703) );
  NAND U3349 ( .A(n2704), .B(n2703), .Z(n2706) );
  XNOR U3350 ( .A(n2705), .B(n2706), .Z(n2707) );
  XNOR U3351 ( .A(n2708), .B(n2707), .Z(n2723) );
  XNOR U3352 ( .A(n2723), .B(sreg[1064]), .Z(n2725) );
  XNOR U3353 ( .A(n2724), .B(n2725), .Z(c[1064]) );
  NANDN U3354 ( .A(n2706), .B(n2705), .Z(n2710) );
  NAND U3355 ( .A(n2708), .B(n2707), .Z(n2709) );
  NAND U3356 ( .A(n2710), .B(n2709), .Z(n2731) );
  AND U3357 ( .A(b[2]), .B(a[43]), .Z(n2737) );
  AND U3358 ( .A(a[44]), .B(b[1]), .Z(n2735) );
  AND U3359 ( .A(a[42]), .B(b[3]), .Z(n2734) );
  XOR U3360 ( .A(n2735), .B(n2734), .Z(n2736) );
  XOR U3361 ( .A(n2737), .B(n2736), .Z(n2740) );
  NAND U3362 ( .A(b[0]), .B(a[45]), .Z(n2741) );
  XOR U3363 ( .A(n2740), .B(n2741), .Z(n2743) );
  OR U3364 ( .A(n2712), .B(n2711), .Z(n2716) );
  NANDN U3365 ( .A(n2714), .B(n2713), .Z(n2715) );
  NAND U3366 ( .A(n2716), .B(n2715), .Z(n2742) );
  XNOR U3367 ( .A(n2743), .B(n2742), .Z(n2728) );
  NANDN U3368 ( .A(n2718), .B(n2717), .Z(n2722) );
  OR U3369 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U3370 ( .A(n2722), .B(n2721), .Z(n2729) );
  XNOR U3371 ( .A(n2728), .B(n2729), .Z(n2730) );
  XNOR U3372 ( .A(n2731), .B(n2730), .Z(n2746) );
  XNOR U3373 ( .A(n2746), .B(sreg[1065]), .Z(n2748) );
  NAND U3374 ( .A(n2723), .B(sreg[1064]), .Z(n2727) );
  NANDN U3375 ( .A(n2725), .B(n2724), .Z(n2726) );
  AND U3376 ( .A(n2727), .B(n2726), .Z(n2747) );
  XOR U3377 ( .A(n2748), .B(n2747), .Z(c[1065]) );
  NANDN U3378 ( .A(n2729), .B(n2728), .Z(n2733) );
  NAND U3379 ( .A(n2731), .B(n2730), .Z(n2732) );
  NAND U3380 ( .A(n2733), .B(n2732), .Z(n2757) );
  AND U3381 ( .A(b[2]), .B(a[44]), .Z(n2763) );
  AND U3382 ( .A(a[45]), .B(b[1]), .Z(n2761) );
  AND U3383 ( .A(a[43]), .B(b[3]), .Z(n2760) );
  XOR U3384 ( .A(n2761), .B(n2760), .Z(n2762) );
  XOR U3385 ( .A(n2763), .B(n2762), .Z(n2766) );
  NAND U3386 ( .A(b[0]), .B(a[46]), .Z(n2767) );
  XOR U3387 ( .A(n2766), .B(n2767), .Z(n2769) );
  OR U3388 ( .A(n2735), .B(n2734), .Z(n2739) );
  NANDN U3389 ( .A(n2737), .B(n2736), .Z(n2738) );
  NAND U3390 ( .A(n2739), .B(n2738), .Z(n2768) );
  XNOR U3391 ( .A(n2769), .B(n2768), .Z(n2754) );
  NANDN U3392 ( .A(n2741), .B(n2740), .Z(n2745) );
  OR U3393 ( .A(n2743), .B(n2742), .Z(n2744) );
  NAND U3394 ( .A(n2745), .B(n2744), .Z(n2755) );
  XNOR U3395 ( .A(n2754), .B(n2755), .Z(n2756) );
  XNOR U3396 ( .A(n2757), .B(n2756), .Z(n2753) );
  NAND U3397 ( .A(n2746), .B(sreg[1065]), .Z(n2750) );
  OR U3398 ( .A(n2748), .B(n2747), .Z(n2749) );
  AND U3399 ( .A(n2750), .B(n2749), .Z(n2752) );
  XNOR U3400 ( .A(n2752), .B(sreg[1066]), .Z(n2751) );
  XOR U3401 ( .A(n2753), .B(n2751), .Z(c[1066]) );
  NANDN U3402 ( .A(n2755), .B(n2754), .Z(n2759) );
  NAND U3403 ( .A(n2757), .B(n2756), .Z(n2758) );
  NAND U3404 ( .A(n2759), .B(n2758), .Z(n2775) );
  AND U3405 ( .A(b[2]), .B(a[45]), .Z(n2781) );
  AND U3406 ( .A(a[46]), .B(b[1]), .Z(n2779) );
  AND U3407 ( .A(a[44]), .B(b[3]), .Z(n2778) );
  XOR U3408 ( .A(n2779), .B(n2778), .Z(n2780) );
  XOR U3409 ( .A(n2781), .B(n2780), .Z(n2784) );
  NAND U3410 ( .A(b[0]), .B(a[47]), .Z(n2785) );
  XOR U3411 ( .A(n2784), .B(n2785), .Z(n2787) );
  OR U3412 ( .A(n2761), .B(n2760), .Z(n2765) );
  NANDN U3413 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U3414 ( .A(n2765), .B(n2764), .Z(n2786) );
  XNOR U3415 ( .A(n2787), .B(n2786), .Z(n2772) );
  NANDN U3416 ( .A(n2767), .B(n2766), .Z(n2771) );
  OR U3417 ( .A(n2769), .B(n2768), .Z(n2770) );
  NAND U3418 ( .A(n2771), .B(n2770), .Z(n2773) );
  XNOR U3419 ( .A(n2772), .B(n2773), .Z(n2774) );
  XNOR U3420 ( .A(n2775), .B(n2774), .Z(n2790) );
  XNOR U3421 ( .A(n2790), .B(sreg[1067]), .Z(n2792) );
  XNOR U3422 ( .A(n2791), .B(n2792), .Z(c[1067]) );
  NANDN U3423 ( .A(n2773), .B(n2772), .Z(n2777) );
  NAND U3424 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3425 ( .A(n2777), .B(n2776), .Z(n2798) );
  AND U3426 ( .A(b[2]), .B(a[46]), .Z(n2804) );
  AND U3427 ( .A(a[47]), .B(b[1]), .Z(n2802) );
  AND U3428 ( .A(a[45]), .B(b[3]), .Z(n2801) );
  XOR U3429 ( .A(n2802), .B(n2801), .Z(n2803) );
  XOR U3430 ( .A(n2804), .B(n2803), .Z(n2807) );
  NAND U3431 ( .A(b[0]), .B(a[48]), .Z(n2808) );
  XOR U3432 ( .A(n2807), .B(n2808), .Z(n2810) );
  OR U3433 ( .A(n2779), .B(n2778), .Z(n2783) );
  NANDN U3434 ( .A(n2781), .B(n2780), .Z(n2782) );
  NAND U3435 ( .A(n2783), .B(n2782), .Z(n2809) );
  XNOR U3436 ( .A(n2810), .B(n2809), .Z(n2795) );
  NANDN U3437 ( .A(n2785), .B(n2784), .Z(n2789) );
  OR U3438 ( .A(n2787), .B(n2786), .Z(n2788) );
  NAND U3439 ( .A(n2789), .B(n2788), .Z(n2796) );
  XNOR U3440 ( .A(n2795), .B(n2796), .Z(n2797) );
  XNOR U3441 ( .A(n2798), .B(n2797), .Z(n2813) );
  XNOR U3442 ( .A(n2813), .B(sreg[1068]), .Z(n2815) );
  NAND U3443 ( .A(n2790), .B(sreg[1067]), .Z(n2794) );
  NANDN U3444 ( .A(n2792), .B(n2791), .Z(n2793) );
  AND U3445 ( .A(n2794), .B(n2793), .Z(n2814) );
  XOR U3446 ( .A(n2815), .B(n2814), .Z(c[1068]) );
  NANDN U3447 ( .A(n2796), .B(n2795), .Z(n2800) );
  NAND U3448 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U3449 ( .A(n2800), .B(n2799), .Z(n2821) );
  AND U3450 ( .A(b[2]), .B(a[47]), .Z(n2827) );
  AND U3451 ( .A(a[48]), .B(b[1]), .Z(n2825) );
  AND U3452 ( .A(a[46]), .B(b[3]), .Z(n2824) );
  XOR U3453 ( .A(n2825), .B(n2824), .Z(n2826) );
  XOR U3454 ( .A(n2827), .B(n2826), .Z(n2830) );
  NAND U3455 ( .A(b[0]), .B(a[49]), .Z(n2831) );
  XOR U3456 ( .A(n2830), .B(n2831), .Z(n2833) );
  OR U3457 ( .A(n2802), .B(n2801), .Z(n2806) );
  NANDN U3458 ( .A(n2804), .B(n2803), .Z(n2805) );
  NAND U3459 ( .A(n2806), .B(n2805), .Z(n2832) );
  XNOR U3460 ( .A(n2833), .B(n2832), .Z(n2818) );
  NANDN U3461 ( .A(n2808), .B(n2807), .Z(n2812) );
  OR U3462 ( .A(n2810), .B(n2809), .Z(n2811) );
  NAND U3463 ( .A(n2812), .B(n2811), .Z(n2819) );
  XNOR U3464 ( .A(n2818), .B(n2819), .Z(n2820) );
  XNOR U3465 ( .A(n2821), .B(n2820), .Z(n2836) );
  XNOR U3466 ( .A(n2836), .B(sreg[1069]), .Z(n2838) );
  NAND U3467 ( .A(n2813), .B(sreg[1068]), .Z(n2817) );
  OR U3468 ( .A(n2815), .B(n2814), .Z(n2816) );
  AND U3469 ( .A(n2817), .B(n2816), .Z(n2837) );
  XOR U3470 ( .A(n2838), .B(n2837), .Z(c[1069]) );
  NANDN U3471 ( .A(n2819), .B(n2818), .Z(n2823) );
  NAND U3472 ( .A(n2821), .B(n2820), .Z(n2822) );
  NAND U3473 ( .A(n2823), .B(n2822), .Z(n2844) );
  AND U3474 ( .A(b[2]), .B(a[48]), .Z(n2850) );
  AND U3475 ( .A(a[49]), .B(b[1]), .Z(n2848) );
  AND U3476 ( .A(a[47]), .B(b[3]), .Z(n2847) );
  XOR U3477 ( .A(n2848), .B(n2847), .Z(n2849) );
  XOR U3478 ( .A(n2850), .B(n2849), .Z(n2853) );
  NAND U3479 ( .A(b[0]), .B(a[50]), .Z(n2854) );
  XOR U3480 ( .A(n2853), .B(n2854), .Z(n2856) );
  OR U3481 ( .A(n2825), .B(n2824), .Z(n2829) );
  NANDN U3482 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U3483 ( .A(n2829), .B(n2828), .Z(n2855) );
  XNOR U3484 ( .A(n2856), .B(n2855), .Z(n2841) );
  NANDN U3485 ( .A(n2831), .B(n2830), .Z(n2835) );
  OR U3486 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U3487 ( .A(n2835), .B(n2834), .Z(n2842) );
  XNOR U3488 ( .A(n2841), .B(n2842), .Z(n2843) );
  XNOR U3489 ( .A(n2844), .B(n2843), .Z(n2859) );
  XNOR U3490 ( .A(n2859), .B(sreg[1070]), .Z(n2861) );
  NAND U3491 ( .A(n2836), .B(sreg[1069]), .Z(n2840) );
  OR U3492 ( .A(n2838), .B(n2837), .Z(n2839) );
  AND U3493 ( .A(n2840), .B(n2839), .Z(n2860) );
  XOR U3494 ( .A(n2861), .B(n2860), .Z(c[1070]) );
  NANDN U3495 ( .A(n2842), .B(n2841), .Z(n2846) );
  NAND U3496 ( .A(n2844), .B(n2843), .Z(n2845) );
  NAND U3497 ( .A(n2846), .B(n2845), .Z(n2868) );
  AND U3498 ( .A(b[2]), .B(a[49]), .Z(n2874) );
  AND U3499 ( .A(a[50]), .B(b[1]), .Z(n2872) );
  AND U3500 ( .A(a[48]), .B(b[3]), .Z(n2871) );
  XOR U3501 ( .A(n2872), .B(n2871), .Z(n2873) );
  XOR U3502 ( .A(n2874), .B(n2873), .Z(n2877) );
  NAND U3503 ( .A(b[0]), .B(a[51]), .Z(n2878) );
  XOR U3504 ( .A(n2877), .B(n2878), .Z(n2880) );
  OR U3505 ( .A(n2848), .B(n2847), .Z(n2852) );
  NANDN U3506 ( .A(n2850), .B(n2849), .Z(n2851) );
  NAND U3507 ( .A(n2852), .B(n2851), .Z(n2879) );
  XNOR U3508 ( .A(n2880), .B(n2879), .Z(n2865) );
  NANDN U3509 ( .A(n2854), .B(n2853), .Z(n2858) );
  OR U3510 ( .A(n2856), .B(n2855), .Z(n2857) );
  NAND U3511 ( .A(n2858), .B(n2857), .Z(n2866) );
  XNOR U3512 ( .A(n2865), .B(n2866), .Z(n2867) );
  XNOR U3513 ( .A(n2868), .B(n2867), .Z(n2884) );
  NAND U3514 ( .A(n2859), .B(sreg[1070]), .Z(n2863) );
  OR U3515 ( .A(n2861), .B(n2860), .Z(n2862) );
  AND U3516 ( .A(n2863), .B(n2862), .Z(n2883) );
  XNOR U3517 ( .A(n2883), .B(sreg[1071]), .Z(n2864) );
  XOR U3518 ( .A(n2884), .B(n2864), .Z(c[1071]) );
  NANDN U3519 ( .A(n2866), .B(n2865), .Z(n2870) );
  NAND U3520 ( .A(n2868), .B(n2867), .Z(n2869) );
  NAND U3521 ( .A(n2870), .B(n2869), .Z(n2891) );
  AND U3522 ( .A(b[2]), .B(a[50]), .Z(n2897) );
  AND U3523 ( .A(a[51]), .B(b[1]), .Z(n2895) );
  AND U3524 ( .A(a[49]), .B(b[3]), .Z(n2894) );
  XOR U3525 ( .A(n2895), .B(n2894), .Z(n2896) );
  XOR U3526 ( .A(n2897), .B(n2896), .Z(n2900) );
  NAND U3527 ( .A(b[0]), .B(a[52]), .Z(n2901) );
  XOR U3528 ( .A(n2900), .B(n2901), .Z(n2903) );
  OR U3529 ( .A(n2872), .B(n2871), .Z(n2876) );
  NANDN U3530 ( .A(n2874), .B(n2873), .Z(n2875) );
  NAND U3531 ( .A(n2876), .B(n2875), .Z(n2902) );
  XNOR U3532 ( .A(n2903), .B(n2902), .Z(n2888) );
  NANDN U3533 ( .A(n2878), .B(n2877), .Z(n2882) );
  OR U3534 ( .A(n2880), .B(n2879), .Z(n2881) );
  NAND U3535 ( .A(n2882), .B(n2881), .Z(n2889) );
  XNOR U3536 ( .A(n2888), .B(n2889), .Z(n2890) );
  XOR U3537 ( .A(n2891), .B(n2890), .Z(n2887) );
  XOR U3538 ( .A(sreg[1072]), .B(n2886), .Z(n2885) );
  XOR U3539 ( .A(n2887), .B(n2885), .Z(c[1072]) );
  NANDN U3540 ( .A(n2889), .B(n2888), .Z(n2893) );
  NAND U3541 ( .A(n2891), .B(n2890), .Z(n2892) );
  NAND U3542 ( .A(n2893), .B(n2892), .Z(n2909) );
  AND U3543 ( .A(b[2]), .B(a[51]), .Z(n2915) );
  AND U3544 ( .A(a[52]), .B(b[1]), .Z(n2913) );
  AND U3545 ( .A(a[50]), .B(b[3]), .Z(n2912) );
  XOR U3546 ( .A(n2913), .B(n2912), .Z(n2914) );
  XOR U3547 ( .A(n2915), .B(n2914), .Z(n2918) );
  NAND U3548 ( .A(b[0]), .B(a[53]), .Z(n2919) );
  XOR U3549 ( .A(n2918), .B(n2919), .Z(n2921) );
  OR U3550 ( .A(n2895), .B(n2894), .Z(n2899) );
  NANDN U3551 ( .A(n2897), .B(n2896), .Z(n2898) );
  NAND U3552 ( .A(n2899), .B(n2898), .Z(n2920) );
  XNOR U3553 ( .A(n2921), .B(n2920), .Z(n2906) );
  NANDN U3554 ( .A(n2901), .B(n2900), .Z(n2905) );
  OR U3555 ( .A(n2903), .B(n2902), .Z(n2904) );
  NAND U3556 ( .A(n2905), .B(n2904), .Z(n2907) );
  XNOR U3557 ( .A(n2906), .B(n2907), .Z(n2908) );
  XNOR U3558 ( .A(n2909), .B(n2908), .Z(n2924) );
  XNOR U3559 ( .A(n2924), .B(sreg[1073]), .Z(n2925) );
  XOR U3560 ( .A(n2926), .B(n2925), .Z(c[1073]) );
  NANDN U3561 ( .A(n2907), .B(n2906), .Z(n2911) );
  NAND U3562 ( .A(n2909), .B(n2908), .Z(n2910) );
  NAND U3563 ( .A(n2911), .B(n2910), .Z(n2932) );
  AND U3564 ( .A(b[2]), .B(a[52]), .Z(n2938) );
  AND U3565 ( .A(a[53]), .B(b[1]), .Z(n2936) );
  AND U3566 ( .A(a[51]), .B(b[3]), .Z(n2935) );
  XOR U3567 ( .A(n2936), .B(n2935), .Z(n2937) );
  XOR U3568 ( .A(n2938), .B(n2937), .Z(n2941) );
  NAND U3569 ( .A(b[0]), .B(a[54]), .Z(n2942) );
  XOR U3570 ( .A(n2941), .B(n2942), .Z(n2944) );
  OR U3571 ( .A(n2913), .B(n2912), .Z(n2917) );
  NANDN U3572 ( .A(n2915), .B(n2914), .Z(n2916) );
  NAND U3573 ( .A(n2917), .B(n2916), .Z(n2943) );
  XNOR U3574 ( .A(n2944), .B(n2943), .Z(n2929) );
  NANDN U3575 ( .A(n2919), .B(n2918), .Z(n2923) );
  OR U3576 ( .A(n2921), .B(n2920), .Z(n2922) );
  NAND U3577 ( .A(n2923), .B(n2922), .Z(n2930) );
  XNOR U3578 ( .A(n2929), .B(n2930), .Z(n2931) );
  XNOR U3579 ( .A(n2932), .B(n2931), .Z(n2947) );
  XOR U3580 ( .A(sreg[1074]), .B(n2947), .Z(n2948) );
  NAND U3581 ( .A(n2924), .B(sreg[1073]), .Z(n2928) );
  OR U3582 ( .A(n2926), .B(n2925), .Z(n2927) );
  NAND U3583 ( .A(n2928), .B(n2927), .Z(n2949) );
  XOR U3584 ( .A(n2948), .B(n2949), .Z(c[1074]) );
  NANDN U3585 ( .A(n2930), .B(n2929), .Z(n2934) );
  NAND U3586 ( .A(n2932), .B(n2931), .Z(n2933) );
  NAND U3587 ( .A(n2934), .B(n2933), .Z(n2958) );
  AND U3588 ( .A(b[2]), .B(a[53]), .Z(n2964) );
  AND U3589 ( .A(a[54]), .B(b[1]), .Z(n2962) );
  AND U3590 ( .A(a[52]), .B(b[3]), .Z(n2961) );
  XOR U3591 ( .A(n2962), .B(n2961), .Z(n2963) );
  XOR U3592 ( .A(n2964), .B(n2963), .Z(n2967) );
  NAND U3593 ( .A(b[0]), .B(a[55]), .Z(n2968) );
  XOR U3594 ( .A(n2967), .B(n2968), .Z(n2970) );
  OR U3595 ( .A(n2936), .B(n2935), .Z(n2940) );
  NANDN U3596 ( .A(n2938), .B(n2937), .Z(n2939) );
  NAND U3597 ( .A(n2940), .B(n2939), .Z(n2969) );
  XNOR U3598 ( .A(n2970), .B(n2969), .Z(n2955) );
  NANDN U3599 ( .A(n2942), .B(n2941), .Z(n2946) );
  OR U3600 ( .A(n2944), .B(n2943), .Z(n2945) );
  NAND U3601 ( .A(n2946), .B(n2945), .Z(n2956) );
  XNOR U3602 ( .A(n2955), .B(n2956), .Z(n2957) );
  XOR U3603 ( .A(n2958), .B(n2957), .Z(n2954) );
  OR U3604 ( .A(n2947), .B(sreg[1074]), .Z(n2951) );
  NANDN U3605 ( .A(n2949), .B(n2948), .Z(n2950) );
  AND U3606 ( .A(n2951), .B(n2950), .Z(n2953) );
  XNOR U3607 ( .A(sreg[1075]), .B(n2953), .Z(n2952) );
  XOR U3608 ( .A(n2954), .B(n2952), .Z(c[1075]) );
  NANDN U3609 ( .A(n2956), .B(n2955), .Z(n2960) );
  NAND U3610 ( .A(n2958), .B(n2957), .Z(n2959) );
  NAND U3611 ( .A(n2960), .B(n2959), .Z(n2976) );
  AND U3612 ( .A(b[2]), .B(a[54]), .Z(n2982) );
  AND U3613 ( .A(a[55]), .B(b[1]), .Z(n2980) );
  AND U3614 ( .A(a[53]), .B(b[3]), .Z(n2979) );
  XOR U3615 ( .A(n2980), .B(n2979), .Z(n2981) );
  XOR U3616 ( .A(n2982), .B(n2981), .Z(n2985) );
  NAND U3617 ( .A(b[0]), .B(a[56]), .Z(n2986) );
  XOR U3618 ( .A(n2985), .B(n2986), .Z(n2988) );
  OR U3619 ( .A(n2962), .B(n2961), .Z(n2966) );
  NANDN U3620 ( .A(n2964), .B(n2963), .Z(n2965) );
  NAND U3621 ( .A(n2966), .B(n2965), .Z(n2987) );
  XNOR U3622 ( .A(n2988), .B(n2987), .Z(n2973) );
  NANDN U3623 ( .A(n2968), .B(n2967), .Z(n2972) );
  OR U3624 ( .A(n2970), .B(n2969), .Z(n2971) );
  NAND U3625 ( .A(n2972), .B(n2971), .Z(n2974) );
  XNOR U3626 ( .A(n2973), .B(n2974), .Z(n2975) );
  XNOR U3627 ( .A(n2976), .B(n2975), .Z(n2991) );
  XNOR U3628 ( .A(n2991), .B(sreg[1076]), .Z(n2992) );
  XOR U3629 ( .A(n2993), .B(n2992), .Z(c[1076]) );
  NANDN U3630 ( .A(n2974), .B(n2973), .Z(n2978) );
  NAND U3631 ( .A(n2976), .B(n2975), .Z(n2977) );
  NAND U3632 ( .A(n2978), .B(n2977), .Z(n2999) );
  AND U3633 ( .A(b[2]), .B(a[55]), .Z(n3005) );
  AND U3634 ( .A(a[56]), .B(b[1]), .Z(n3003) );
  AND U3635 ( .A(a[54]), .B(b[3]), .Z(n3002) );
  XOR U3636 ( .A(n3003), .B(n3002), .Z(n3004) );
  XOR U3637 ( .A(n3005), .B(n3004), .Z(n3008) );
  NAND U3638 ( .A(b[0]), .B(a[57]), .Z(n3009) );
  XOR U3639 ( .A(n3008), .B(n3009), .Z(n3011) );
  OR U3640 ( .A(n2980), .B(n2979), .Z(n2984) );
  NANDN U3641 ( .A(n2982), .B(n2981), .Z(n2983) );
  NAND U3642 ( .A(n2984), .B(n2983), .Z(n3010) );
  XNOR U3643 ( .A(n3011), .B(n3010), .Z(n2996) );
  NANDN U3644 ( .A(n2986), .B(n2985), .Z(n2990) );
  OR U3645 ( .A(n2988), .B(n2987), .Z(n2989) );
  NAND U3646 ( .A(n2990), .B(n2989), .Z(n2997) );
  XNOR U3647 ( .A(n2996), .B(n2997), .Z(n2998) );
  XNOR U3648 ( .A(n2999), .B(n2998), .Z(n3014) );
  XNOR U3649 ( .A(n3014), .B(sreg[1077]), .Z(n3016) );
  NAND U3650 ( .A(n2991), .B(sreg[1076]), .Z(n2995) );
  OR U3651 ( .A(n2993), .B(n2992), .Z(n2994) );
  AND U3652 ( .A(n2995), .B(n2994), .Z(n3015) );
  XOR U3653 ( .A(n3016), .B(n3015), .Z(c[1077]) );
  NANDN U3654 ( .A(n2997), .B(n2996), .Z(n3001) );
  NAND U3655 ( .A(n2999), .B(n2998), .Z(n3000) );
  NAND U3656 ( .A(n3001), .B(n3000), .Z(n3023) );
  AND U3657 ( .A(b[2]), .B(a[56]), .Z(n3029) );
  AND U3658 ( .A(a[57]), .B(b[1]), .Z(n3027) );
  AND U3659 ( .A(a[55]), .B(b[3]), .Z(n3026) );
  XOR U3660 ( .A(n3027), .B(n3026), .Z(n3028) );
  XOR U3661 ( .A(n3029), .B(n3028), .Z(n3032) );
  NAND U3662 ( .A(b[0]), .B(a[58]), .Z(n3033) );
  XOR U3663 ( .A(n3032), .B(n3033), .Z(n3035) );
  OR U3664 ( .A(n3003), .B(n3002), .Z(n3007) );
  NANDN U3665 ( .A(n3005), .B(n3004), .Z(n3006) );
  NAND U3666 ( .A(n3007), .B(n3006), .Z(n3034) );
  XNOR U3667 ( .A(n3035), .B(n3034), .Z(n3020) );
  NANDN U3668 ( .A(n3009), .B(n3008), .Z(n3013) );
  OR U3669 ( .A(n3011), .B(n3010), .Z(n3012) );
  NAND U3670 ( .A(n3013), .B(n3012), .Z(n3021) );
  XNOR U3671 ( .A(n3020), .B(n3021), .Z(n3022) );
  XOR U3672 ( .A(n3023), .B(n3022), .Z(n3039) );
  NAND U3673 ( .A(n3014), .B(sreg[1077]), .Z(n3018) );
  OR U3674 ( .A(n3016), .B(n3015), .Z(n3017) );
  NAND U3675 ( .A(n3018), .B(n3017), .Z(n3038) );
  XNOR U3676 ( .A(sreg[1078]), .B(n3038), .Z(n3019) );
  XOR U3677 ( .A(n3039), .B(n3019), .Z(c[1078]) );
  NANDN U3678 ( .A(n3021), .B(n3020), .Z(n3025) );
  NAND U3679 ( .A(n3023), .B(n3022), .Z(n3024) );
  NAND U3680 ( .A(n3025), .B(n3024), .Z(n3046) );
  AND U3681 ( .A(b[2]), .B(a[57]), .Z(n3052) );
  AND U3682 ( .A(a[58]), .B(b[1]), .Z(n3050) );
  AND U3683 ( .A(a[56]), .B(b[3]), .Z(n3049) );
  XOR U3684 ( .A(n3050), .B(n3049), .Z(n3051) );
  XOR U3685 ( .A(n3052), .B(n3051), .Z(n3055) );
  NAND U3686 ( .A(b[0]), .B(a[59]), .Z(n3056) );
  XOR U3687 ( .A(n3055), .B(n3056), .Z(n3058) );
  OR U3688 ( .A(n3027), .B(n3026), .Z(n3031) );
  NANDN U3689 ( .A(n3029), .B(n3028), .Z(n3030) );
  NAND U3690 ( .A(n3031), .B(n3030), .Z(n3057) );
  XNOR U3691 ( .A(n3058), .B(n3057), .Z(n3043) );
  NANDN U3692 ( .A(n3033), .B(n3032), .Z(n3037) );
  OR U3693 ( .A(n3035), .B(n3034), .Z(n3036) );
  NAND U3694 ( .A(n3037), .B(n3036), .Z(n3044) );
  XNOR U3695 ( .A(n3043), .B(n3044), .Z(n3045) );
  XOR U3696 ( .A(n3046), .B(n3045), .Z(n3042) );
  XNOR U3697 ( .A(sreg[1079]), .B(n3041), .Z(n3040) );
  XOR U3698 ( .A(n3042), .B(n3040), .Z(c[1079]) );
  NANDN U3699 ( .A(n3044), .B(n3043), .Z(n3048) );
  NAND U3700 ( .A(n3046), .B(n3045), .Z(n3047) );
  NAND U3701 ( .A(n3048), .B(n3047), .Z(n3064) );
  AND U3702 ( .A(b[2]), .B(a[58]), .Z(n3070) );
  AND U3703 ( .A(a[59]), .B(b[1]), .Z(n3068) );
  AND U3704 ( .A(a[57]), .B(b[3]), .Z(n3067) );
  XOR U3705 ( .A(n3068), .B(n3067), .Z(n3069) );
  XOR U3706 ( .A(n3070), .B(n3069), .Z(n3073) );
  NAND U3707 ( .A(b[0]), .B(a[60]), .Z(n3074) );
  XOR U3708 ( .A(n3073), .B(n3074), .Z(n3076) );
  OR U3709 ( .A(n3050), .B(n3049), .Z(n3054) );
  NANDN U3710 ( .A(n3052), .B(n3051), .Z(n3053) );
  NAND U3711 ( .A(n3054), .B(n3053), .Z(n3075) );
  XNOR U3712 ( .A(n3076), .B(n3075), .Z(n3061) );
  NANDN U3713 ( .A(n3056), .B(n3055), .Z(n3060) );
  OR U3714 ( .A(n3058), .B(n3057), .Z(n3059) );
  NAND U3715 ( .A(n3060), .B(n3059), .Z(n3062) );
  XNOR U3716 ( .A(n3061), .B(n3062), .Z(n3063) );
  XNOR U3717 ( .A(n3064), .B(n3063), .Z(n3079) );
  XNOR U3718 ( .A(n3079), .B(sreg[1080]), .Z(n3080) );
  XOR U3719 ( .A(n3081), .B(n3080), .Z(c[1080]) );
  NANDN U3720 ( .A(n3062), .B(n3061), .Z(n3066) );
  NAND U3721 ( .A(n3064), .B(n3063), .Z(n3065) );
  NAND U3722 ( .A(n3066), .B(n3065), .Z(n3088) );
  AND U3723 ( .A(b[2]), .B(a[59]), .Z(n3094) );
  AND U3724 ( .A(a[60]), .B(b[1]), .Z(n3092) );
  AND U3725 ( .A(a[58]), .B(b[3]), .Z(n3091) );
  XOR U3726 ( .A(n3092), .B(n3091), .Z(n3093) );
  XOR U3727 ( .A(n3094), .B(n3093), .Z(n3097) );
  NAND U3728 ( .A(b[0]), .B(a[61]), .Z(n3098) );
  XOR U3729 ( .A(n3097), .B(n3098), .Z(n3100) );
  OR U3730 ( .A(n3068), .B(n3067), .Z(n3072) );
  NANDN U3731 ( .A(n3070), .B(n3069), .Z(n3071) );
  NAND U3732 ( .A(n3072), .B(n3071), .Z(n3099) );
  XNOR U3733 ( .A(n3100), .B(n3099), .Z(n3085) );
  NANDN U3734 ( .A(n3074), .B(n3073), .Z(n3078) );
  OR U3735 ( .A(n3076), .B(n3075), .Z(n3077) );
  NAND U3736 ( .A(n3078), .B(n3077), .Z(n3086) );
  XNOR U3737 ( .A(n3085), .B(n3086), .Z(n3087) );
  XOR U3738 ( .A(n3088), .B(n3087), .Z(n3104) );
  NAND U3739 ( .A(n3079), .B(sreg[1080]), .Z(n3083) );
  OR U3740 ( .A(n3081), .B(n3080), .Z(n3082) );
  NAND U3741 ( .A(n3083), .B(n3082), .Z(n3103) );
  XNOR U3742 ( .A(sreg[1081]), .B(n3103), .Z(n3084) );
  XOR U3743 ( .A(n3104), .B(n3084), .Z(c[1081]) );
  NANDN U3744 ( .A(n3086), .B(n3085), .Z(n3090) );
  NAND U3745 ( .A(n3088), .B(n3087), .Z(n3089) );
  NAND U3746 ( .A(n3090), .B(n3089), .Z(n3111) );
  AND U3747 ( .A(b[2]), .B(a[60]), .Z(n3117) );
  AND U3748 ( .A(a[61]), .B(b[1]), .Z(n3115) );
  AND U3749 ( .A(a[59]), .B(b[3]), .Z(n3114) );
  XOR U3750 ( .A(n3115), .B(n3114), .Z(n3116) );
  XOR U3751 ( .A(n3117), .B(n3116), .Z(n3120) );
  NAND U3752 ( .A(b[0]), .B(a[62]), .Z(n3121) );
  XOR U3753 ( .A(n3120), .B(n3121), .Z(n3123) );
  OR U3754 ( .A(n3092), .B(n3091), .Z(n3096) );
  NANDN U3755 ( .A(n3094), .B(n3093), .Z(n3095) );
  NAND U3756 ( .A(n3096), .B(n3095), .Z(n3122) );
  XNOR U3757 ( .A(n3123), .B(n3122), .Z(n3108) );
  NANDN U3758 ( .A(n3098), .B(n3097), .Z(n3102) );
  OR U3759 ( .A(n3100), .B(n3099), .Z(n3101) );
  NAND U3760 ( .A(n3102), .B(n3101), .Z(n3109) );
  XNOR U3761 ( .A(n3108), .B(n3109), .Z(n3110) );
  XOR U3762 ( .A(n3111), .B(n3110), .Z(n3107) );
  XNOR U3763 ( .A(sreg[1082]), .B(n3106), .Z(n3105) );
  XOR U3764 ( .A(n3107), .B(n3105), .Z(c[1082]) );
  NANDN U3765 ( .A(n3109), .B(n3108), .Z(n3113) );
  NAND U3766 ( .A(n3111), .B(n3110), .Z(n3112) );
  NAND U3767 ( .A(n3113), .B(n3112), .Z(n3129) );
  AND U3768 ( .A(b[2]), .B(a[61]), .Z(n3135) );
  AND U3769 ( .A(a[62]), .B(b[1]), .Z(n3133) );
  AND U3770 ( .A(a[60]), .B(b[3]), .Z(n3132) );
  XOR U3771 ( .A(n3133), .B(n3132), .Z(n3134) );
  XOR U3772 ( .A(n3135), .B(n3134), .Z(n3138) );
  NAND U3773 ( .A(b[0]), .B(a[63]), .Z(n3139) );
  XOR U3774 ( .A(n3138), .B(n3139), .Z(n3141) );
  OR U3775 ( .A(n3115), .B(n3114), .Z(n3119) );
  NANDN U3776 ( .A(n3117), .B(n3116), .Z(n3118) );
  NAND U3777 ( .A(n3119), .B(n3118), .Z(n3140) );
  XNOR U3778 ( .A(n3141), .B(n3140), .Z(n3126) );
  NANDN U3779 ( .A(n3121), .B(n3120), .Z(n3125) );
  OR U3780 ( .A(n3123), .B(n3122), .Z(n3124) );
  NAND U3781 ( .A(n3125), .B(n3124), .Z(n3127) );
  XNOR U3782 ( .A(n3126), .B(n3127), .Z(n3128) );
  XNOR U3783 ( .A(n3129), .B(n3128), .Z(n3144) );
  XNOR U3784 ( .A(n3144), .B(sreg[1083]), .Z(n3145) );
  XOR U3785 ( .A(n3146), .B(n3145), .Z(c[1083]) );
  NANDN U3786 ( .A(n3127), .B(n3126), .Z(n3131) );
  NAND U3787 ( .A(n3129), .B(n3128), .Z(n3130) );
  NAND U3788 ( .A(n3131), .B(n3130), .Z(n3152) );
  AND U3789 ( .A(b[2]), .B(a[62]), .Z(n3164) );
  AND U3790 ( .A(a[63]), .B(b[1]), .Z(n3162) );
  AND U3791 ( .A(a[61]), .B(b[3]), .Z(n3161) );
  XOR U3792 ( .A(n3162), .B(n3161), .Z(n3163) );
  XOR U3793 ( .A(n3164), .B(n3163), .Z(n3155) );
  NAND U3794 ( .A(b[0]), .B(a[64]), .Z(n3156) );
  XOR U3795 ( .A(n3155), .B(n3156), .Z(n3158) );
  OR U3796 ( .A(n3133), .B(n3132), .Z(n3137) );
  NANDN U3797 ( .A(n3135), .B(n3134), .Z(n3136) );
  NAND U3798 ( .A(n3137), .B(n3136), .Z(n3157) );
  XNOR U3799 ( .A(n3158), .B(n3157), .Z(n3149) );
  NANDN U3800 ( .A(n3139), .B(n3138), .Z(n3143) );
  OR U3801 ( .A(n3141), .B(n3140), .Z(n3142) );
  NAND U3802 ( .A(n3143), .B(n3142), .Z(n3150) );
  XNOR U3803 ( .A(n3149), .B(n3150), .Z(n3151) );
  XNOR U3804 ( .A(n3152), .B(n3151), .Z(n3168) );
  XOR U3805 ( .A(sreg[1084]), .B(n3168), .Z(n3169) );
  NAND U3806 ( .A(n3144), .B(sreg[1083]), .Z(n3148) );
  OR U3807 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U3808 ( .A(n3148), .B(n3147), .Z(n3170) );
  XOR U3809 ( .A(n3169), .B(n3170), .Z(c[1084]) );
  NANDN U3810 ( .A(n3150), .B(n3149), .Z(n3154) );
  NAND U3811 ( .A(n3152), .B(n3151), .Z(n3153) );
  AND U3812 ( .A(n3154), .B(n3153), .Z(n3176) );
  NANDN U3813 ( .A(n3156), .B(n3155), .Z(n3160) );
  OR U3814 ( .A(n3158), .B(n3157), .Z(n3159) );
  AND U3815 ( .A(n3160), .B(n3159), .Z(n3175) );
  AND U3816 ( .A(b[2]), .B(a[63]), .Z(n3180) );
  AND U3817 ( .A(a[64]), .B(b[1]), .Z(n3178) );
  AND U3818 ( .A(a[62]), .B(b[3]), .Z(n3177) );
  XOR U3819 ( .A(n3178), .B(n3177), .Z(n3179) );
  XOR U3820 ( .A(n3180), .B(n3179), .Z(n3183) );
  NAND U3821 ( .A(b[0]), .B(a[65]), .Z(n3184) );
  XOR U3822 ( .A(n3183), .B(n3184), .Z(n3186) );
  OR U3823 ( .A(n3162), .B(n3161), .Z(n3166) );
  NANDN U3824 ( .A(n3164), .B(n3163), .Z(n3165) );
  NAND U3825 ( .A(n3166), .B(n3165), .Z(n3185) );
  XOR U3826 ( .A(n3186), .B(n3185), .Z(n3174) );
  XNOR U3827 ( .A(n3175), .B(n3174), .Z(n3167) );
  XOR U3828 ( .A(n3176), .B(n3167), .Z(n3190) );
  OR U3829 ( .A(n3168), .B(sreg[1084]), .Z(n3172) );
  NANDN U3830 ( .A(n3170), .B(n3169), .Z(n3171) );
  AND U3831 ( .A(n3172), .B(n3171), .Z(n3189) );
  XNOR U3832 ( .A(sreg[1085]), .B(n3189), .Z(n3173) );
  XNOR U3833 ( .A(n3190), .B(n3173), .Z(c[1085]) );
  AND U3834 ( .A(b[2]), .B(a[64]), .Z(n3203) );
  AND U3835 ( .A(a[65]), .B(b[1]), .Z(n3201) );
  AND U3836 ( .A(a[63]), .B(b[3]), .Z(n3200) );
  XOR U3837 ( .A(n3201), .B(n3200), .Z(n3202) );
  XOR U3838 ( .A(n3203), .B(n3202), .Z(n3206) );
  NAND U3839 ( .A(b[0]), .B(a[66]), .Z(n3207) );
  XOR U3840 ( .A(n3206), .B(n3207), .Z(n3209) );
  OR U3841 ( .A(n3178), .B(n3177), .Z(n3182) );
  NANDN U3842 ( .A(n3180), .B(n3179), .Z(n3181) );
  NAND U3843 ( .A(n3182), .B(n3181), .Z(n3208) );
  XNOR U3844 ( .A(n3209), .B(n3208), .Z(n3194) );
  NANDN U3845 ( .A(n3184), .B(n3183), .Z(n3188) );
  OR U3846 ( .A(n3186), .B(n3185), .Z(n3187) );
  NAND U3847 ( .A(n3188), .B(n3187), .Z(n3195) );
  XNOR U3848 ( .A(n3194), .B(n3195), .Z(n3196) );
  XNOR U3849 ( .A(n3197), .B(n3196), .Z(n3193) );
  XOR U3850 ( .A(n3192), .B(sreg[1086]), .Z(n3191) );
  XNOR U3851 ( .A(n3193), .B(n3191), .Z(c[1086]) );
  NANDN U3852 ( .A(n3195), .B(n3194), .Z(n3199) );
  NANDN U3853 ( .A(n3197), .B(n3196), .Z(n3198) );
  NAND U3854 ( .A(n3199), .B(n3198), .Z(n3215) );
  AND U3855 ( .A(b[2]), .B(a[65]), .Z(n3221) );
  AND U3856 ( .A(a[66]), .B(b[1]), .Z(n3219) );
  AND U3857 ( .A(a[64]), .B(b[3]), .Z(n3218) );
  XOR U3858 ( .A(n3219), .B(n3218), .Z(n3220) );
  XOR U3859 ( .A(n3221), .B(n3220), .Z(n3224) );
  NAND U3860 ( .A(b[0]), .B(a[67]), .Z(n3225) );
  XOR U3861 ( .A(n3224), .B(n3225), .Z(n3227) );
  OR U3862 ( .A(n3201), .B(n3200), .Z(n3205) );
  NANDN U3863 ( .A(n3203), .B(n3202), .Z(n3204) );
  NAND U3864 ( .A(n3205), .B(n3204), .Z(n3226) );
  XNOR U3865 ( .A(n3227), .B(n3226), .Z(n3212) );
  NANDN U3866 ( .A(n3207), .B(n3206), .Z(n3211) );
  OR U3867 ( .A(n3209), .B(n3208), .Z(n3210) );
  NAND U3868 ( .A(n3211), .B(n3210), .Z(n3213) );
  XNOR U3869 ( .A(n3212), .B(n3213), .Z(n3214) );
  XNOR U3870 ( .A(n3215), .B(n3214), .Z(n3231) );
  XNOR U3871 ( .A(n3231), .B(sreg[1087]), .Z(n3233) );
  XNOR U3872 ( .A(n3232), .B(n3233), .Z(c[1087]) );
  NANDN U3873 ( .A(n3213), .B(n3212), .Z(n3217) );
  NAND U3874 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U3875 ( .A(n3217), .B(n3216), .Z(n3238) );
  AND U3876 ( .A(b[2]), .B(a[66]), .Z(n3242) );
  AND U3877 ( .A(a[67]), .B(b[1]), .Z(n3240) );
  AND U3878 ( .A(a[65]), .B(b[3]), .Z(n3239) );
  XOR U3879 ( .A(n3240), .B(n3239), .Z(n3241) );
  XOR U3880 ( .A(n3242), .B(n3241), .Z(n3245) );
  NAND U3881 ( .A(b[0]), .B(a[68]), .Z(n3246) );
  XOR U3882 ( .A(n3245), .B(n3246), .Z(n3247) );
  OR U3883 ( .A(n3219), .B(n3218), .Z(n3223) );
  NANDN U3884 ( .A(n3221), .B(n3220), .Z(n3222) );
  AND U3885 ( .A(n3223), .B(n3222), .Z(n3248) );
  XOR U3886 ( .A(n3247), .B(n3248), .Z(n3236) );
  NANDN U3887 ( .A(n3225), .B(n3224), .Z(n3229) );
  OR U3888 ( .A(n3227), .B(n3226), .Z(n3228) );
  AND U3889 ( .A(n3229), .B(n3228), .Z(n3237) );
  XOR U3890 ( .A(n3236), .B(n3237), .Z(n3230) );
  XOR U3891 ( .A(n3238), .B(n3230), .Z(n3249) );
  XNOR U3892 ( .A(sreg[1088]), .B(n3249), .Z(n3251) );
  NAND U3893 ( .A(n3231), .B(sreg[1087]), .Z(n3235) );
  NANDN U3894 ( .A(n3233), .B(n3232), .Z(n3234) );
  AND U3895 ( .A(n3235), .B(n3234), .Z(n3250) );
  XOR U3896 ( .A(n3251), .B(n3250), .Z(c[1088]) );
  AND U3897 ( .A(b[2]), .B(a[67]), .Z(n3264) );
  AND U3898 ( .A(a[68]), .B(b[1]), .Z(n3262) );
  AND U3899 ( .A(a[66]), .B(b[3]), .Z(n3261) );
  XOR U3900 ( .A(n3262), .B(n3261), .Z(n3263) );
  XOR U3901 ( .A(n3264), .B(n3263), .Z(n3267) );
  NAND U3902 ( .A(b[0]), .B(a[69]), .Z(n3268) );
  XOR U3903 ( .A(n3267), .B(n3268), .Z(n3270) );
  OR U3904 ( .A(n3240), .B(n3239), .Z(n3244) );
  NANDN U3905 ( .A(n3242), .B(n3241), .Z(n3243) );
  NAND U3906 ( .A(n3244), .B(n3243), .Z(n3269) );
  XNOR U3907 ( .A(n3270), .B(n3269), .Z(n3255) );
  XNOR U3908 ( .A(n3255), .B(n3256), .Z(n3258) );
  XOR U3909 ( .A(n3257), .B(n3258), .Z(n3274) );
  NAND U3910 ( .A(sreg[1088]), .B(n3249), .Z(n3253) );
  OR U3911 ( .A(n3251), .B(n3250), .Z(n3252) );
  AND U3912 ( .A(n3253), .B(n3252), .Z(n3273) );
  XNOR U3913 ( .A(n3273), .B(sreg[1089]), .Z(n3254) );
  XNOR U3914 ( .A(n3274), .B(n3254), .Z(c[1089]) );
  NANDN U3915 ( .A(n3256), .B(n3255), .Z(n3260) );
  NAND U3916 ( .A(n3258), .B(n3257), .Z(n3259) );
  NAND U3917 ( .A(n3260), .B(n3259), .Z(n3281) );
  AND U3918 ( .A(b[2]), .B(a[68]), .Z(n3287) );
  AND U3919 ( .A(a[69]), .B(b[1]), .Z(n3285) );
  AND U3920 ( .A(a[67]), .B(b[3]), .Z(n3284) );
  XOR U3921 ( .A(n3285), .B(n3284), .Z(n3286) );
  XOR U3922 ( .A(n3287), .B(n3286), .Z(n3290) );
  NAND U3923 ( .A(b[0]), .B(a[70]), .Z(n3291) );
  XOR U3924 ( .A(n3290), .B(n3291), .Z(n3293) );
  OR U3925 ( .A(n3262), .B(n3261), .Z(n3266) );
  NANDN U3926 ( .A(n3264), .B(n3263), .Z(n3265) );
  NAND U3927 ( .A(n3266), .B(n3265), .Z(n3292) );
  XNOR U3928 ( .A(n3293), .B(n3292), .Z(n3278) );
  NANDN U3929 ( .A(n3268), .B(n3267), .Z(n3272) );
  OR U3930 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U3931 ( .A(n3272), .B(n3271), .Z(n3279) );
  XNOR U3932 ( .A(n3278), .B(n3279), .Z(n3280) );
  XOR U3933 ( .A(n3281), .B(n3280), .Z(n3277) );
  XOR U3934 ( .A(sreg[1090]), .B(n3276), .Z(n3275) );
  XOR U3935 ( .A(n3277), .B(n3275), .Z(c[1090]) );
  NANDN U3936 ( .A(n3279), .B(n3278), .Z(n3283) );
  NAND U3937 ( .A(n3281), .B(n3280), .Z(n3282) );
  NAND U3938 ( .A(n3283), .B(n3282), .Z(n3304) );
  AND U3939 ( .A(b[2]), .B(a[69]), .Z(n3310) );
  AND U3940 ( .A(a[70]), .B(b[1]), .Z(n3308) );
  AND U3941 ( .A(a[68]), .B(b[3]), .Z(n3307) );
  XOR U3942 ( .A(n3308), .B(n3307), .Z(n3309) );
  XOR U3943 ( .A(n3310), .B(n3309), .Z(n3313) );
  NAND U3944 ( .A(b[0]), .B(a[71]), .Z(n3314) );
  XOR U3945 ( .A(n3313), .B(n3314), .Z(n3316) );
  OR U3946 ( .A(n3285), .B(n3284), .Z(n3289) );
  NANDN U3947 ( .A(n3287), .B(n3286), .Z(n3288) );
  NAND U3948 ( .A(n3289), .B(n3288), .Z(n3315) );
  XNOR U3949 ( .A(n3316), .B(n3315), .Z(n3301) );
  NANDN U3950 ( .A(n3291), .B(n3290), .Z(n3295) );
  OR U3951 ( .A(n3293), .B(n3292), .Z(n3294) );
  NAND U3952 ( .A(n3295), .B(n3294), .Z(n3302) );
  XNOR U3953 ( .A(n3301), .B(n3302), .Z(n3303) );
  XNOR U3954 ( .A(n3304), .B(n3303), .Z(n3296) );
  XNOR U3955 ( .A(n3296), .B(sreg[1091]), .Z(n3297) );
  XOR U3956 ( .A(n3298), .B(n3297), .Z(c[1091]) );
  NAND U3957 ( .A(n3296), .B(sreg[1091]), .Z(n3300) );
  OR U3958 ( .A(n3298), .B(n3297), .Z(n3299) );
  AND U3959 ( .A(n3300), .B(n3299), .Z(n3339) );
  NANDN U3960 ( .A(n3302), .B(n3301), .Z(n3306) );
  NAND U3961 ( .A(n3304), .B(n3303), .Z(n3305) );
  NAND U3962 ( .A(n3306), .B(n3305), .Z(n3323) );
  AND U3963 ( .A(b[2]), .B(a[70]), .Z(n3329) );
  AND U3964 ( .A(a[71]), .B(b[1]), .Z(n3327) );
  AND U3965 ( .A(a[69]), .B(b[3]), .Z(n3326) );
  XOR U3966 ( .A(n3327), .B(n3326), .Z(n3328) );
  XOR U3967 ( .A(n3329), .B(n3328), .Z(n3332) );
  NAND U3968 ( .A(b[0]), .B(a[72]), .Z(n3333) );
  XOR U3969 ( .A(n3332), .B(n3333), .Z(n3335) );
  OR U3970 ( .A(n3308), .B(n3307), .Z(n3312) );
  NANDN U3971 ( .A(n3310), .B(n3309), .Z(n3311) );
  NAND U3972 ( .A(n3312), .B(n3311), .Z(n3334) );
  XNOR U3973 ( .A(n3335), .B(n3334), .Z(n3320) );
  NANDN U3974 ( .A(n3314), .B(n3313), .Z(n3318) );
  OR U3975 ( .A(n3316), .B(n3315), .Z(n3317) );
  NAND U3976 ( .A(n3318), .B(n3317), .Z(n3321) );
  XNOR U3977 ( .A(n3320), .B(n3321), .Z(n3322) );
  XNOR U3978 ( .A(n3323), .B(n3322), .Z(n3338) );
  XNOR U3979 ( .A(sreg[1092]), .B(n3338), .Z(n3319) );
  XOR U3980 ( .A(n3339), .B(n3319), .Z(c[1092]) );
  NANDN U3981 ( .A(n3321), .B(n3320), .Z(n3325) );
  NAND U3982 ( .A(n3323), .B(n3322), .Z(n3324) );
  NAND U3983 ( .A(n3325), .B(n3324), .Z(n3346) );
  AND U3984 ( .A(b[2]), .B(a[71]), .Z(n3352) );
  AND U3985 ( .A(a[72]), .B(b[1]), .Z(n3350) );
  AND U3986 ( .A(a[70]), .B(b[3]), .Z(n3349) );
  XOR U3987 ( .A(n3350), .B(n3349), .Z(n3351) );
  XOR U3988 ( .A(n3352), .B(n3351), .Z(n3355) );
  NAND U3989 ( .A(b[0]), .B(a[73]), .Z(n3356) );
  XOR U3990 ( .A(n3355), .B(n3356), .Z(n3358) );
  OR U3991 ( .A(n3327), .B(n3326), .Z(n3331) );
  NANDN U3992 ( .A(n3329), .B(n3328), .Z(n3330) );
  NAND U3993 ( .A(n3331), .B(n3330), .Z(n3357) );
  XNOR U3994 ( .A(n3358), .B(n3357), .Z(n3343) );
  NANDN U3995 ( .A(n3333), .B(n3332), .Z(n3337) );
  OR U3996 ( .A(n3335), .B(n3334), .Z(n3336) );
  NAND U3997 ( .A(n3337), .B(n3336), .Z(n3344) );
  XNOR U3998 ( .A(n3343), .B(n3344), .Z(n3345) );
  XOR U3999 ( .A(n3346), .B(n3345), .Z(n3342) );
  XNOR U4000 ( .A(sreg[1093]), .B(n3341), .Z(n3340) );
  XOR U4001 ( .A(n3342), .B(n3340), .Z(c[1093]) );
  NANDN U4002 ( .A(n3344), .B(n3343), .Z(n3348) );
  NAND U4003 ( .A(n3346), .B(n3345), .Z(n3347) );
  NAND U4004 ( .A(n3348), .B(n3347), .Z(n3364) );
  AND U4005 ( .A(b[2]), .B(a[72]), .Z(n3370) );
  AND U4006 ( .A(a[73]), .B(b[1]), .Z(n3368) );
  AND U4007 ( .A(a[71]), .B(b[3]), .Z(n3367) );
  XOR U4008 ( .A(n3368), .B(n3367), .Z(n3369) );
  XOR U4009 ( .A(n3370), .B(n3369), .Z(n3373) );
  NAND U4010 ( .A(b[0]), .B(a[74]), .Z(n3374) );
  XOR U4011 ( .A(n3373), .B(n3374), .Z(n3376) );
  OR U4012 ( .A(n3350), .B(n3349), .Z(n3354) );
  NANDN U4013 ( .A(n3352), .B(n3351), .Z(n3353) );
  NAND U4014 ( .A(n3354), .B(n3353), .Z(n3375) );
  XNOR U4015 ( .A(n3376), .B(n3375), .Z(n3361) );
  NANDN U4016 ( .A(n3356), .B(n3355), .Z(n3360) );
  OR U4017 ( .A(n3358), .B(n3357), .Z(n3359) );
  NAND U4018 ( .A(n3360), .B(n3359), .Z(n3362) );
  XNOR U4019 ( .A(n3361), .B(n3362), .Z(n3363) );
  XNOR U4020 ( .A(n3364), .B(n3363), .Z(n3379) );
  XNOR U4021 ( .A(n3379), .B(sreg[1094]), .Z(n3380) );
  XOR U4022 ( .A(n3381), .B(n3380), .Z(c[1094]) );
  NANDN U4023 ( .A(n3362), .B(n3361), .Z(n3366) );
  NAND U4024 ( .A(n3364), .B(n3363), .Z(n3365) );
  NAND U4025 ( .A(n3366), .B(n3365), .Z(n3388) );
  AND U4026 ( .A(b[2]), .B(a[73]), .Z(n3394) );
  AND U4027 ( .A(a[74]), .B(b[1]), .Z(n3392) );
  AND U4028 ( .A(a[72]), .B(b[3]), .Z(n3391) );
  XOR U4029 ( .A(n3392), .B(n3391), .Z(n3393) );
  XOR U4030 ( .A(n3394), .B(n3393), .Z(n3397) );
  NAND U4031 ( .A(b[0]), .B(a[75]), .Z(n3398) );
  XOR U4032 ( .A(n3397), .B(n3398), .Z(n3400) );
  OR U4033 ( .A(n3368), .B(n3367), .Z(n3372) );
  NANDN U4034 ( .A(n3370), .B(n3369), .Z(n3371) );
  NAND U4035 ( .A(n3372), .B(n3371), .Z(n3399) );
  XNOR U4036 ( .A(n3400), .B(n3399), .Z(n3385) );
  NANDN U4037 ( .A(n3374), .B(n3373), .Z(n3378) );
  OR U4038 ( .A(n3376), .B(n3375), .Z(n3377) );
  NAND U4039 ( .A(n3378), .B(n3377), .Z(n3386) );
  XNOR U4040 ( .A(n3385), .B(n3386), .Z(n3387) );
  XNOR U4041 ( .A(n3388), .B(n3387), .Z(n3404) );
  NAND U4042 ( .A(n3379), .B(sreg[1094]), .Z(n3383) );
  OR U4043 ( .A(n3381), .B(n3380), .Z(n3382) );
  AND U4044 ( .A(n3383), .B(n3382), .Z(n3403) );
  XNOR U4045 ( .A(n3403), .B(sreg[1095]), .Z(n3384) );
  XOR U4046 ( .A(n3404), .B(n3384), .Z(c[1095]) );
  NANDN U4047 ( .A(n3386), .B(n3385), .Z(n3390) );
  NAND U4048 ( .A(n3388), .B(n3387), .Z(n3389) );
  NAND U4049 ( .A(n3390), .B(n3389), .Z(n3411) );
  AND U4050 ( .A(b[2]), .B(a[74]), .Z(n3417) );
  AND U4051 ( .A(a[75]), .B(b[1]), .Z(n3415) );
  AND U4052 ( .A(a[73]), .B(b[3]), .Z(n3414) );
  XOR U4053 ( .A(n3415), .B(n3414), .Z(n3416) );
  XOR U4054 ( .A(n3417), .B(n3416), .Z(n3420) );
  NAND U4055 ( .A(b[0]), .B(a[76]), .Z(n3421) );
  XOR U4056 ( .A(n3420), .B(n3421), .Z(n3423) );
  OR U4057 ( .A(n3392), .B(n3391), .Z(n3396) );
  NANDN U4058 ( .A(n3394), .B(n3393), .Z(n3395) );
  NAND U4059 ( .A(n3396), .B(n3395), .Z(n3422) );
  XNOR U4060 ( .A(n3423), .B(n3422), .Z(n3408) );
  NANDN U4061 ( .A(n3398), .B(n3397), .Z(n3402) );
  OR U4062 ( .A(n3400), .B(n3399), .Z(n3401) );
  NAND U4063 ( .A(n3402), .B(n3401), .Z(n3409) );
  XNOR U4064 ( .A(n3408), .B(n3409), .Z(n3410) );
  XOR U4065 ( .A(n3411), .B(n3410), .Z(n3407) );
  XOR U4066 ( .A(sreg[1096]), .B(n3406), .Z(n3405) );
  XOR U4067 ( .A(n3407), .B(n3405), .Z(c[1096]) );
  NANDN U4068 ( .A(n3409), .B(n3408), .Z(n3413) );
  NAND U4069 ( .A(n3411), .B(n3410), .Z(n3412) );
  NAND U4070 ( .A(n3413), .B(n3412), .Z(n3434) );
  AND U4071 ( .A(b[2]), .B(a[75]), .Z(n3440) );
  AND U4072 ( .A(a[76]), .B(b[1]), .Z(n3438) );
  AND U4073 ( .A(a[74]), .B(b[3]), .Z(n3437) );
  XOR U4074 ( .A(n3438), .B(n3437), .Z(n3439) );
  XOR U4075 ( .A(n3440), .B(n3439), .Z(n3443) );
  NAND U4076 ( .A(b[0]), .B(a[77]), .Z(n3444) );
  XOR U4077 ( .A(n3443), .B(n3444), .Z(n3446) );
  OR U4078 ( .A(n3415), .B(n3414), .Z(n3419) );
  NANDN U4079 ( .A(n3417), .B(n3416), .Z(n3418) );
  NAND U4080 ( .A(n3419), .B(n3418), .Z(n3445) );
  XNOR U4081 ( .A(n3446), .B(n3445), .Z(n3431) );
  NANDN U4082 ( .A(n3421), .B(n3420), .Z(n3425) );
  OR U4083 ( .A(n3423), .B(n3422), .Z(n3424) );
  NAND U4084 ( .A(n3425), .B(n3424), .Z(n3432) );
  XNOR U4085 ( .A(n3431), .B(n3432), .Z(n3433) );
  XNOR U4086 ( .A(n3434), .B(n3433), .Z(n3426) );
  XNOR U4087 ( .A(n3426), .B(sreg[1097]), .Z(n3427) );
  XOR U4088 ( .A(n3428), .B(n3427), .Z(c[1097]) );
  NAND U4089 ( .A(n3426), .B(sreg[1097]), .Z(n3430) );
  OR U4090 ( .A(n3428), .B(n3427), .Z(n3429) );
  AND U4091 ( .A(n3430), .B(n3429), .Z(n3469) );
  NANDN U4092 ( .A(n3432), .B(n3431), .Z(n3436) );
  NAND U4093 ( .A(n3434), .B(n3433), .Z(n3435) );
  NAND U4094 ( .A(n3436), .B(n3435), .Z(n3453) );
  AND U4095 ( .A(b[2]), .B(a[76]), .Z(n3459) );
  AND U4096 ( .A(a[77]), .B(b[1]), .Z(n3457) );
  AND U4097 ( .A(a[75]), .B(b[3]), .Z(n3456) );
  XOR U4098 ( .A(n3457), .B(n3456), .Z(n3458) );
  XOR U4099 ( .A(n3459), .B(n3458), .Z(n3462) );
  NAND U4100 ( .A(b[0]), .B(a[78]), .Z(n3463) );
  XOR U4101 ( .A(n3462), .B(n3463), .Z(n3465) );
  OR U4102 ( .A(n3438), .B(n3437), .Z(n3442) );
  NANDN U4103 ( .A(n3440), .B(n3439), .Z(n3441) );
  NAND U4104 ( .A(n3442), .B(n3441), .Z(n3464) );
  XNOR U4105 ( .A(n3465), .B(n3464), .Z(n3450) );
  NANDN U4106 ( .A(n3444), .B(n3443), .Z(n3448) );
  OR U4107 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U4108 ( .A(n3448), .B(n3447), .Z(n3451) );
  XNOR U4109 ( .A(n3450), .B(n3451), .Z(n3452) );
  XNOR U4110 ( .A(n3453), .B(n3452), .Z(n3468) );
  XNOR U4111 ( .A(sreg[1098]), .B(n3468), .Z(n3449) );
  XOR U4112 ( .A(n3469), .B(n3449), .Z(c[1098]) );
  NANDN U4113 ( .A(n3451), .B(n3450), .Z(n3455) );
  NAND U4114 ( .A(n3453), .B(n3452), .Z(n3454) );
  NAND U4115 ( .A(n3455), .B(n3454), .Z(n3474) );
  AND U4116 ( .A(b[2]), .B(a[77]), .Z(n3480) );
  AND U4117 ( .A(a[78]), .B(b[1]), .Z(n3478) );
  AND U4118 ( .A(a[76]), .B(b[3]), .Z(n3477) );
  XOR U4119 ( .A(n3478), .B(n3477), .Z(n3479) );
  XOR U4120 ( .A(n3480), .B(n3479), .Z(n3483) );
  NAND U4121 ( .A(b[0]), .B(a[79]), .Z(n3484) );
  XOR U4122 ( .A(n3483), .B(n3484), .Z(n3486) );
  OR U4123 ( .A(n3457), .B(n3456), .Z(n3461) );
  NANDN U4124 ( .A(n3459), .B(n3458), .Z(n3460) );
  NAND U4125 ( .A(n3461), .B(n3460), .Z(n3485) );
  XNOR U4126 ( .A(n3486), .B(n3485), .Z(n3471) );
  NANDN U4127 ( .A(n3463), .B(n3462), .Z(n3467) );
  OR U4128 ( .A(n3465), .B(n3464), .Z(n3466) );
  NAND U4129 ( .A(n3467), .B(n3466), .Z(n3472) );
  XNOR U4130 ( .A(n3471), .B(n3472), .Z(n3473) );
  XOR U4131 ( .A(n3474), .B(n3473), .Z(n3490) );
  XNOR U4132 ( .A(sreg[1099]), .B(n3489), .Z(n3470) );
  XOR U4133 ( .A(n3490), .B(n3470), .Z(c[1099]) );
  NANDN U4134 ( .A(n3472), .B(n3471), .Z(n3476) );
  NAND U4135 ( .A(n3474), .B(n3473), .Z(n3475) );
  NAND U4136 ( .A(n3476), .B(n3475), .Z(n3495) );
  AND U4137 ( .A(b[2]), .B(a[78]), .Z(n3501) );
  AND U4138 ( .A(a[79]), .B(b[1]), .Z(n3499) );
  AND U4139 ( .A(a[77]), .B(b[3]), .Z(n3498) );
  XOR U4140 ( .A(n3499), .B(n3498), .Z(n3500) );
  XOR U4141 ( .A(n3501), .B(n3500), .Z(n3504) );
  NAND U4142 ( .A(b[0]), .B(a[80]), .Z(n3505) );
  XOR U4143 ( .A(n3504), .B(n3505), .Z(n3507) );
  OR U4144 ( .A(n3478), .B(n3477), .Z(n3482) );
  NANDN U4145 ( .A(n3480), .B(n3479), .Z(n3481) );
  NAND U4146 ( .A(n3482), .B(n3481), .Z(n3506) );
  XNOR U4147 ( .A(n3507), .B(n3506), .Z(n3492) );
  NANDN U4148 ( .A(n3484), .B(n3483), .Z(n3488) );
  OR U4149 ( .A(n3486), .B(n3485), .Z(n3487) );
  NAND U4150 ( .A(n3488), .B(n3487), .Z(n3493) );
  XNOR U4151 ( .A(n3492), .B(n3493), .Z(n3494) );
  XOR U4152 ( .A(n3495), .B(n3494), .Z(n3511) );
  XNOR U4153 ( .A(sreg[1100]), .B(n3510), .Z(n3491) );
  XOR U4154 ( .A(n3511), .B(n3491), .Z(c[1100]) );
  NANDN U4155 ( .A(n3493), .B(n3492), .Z(n3497) );
  NAND U4156 ( .A(n3495), .B(n3494), .Z(n3496) );
  NAND U4157 ( .A(n3497), .B(n3496), .Z(n3516) );
  AND U4158 ( .A(b[2]), .B(a[79]), .Z(n3522) );
  AND U4159 ( .A(a[80]), .B(b[1]), .Z(n3520) );
  AND U4160 ( .A(a[78]), .B(b[3]), .Z(n3519) );
  XOR U4161 ( .A(n3520), .B(n3519), .Z(n3521) );
  XOR U4162 ( .A(n3522), .B(n3521), .Z(n3525) );
  NAND U4163 ( .A(b[0]), .B(a[81]), .Z(n3526) );
  XOR U4164 ( .A(n3525), .B(n3526), .Z(n3528) );
  OR U4165 ( .A(n3499), .B(n3498), .Z(n3503) );
  NANDN U4166 ( .A(n3501), .B(n3500), .Z(n3502) );
  NAND U4167 ( .A(n3503), .B(n3502), .Z(n3527) );
  XNOR U4168 ( .A(n3528), .B(n3527), .Z(n3513) );
  NANDN U4169 ( .A(n3505), .B(n3504), .Z(n3509) );
  OR U4170 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U4171 ( .A(n3509), .B(n3508), .Z(n3514) );
  XNOR U4172 ( .A(n3513), .B(n3514), .Z(n3515) );
  XNOR U4173 ( .A(n3516), .B(n3515), .Z(n3532) );
  XOR U4174 ( .A(n3531), .B(sreg[1101]), .Z(n3512) );
  XOR U4175 ( .A(n3532), .B(n3512), .Z(c[1101]) );
  NANDN U4176 ( .A(n3514), .B(n3513), .Z(n3518) );
  NAND U4177 ( .A(n3516), .B(n3515), .Z(n3517) );
  NAND U4178 ( .A(n3518), .B(n3517), .Z(n3539) );
  AND U4179 ( .A(b[2]), .B(a[80]), .Z(n3545) );
  AND U4180 ( .A(a[81]), .B(b[1]), .Z(n3543) );
  AND U4181 ( .A(a[79]), .B(b[3]), .Z(n3542) );
  XOR U4182 ( .A(n3543), .B(n3542), .Z(n3544) );
  XOR U4183 ( .A(n3545), .B(n3544), .Z(n3548) );
  NAND U4184 ( .A(b[0]), .B(a[82]), .Z(n3549) );
  XOR U4185 ( .A(n3548), .B(n3549), .Z(n3551) );
  OR U4186 ( .A(n3520), .B(n3519), .Z(n3524) );
  NANDN U4187 ( .A(n3522), .B(n3521), .Z(n3523) );
  NAND U4188 ( .A(n3524), .B(n3523), .Z(n3550) );
  XNOR U4189 ( .A(n3551), .B(n3550), .Z(n3536) );
  NANDN U4190 ( .A(n3526), .B(n3525), .Z(n3530) );
  OR U4191 ( .A(n3528), .B(n3527), .Z(n3529) );
  NAND U4192 ( .A(n3530), .B(n3529), .Z(n3537) );
  XNOR U4193 ( .A(n3536), .B(n3537), .Z(n3538) );
  XOR U4194 ( .A(n3539), .B(n3538), .Z(n3535) );
  XOR U4195 ( .A(sreg[1102]), .B(n3534), .Z(n3533) );
  XOR U4196 ( .A(n3535), .B(n3533), .Z(c[1102]) );
  NANDN U4197 ( .A(n3537), .B(n3536), .Z(n3541) );
  NAND U4198 ( .A(n3539), .B(n3538), .Z(n3540) );
  NAND U4199 ( .A(n3541), .B(n3540), .Z(n3557) );
  AND U4200 ( .A(b[2]), .B(a[81]), .Z(n3563) );
  AND U4201 ( .A(a[82]), .B(b[1]), .Z(n3561) );
  AND U4202 ( .A(a[80]), .B(b[3]), .Z(n3560) );
  XOR U4203 ( .A(n3561), .B(n3560), .Z(n3562) );
  XOR U4204 ( .A(n3563), .B(n3562), .Z(n3566) );
  NAND U4205 ( .A(b[0]), .B(a[83]), .Z(n3567) );
  XOR U4206 ( .A(n3566), .B(n3567), .Z(n3569) );
  OR U4207 ( .A(n3543), .B(n3542), .Z(n3547) );
  NANDN U4208 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U4209 ( .A(n3547), .B(n3546), .Z(n3568) );
  XNOR U4210 ( .A(n3569), .B(n3568), .Z(n3554) );
  NANDN U4211 ( .A(n3549), .B(n3548), .Z(n3553) );
  OR U4212 ( .A(n3551), .B(n3550), .Z(n3552) );
  NAND U4213 ( .A(n3553), .B(n3552), .Z(n3555) );
  XNOR U4214 ( .A(n3554), .B(n3555), .Z(n3556) );
  XNOR U4215 ( .A(n3557), .B(n3556), .Z(n3572) );
  XNOR U4216 ( .A(n3572), .B(sreg[1103]), .Z(n3573) );
  XOR U4217 ( .A(n3574), .B(n3573), .Z(c[1103]) );
  NANDN U4218 ( .A(n3555), .B(n3554), .Z(n3559) );
  NAND U4219 ( .A(n3557), .B(n3556), .Z(n3558) );
  NAND U4220 ( .A(n3559), .B(n3558), .Z(n3583) );
  AND U4221 ( .A(b[2]), .B(a[82]), .Z(n3595) );
  AND U4222 ( .A(a[83]), .B(b[1]), .Z(n3593) );
  AND U4223 ( .A(a[81]), .B(b[3]), .Z(n3592) );
  XOR U4224 ( .A(n3593), .B(n3592), .Z(n3594) );
  XOR U4225 ( .A(n3595), .B(n3594), .Z(n3586) );
  NAND U4226 ( .A(b[0]), .B(a[84]), .Z(n3587) );
  XOR U4227 ( .A(n3586), .B(n3587), .Z(n3589) );
  OR U4228 ( .A(n3561), .B(n3560), .Z(n3565) );
  NANDN U4229 ( .A(n3563), .B(n3562), .Z(n3564) );
  NAND U4230 ( .A(n3565), .B(n3564), .Z(n3588) );
  XNOR U4231 ( .A(n3589), .B(n3588), .Z(n3580) );
  NANDN U4232 ( .A(n3567), .B(n3566), .Z(n3571) );
  OR U4233 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U4234 ( .A(n3571), .B(n3570), .Z(n3581) );
  XNOR U4235 ( .A(n3580), .B(n3581), .Z(n3582) );
  XNOR U4236 ( .A(n3583), .B(n3582), .Z(n3579) );
  NAND U4237 ( .A(n3572), .B(sreg[1103]), .Z(n3576) );
  OR U4238 ( .A(n3574), .B(n3573), .Z(n3575) );
  AND U4239 ( .A(n3576), .B(n3575), .Z(n3578) );
  XNOR U4240 ( .A(n3578), .B(sreg[1104]), .Z(n3577) );
  XOR U4241 ( .A(n3579), .B(n3577), .Z(c[1104]) );
  NANDN U4242 ( .A(n3581), .B(n3580), .Z(n3585) );
  NAND U4243 ( .A(n3583), .B(n3582), .Z(n3584) );
  NAND U4244 ( .A(n3585), .B(n3584), .Z(n3613) );
  NANDN U4245 ( .A(n3587), .B(n3586), .Z(n3591) );
  OR U4246 ( .A(n3589), .B(n3588), .Z(n3590) );
  NAND U4247 ( .A(n3591), .B(n3590), .Z(n3610) );
  AND U4248 ( .A(b[2]), .B(a[83]), .Z(n3601) );
  AND U4249 ( .A(a[84]), .B(b[1]), .Z(n3599) );
  AND U4250 ( .A(a[82]), .B(b[3]), .Z(n3598) );
  XOR U4251 ( .A(n3599), .B(n3598), .Z(n3600) );
  XOR U4252 ( .A(n3601), .B(n3600), .Z(n3604) );
  NAND U4253 ( .A(b[0]), .B(a[85]), .Z(n3605) );
  XNOR U4254 ( .A(n3604), .B(n3605), .Z(n3606) );
  OR U4255 ( .A(n3593), .B(n3592), .Z(n3597) );
  NANDN U4256 ( .A(n3595), .B(n3594), .Z(n3596) );
  AND U4257 ( .A(n3597), .B(n3596), .Z(n3607) );
  XNOR U4258 ( .A(n3606), .B(n3607), .Z(n3611) );
  XNOR U4259 ( .A(n3610), .B(n3611), .Z(n3612) );
  XNOR U4260 ( .A(n3613), .B(n3612), .Z(n3616) );
  XNOR U4261 ( .A(sreg[1105]), .B(n3616), .Z(n3618) );
  XNOR U4262 ( .A(n3617), .B(n3618), .Z(c[1105]) );
  AND U4263 ( .A(b[2]), .B(a[84]), .Z(n3631) );
  AND U4264 ( .A(a[85]), .B(b[1]), .Z(n3629) );
  AND U4265 ( .A(a[83]), .B(b[3]), .Z(n3628) );
  XOR U4266 ( .A(n3629), .B(n3628), .Z(n3630) );
  XOR U4267 ( .A(n3631), .B(n3630), .Z(n3634) );
  NAND U4268 ( .A(b[0]), .B(a[86]), .Z(n3635) );
  XOR U4269 ( .A(n3634), .B(n3635), .Z(n3637) );
  OR U4270 ( .A(n3599), .B(n3598), .Z(n3603) );
  NANDN U4271 ( .A(n3601), .B(n3600), .Z(n3602) );
  NAND U4272 ( .A(n3603), .B(n3602), .Z(n3636) );
  XNOR U4273 ( .A(n3637), .B(n3636), .Z(n3622) );
  NANDN U4274 ( .A(n3605), .B(n3604), .Z(n3609) );
  NAND U4275 ( .A(n3607), .B(n3606), .Z(n3608) );
  NAND U4276 ( .A(n3609), .B(n3608), .Z(n3623) );
  XNOR U4277 ( .A(n3622), .B(n3623), .Z(n3624) );
  NANDN U4278 ( .A(n3611), .B(n3610), .Z(n3615) );
  NANDN U4279 ( .A(n3613), .B(n3612), .Z(n3614) );
  NAND U4280 ( .A(n3615), .B(n3614), .Z(n3625) );
  XOR U4281 ( .A(n3624), .B(n3625), .Z(n3641) );
  NAND U4282 ( .A(sreg[1105]), .B(n3616), .Z(n3620) );
  NANDN U4283 ( .A(n3618), .B(n3617), .Z(n3619) );
  NAND U4284 ( .A(n3620), .B(n3619), .Z(n3640) );
  XNOR U4285 ( .A(sreg[1106]), .B(n3640), .Z(n3621) );
  XNOR U4286 ( .A(n3641), .B(n3621), .Z(c[1106]) );
  NANDN U4287 ( .A(n3623), .B(n3622), .Z(n3627) );
  NANDN U4288 ( .A(n3625), .B(n3624), .Z(n3626) );
  NAND U4289 ( .A(n3627), .B(n3626), .Z(n3658) );
  AND U4290 ( .A(b[2]), .B(a[85]), .Z(n3652) );
  AND U4291 ( .A(a[86]), .B(b[1]), .Z(n3650) );
  AND U4292 ( .A(a[84]), .B(b[3]), .Z(n3649) );
  XOR U4293 ( .A(n3650), .B(n3649), .Z(n3651) );
  XOR U4294 ( .A(n3652), .B(n3651), .Z(n3643) );
  NAND U4295 ( .A(b[0]), .B(a[87]), .Z(n3644) );
  XOR U4296 ( .A(n3643), .B(n3644), .Z(n3646) );
  OR U4297 ( .A(n3629), .B(n3628), .Z(n3633) );
  NANDN U4298 ( .A(n3631), .B(n3630), .Z(n3632) );
  NAND U4299 ( .A(n3633), .B(n3632), .Z(n3645) );
  XNOR U4300 ( .A(n3646), .B(n3645), .Z(n3655) );
  NANDN U4301 ( .A(n3635), .B(n3634), .Z(n3639) );
  OR U4302 ( .A(n3637), .B(n3636), .Z(n3638) );
  NAND U4303 ( .A(n3639), .B(n3638), .Z(n3656) );
  XNOR U4304 ( .A(n3655), .B(n3656), .Z(n3657) );
  XOR U4305 ( .A(n3658), .B(n3657), .Z(n3662) );
  XNOR U4306 ( .A(sreg[1107]), .B(n3661), .Z(n3642) );
  XOR U4307 ( .A(n3662), .B(n3642), .Z(c[1107]) );
  NANDN U4308 ( .A(n3644), .B(n3643), .Z(n3648) );
  OR U4309 ( .A(n3646), .B(n3645), .Z(n3647) );
  NAND U4310 ( .A(n3648), .B(n3647), .Z(n3664) );
  AND U4311 ( .A(b[2]), .B(a[86]), .Z(n3673) );
  AND U4312 ( .A(a[87]), .B(b[1]), .Z(n3671) );
  AND U4313 ( .A(a[85]), .B(b[3]), .Z(n3670) );
  XOR U4314 ( .A(n3671), .B(n3670), .Z(n3672) );
  XOR U4315 ( .A(n3673), .B(n3672), .Z(n3676) );
  NAND U4316 ( .A(b[0]), .B(a[88]), .Z(n3677) );
  XNOR U4317 ( .A(n3676), .B(n3677), .Z(n3678) );
  OR U4318 ( .A(n3650), .B(n3649), .Z(n3654) );
  NANDN U4319 ( .A(n3652), .B(n3651), .Z(n3653) );
  AND U4320 ( .A(n3654), .B(n3653), .Z(n3679) );
  XNOR U4321 ( .A(n3678), .B(n3679), .Z(n3665) );
  XNOR U4322 ( .A(n3664), .B(n3665), .Z(n3666) );
  NANDN U4323 ( .A(n3656), .B(n3655), .Z(n3660) );
  NAND U4324 ( .A(n3658), .B(n3657), .Z(n3659) );
  AND U4325 ( .A(n3660), .B(n3659), .Z(n3667) );
  XNOR U4326 ( .A(n3666), .B(n3667), .Z(n3683) );
  XNOR U4327 ( .A(sreg[1108]), .B(n3682), .Z(n3663) );
  XOR U4328 ( .A(n3683), .B(n3663), .Z(c[1108]) );
  NANDN U4329 ( .A(n3665), .B(n3664), .Z(n3669) );
  NAND U4330 ( .A(n3667), .B(n3666), .Z(n3668) );
  NAND U4331 ( .A(n3669), .B(n3668), .Z(n3690) );
  AND U4332 ( .A(b[2]), .B(a[87]), .Z(n3696) );
  AND U4333 ( .A(a[88]), .B(b[1]), .Z(n3694) );
  AND U4334 ( .A(a[86]), .B(b[3]), .Z(n3693) );
  XOR U4335 ( .A(n3694), .B(n3693), .Z(n3695) );
  XOR U4336 ( .A(n3696), .B(n3695), .Z(n3699) );
  NAND U4337 ( .A(b[0]), .B(a[89]), .Z(n3700) );
  XOR U4338 ( .A(n3699), .B(n3700), .Z(n3702) );
  OR U4339 ( .A(n3671), .B(n3670), .Z(n3675) );
  NANDN U4340 ( .A(n3673), .B(n3672), .Z(n3674) );
  NAND U4341 ( .A(n3675), .B(n3674), .Z(n3701) );
  XNOR U4342 ( .A(n3702), .B(n3701), .Z(n3687) );
  NANDN U4343 ( .A(n3677), .B(n3676), .Z(n3681) );
  NAND U4344 ( .A(n3679), .B(n3678), .Z(n3680) );
  NAND U4345 ( .A(n3681), .B(n3680), .Z(n3688) );
  XNOR U4346 ( .A(n3687), .B(n3688), .Z(n3689) );
  XNOR U4347 ( .A(n3690), .B(n3689), .Z(n3686) );
  XOR U4348 ( .A(n3685), .B(sreg[1109]), .Z(n3684) );
  XNOR U4349 ( .A(n3686), .B(n3684), .Z(c[1109]) );
  NANDN U4350 ( .A(n3688), .B(n3687), .Z(n3692) );
  NANDN U4351 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U4352 ( .A(n3692), .B(n3691), .Z(n3720) );
  AND U4353 ( .A(b[2]), .B(a[88]), .Z(n3714) );
  AND U4354 ( .A(a[89]), .B(b[1]), .Z(n3712) );
  AND U4355 ( .A(a[87]), .B(b[3]), .Z(n3711) );
  XOR U4356 ( .A(n3712), .B(n3711), .Z(n3713) );
  XOR U4357 ( .A(n3714), .B(n3713), .Z(n3705) );
  NAND U4358 ( .A(b[0]), .B(a[90]), .Z(n3706) );
  XOR U4359 ( .A(n3705), .B(n3706), .Z(n3708) );
  OR U4360 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U4361 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U4362 ( .A(n3698), .B(n3697), .Z(n3707) );
  XNOR U4363 ( .A(n3708), .B(n3707), .Z(n3717) );
  NANDN U4364 ( .A(n3700), .B(n3699), .Z(n3704) );
  OR U4365 ( .A(n3702), .B(n3701), .Z(n3703) );
  NAND U4366 ( .A(n3704), .B(n3703), .Z(n3718) );
  XNOR U4367 ( .A(n3717), .B(n3718), .Z(n3719) );
  XNOR U4368 ( .A(n3720), .B(n3719), .Z(n3723) );
  XNOR U4369 ( .A(n3723), .B(sreg[1110]), .Z(n3725) );
  XNOR U4370 ( .A(n3724), .B(n3725), .Z(c[1110]) );
  NANDN U4371 ( .A(n3706), .B(n3705), .Z(n3710) );
  OR U4372 ( .A(n3708), .B(n3707), .Z(n3709) );
  NAND U4373 ( .A(n3710), .B(n3709), .Z(n3728) );
  AND U4374 ( .A(b[2]), .B(a[89]), .Z(n3737) );
  AND U4375 ( .A(a[90]), .B(b[1]), .Z(n3735) );
  AND U4376 ( .A(a[88]), .B(b[3]), .Z(n3734) );
  XOR U4377 ( .A(n3735), .B(n3734), .Z(n3736) );
  XOR U4378 ( .A(n3737), .B(n3736), .Z(n3740) );
  NAND U4379 ( .A(b[0]), .B(a[91]), .Z(n3741) );
  XNOR U4380 ( .A(n3740), .B(n3741), .Z(n3742) );
  OR U4381 ( .A(n3712), .B(n3711), .Z(n3716) );
  NANDN U4382 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U4383 ( .A(n3716), .B(n3715), .Z(n3743) );
  XNOR U4384 ( .A(n3742), .B(n3743), .Z(n3729) );
  XNOR U4385 ( .A(n3728), .B(n3729), .Z(n3730) );
  NANDN U4386 ( .A(n3718), .B(n3717), .Z(n3722) );
  NAND U4387 ( .A(n3720), .B(n3719), .Z(n3721) );
  NAND U4388 ( .A(n3722), .B(n3721), .Z(n3731) );
  XNOR U4389 ( .A(n3730), .B(n3731), .Z(n3746) );
  XOR U4390 ( .A(sreg[1111]), .B(n3746), .Z(n3747) );
  NAND U4391 ( .A(n3723), .B(sreg[1110]), .Z(n3727) );
  NANDN U4392 ( .A(n3725), .B(n3724), .Z(n3726) );
  NAND U4393 ( .A(n3727), .B(n3726), .Z(n3748) );
  XOR U4394 ( .A(n3747), .B(n3748), .Z(c[1111]) );
  NANDN U4395 ( .A(n3729), .B(n3728), .Z(n3733) );
  NANDN U4396 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U4397 ( .A(n3733), .B(n3732), .Z(n3757) );
  AND U4398 ( .A(b[2]), .B(a[90]), .Z(n3763) );
  AND U4399 ( .A(a[91]), .B(b[1]), .Z(n3761) );
  AND U4400 ( .A(a[89]), .B(b[3]), .Z(n3760) );
  XOR U4401 ( .A(n3761), .B(n3760), .Z(n3762) );
  XOR U4402 ( .A(n3763), .B(n3762), .Z(n3766) );
  NAND U4403 ( .A(b[0]), .B(a[92]), .Z(n3767) );
  XOR U4404 ( .A(n3766), .B(n3767), .Z(n3769) );
  OR U4405 ( .A(n3735), .B(n3734), .Z(n3739) );
  NANDN U4406 ( .A(n3737), .B(n3736), .Z(n3738) );
  NAND U4407 ( .A(n3739), .B(n3738), .Z(n3768) );
  XNOR U4408 ( .A(n3769), .B(n3768), .Z(n3754) );
  NANDN U4409 ( .A(n3741), .B(n3740), .Z(n3745) );
  NAND U4410 ( .A(n3743), .B(n3742), .Z(n3744) );
  NAND U4411 ( .A(n3745), .B(n3744), .Z(n3755) );
  XNOR U4412 ( .A(n3754), .B(n3755), .Z(n3756) );
  XOR U4413 ( .A(n3757), .B(n3756), .Z(n3753) );
  OR U4414 ( .A(n3746), .B(sreg[1111]), .Z(n3750) );
  NANDN U4415 ( .A(n3748), .B(n3747), .Z(n3749) );
  AND U4416 ( .A(n3750), .B(n3749), .Z(n3752) );
  XNOR U4417 ( .A(sreg[1112]), .B(n3752), .Z(n3751) );
  XNOR U4418 ( .A(n3753), .B(n3751), .Z(c[1112]) );
  NANDN U4419 ( .A(n3755), .B(n3754), .Z(n3759) );
  NANDN U4420 ( .A(n3757), .B(n3756), .Z(n3758) );
  NAND U4421 ( .A(n3759), .B(n3758), .Z(n3787) );
  AND U4422 ( .A(b[2]), .B(a[91]), .Z(n3781) );
  AND U4423 ( .A(a[92]), .B(b[1]), .Z(n3779) );
  AND U4424 ( .A(a[90]), .B(b[3]), .Z(n3778) );
  XOR U4425 ( .A(n3779), .B(n3778), .Z(n3780) );
  XOR U4426 ( .A(n3781), .B(n3780), .Z(n3772) );
  NAND U4427 ( .A(b[0]), .B(a[93]), .Z(n3773) );
  XOR U4428 ( .A(n3772), .B(n3773), .Z(n3775) );
  OR U4429 ( .A(n3761), .B(n3760), .Z(n3765) );
  NANDN U4430 ( .A(n3763), .B(n3762), .Z(n3764) );
  NAND U4431 ( .A(n3765), .B(n3764), .Z(n3774) );
  XNOR U4432 ( .A(n3775), .B(n3774), .Z(n3784) );
  NANDN U4433 ( .A(n3767), .B(n3766), .Z(n3771) );
  OR U4434 ( .A(n3769), .B(n3768), .Z(n3770) );
  NAND U4435 ( .A(n3771), .B(n3770), .Z(n3785) );
  XNOR U4436 ( .A(n3784), .B(n3785), .Z(n3786) );
  XNOR U4437 ( .A(n3787), .B(n3786), .Z(n3790) );
  XNOR U4438 ( .A(n3790), .B(sreg[1113]), .Z(n3791) );
  XOR U4439 ( .A(n3792), .B(n3791), .Z(c[1113]) );
  NANDN U4440 ( .A(n3773), .B(n3772), .Z(n3777) );
  OR U4441 ( .A(n3775), .B(n3774), .Z(n3776) );
  NAND U4442 ( .A(n3777), .B(n3776), .Z(n3798) );
  AND U4443 ( .A(b[2]), .B(a[92]), .Z(n3807) );
  AND U4444 ( .A(a[93]), .B(b[1]), .Z(n3805) );
  AND U4445 ( .A(a[91]), .B(b[3]), .Z(n3804) );
  XOR U4446 ( .A(n3805), .B(n3804), .Z(n3806) );
  XOR U4447 ( .A(n3807), .B(n3806), .Z(n3810) );
  NAND U4448 ( .A(b[0]), .B(a[94]), .Z(n3811) );
  XNOR U4449 ( .A(n3810), .B(n3811), .Z(n3812) );
  OR U4450 ( .A(n3779), .B(n3778), .Z(n3783) );
  NANDN U4451 ( .A(n3781), .B(n3780), .Z(n3782) );
  AND U4452 ( .A(n3783), .B(n3782), .Z(n3813) );
  XNOR U4453 ( .A(n3812), .B(n3813), .Z(n3799) );
  XNOR U4454 ( .A(n3798), .B(n3799), .Z(n3800) );
  NANDN U4455 ( .A(n3785), .B(n3784), .Z(n3789) );
  NAND U4456 ( .A(n3787), .B(n3786), .Z(n3788) );
  NAND U4457 ( .A(n3789), .B(n3788), .Z(n3801) );
  XOR U4458 ( .A(n3800), .B(n3801), .Z(n3797) );
  NAND U4459 ( .A(n3790), .B(sreg[1113]), .Z(n3794) );
  OR U4460 ( .A(n3792), .B(n3791), .Z(n3793) );
  AND U4461 ( .A(n3794), .B(n3793), .Z(n3796) );
  XNOR U4462 ( .A(n3796), .B(sreg[1114]), .Z(n3795) );
  XNOR U4463 ( .A(n3797), .B(n3795), .Z(c[1114]) );
  NANDN U4464 ( .A(n3799), .B(n3798), .Z(n3803) );
  NANDN U4465 ( .A(n3801), .B(n3800), .Z(n3802) );
  NAND U4466 ( .A(n3803), .B(n3802), .Z(n3819) );
  AND U4467 ( .A(b[2]), .B(a[93]), .Z(n3825) );
  AND U4468 ( .A(a[94]), .B(b[1]), .Z(n3823) );
  AND U4469 ( .A(a[92]), .B(b[3]), .Z(n3822) );
  XOR U4470 ( .A(n3823), .B(n3822), .Z(n3824) );
  XOR U4471 ( .A(n3825), .B(n3824), .Z(n3828) );
  NAND U4472 ( .A(b[0]), .B(a[95]), .Z(n3829) );
  XOR U4473 ( .A(n3828), .B(n3829), .Z(n3831) );
  OR U4474 ( .A(n3805), .B(n3804), .Z(n3809) );
  NANDN U4475 ( .A(n3807), .B(n3806), .Z(n3808) );
  NAND U4476 ( .A(n3809), .B(n3808), .Z(n3830) );
  XNOR U4477 ( .A(n3831), .B(n3830), .Z(n3816) );
  NANDN U4478 ( .A(n3811), .B(n3810), .Z(n3815) );
  NAND U4479 ( .A(n3813), .B(n3812), .Z(n3814) );
  NAND U4480 ( .A(n3815), .B(n3814), .Z(n3817) );
  XNOR U4481 ( .A(n3816), .B(n3817), .Z(n3818) );
  XNOR U4482 ( .A(n3819), .B(n3818), .Z(n3834) );
  XOR U4483 ( .A(sreg[1115]), .B(n3834), .Z(n3836) );
  XNOR U4484 ( .A(n3835), .B(n3836), .Z(c[1115]) );
  NANDN U4485 ( .A(n3817), .B(n3816), .Z(n3821) );
  NANDN U4486 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U4487 ( .A(n3821), .B(n3820), .Z(n3854) );
  AND U4488 ( .A(b[2]), .B(a[94]), .Z(n3848) );
  AND U4489 ( .A(a[95]), .B(b[1]), .Z(n3846) );
  AND U4490 ( .A(a[93]), .B(b[3]), .Z(n3845) );
  XOR U4491 ( .A(n3846), .B(n3845), .Z(n3847) );
  XOR U4492 ( .A(n3848), .B(n3847), .Z(n3839) );
  NAND U4493 ( .A(b[0]), .B(a[96]), .Z(n3840) );
  XOR U4494 ( .A(n3839), .B(n3840), .Z(n3842) );
  OR U4495 ( .A(n3823), .B(n3822), .Z(n3827) );
  NANDN U4496 ( .A(n3825), .B(n3824), .Z(n3826) );
  NAND U4497 ( .A(n3827), .B(n3826), .Z(n3841) );
  XNOR U4498 ( .A(n3842), .B(n3841), .Z(n3851) );
  NANDN U4499 ( .A(n3829), .B(n3828), .Z(n3833) );
  OR U4500 ( .A(n3831), .B(n3830), .Z(n3832) );
  NAND U4501 ( .A(n3833), .B(n3832), .Z(n3852) );
  XNOR U4502 ( .A(n3851), .B(n3852), .Z(n3853) );
  XNOR U4503 ( .A(n3854), .B(n3853), .Z(n3857) );
  XOR U4504 ( .A(sreg[1116]), .B(n3857), .Z(n3858) );
  NANDN U4505 ( .A(n3834), .B(sreg[1115]), .Z(n3838) );
  NANDN U4506 ( .A(n3836), .B(n3835), .Z(n3837) );
  NAND U4507 ( .A(n3838), .B(n3837), .Z(n3859) );
  XOR U4508 ( .A(n3858), .B(n3859), .Z(c[1116]) );
  NANDN U4509 ( .A(n3840), .B(n3839), .Z(n3844) );
  OR U4510 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4511 ( .A(n3844), .B(n3843), .Z(n3863) );
  AND U4512 ( .A(b[2]), .B(a[95]), .Z(n3872) );
  AND U4513 ( .A(a[96]), .B(b[1]), .Z(n3870) );
  AND U4514 ( .A(a[94]), .B(b[3]), .Z(n3869) );
  XOR U4515 ( .A(n3870), .B(n3869), .Z(n3871) );
  XOR U4516 ( .A(n3872), .B(n3871), .Z(n3875) );
  NAND U4517 ( .A(b[0]), .B(a[97]), .Z(n3876) );
  XNOR U4518 ( .A(n3875), .B(n3876), .Z(n3877) );
  OR U4519 ( .A(n3846), .B(n3845), .Z(n3850) );
  NANDN U4520 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4521 ( .A(n3850), .B(n3849), .Z(n3878) );
  XNOR U4522 ( .A(n3877), .B(n3878), .Z(n3864) );
  XNOR U4523 ( .A(n3863), .B(n3864), .Z(n3865) );
  NANDN U4524 ( .A(n3852), .B(n3851), .Z(n3856) );
  NAND U4525 ( .A(n3854), .B(n3853), .Z(n3855) );
  AND U4526 ( .A(n3856), .B(n3855), .Z(n3866) );
  XNOR U4527 ( .A(n3865), .B(n3866), .Z(n3882) );
  OR U4528 ( .A(n3857), .B(sreg[1116]), .Z(n3861) );
  NANDN U4529 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U4530 ( .A(n3861), .B(n3860), .Z(n3881) );
  XNOR U4531 ( .A(sreg[1117]), .B(n3881), .Z(n3862) );
  XOR U4532 ( .A(n3882), .B(n3862), .Z(c[1117]) );
  NANDN U4533 ( .A(n3864), .B(n3863), .Z(n3868) );
  NAND U4534 ( .A(n3866), .B(n3865), .Z(n3867) );
  NAND U4535 ( .A(n3868), .B(n3867), .Z(n3887) );
  AND U4536 ( .A(b[2]), .B(a[96]), .Z(n3893) );
  AND U4537 ( .A(a[97]), .B(b[1]), .Z(n3891) );
  AND U4538 ( .A(a[95]), .B(b[3]), .Z(n3890) );
  XOR U4539 ( .A(n3891), .B(n3890), .Z(n3892) );
  XOR U4540 ( .A(n3893), .B(n3892), .Z(n3896) );
  NAND U4541 ( .A(b[0]), .B(a[98]), .Z(n3897) );
  XOR U4542 ( .A(n3896), .B(n3897), .Z(n3899) );
  OR U4543 ( .A(n3870), .B(n3869), .Z(n3874) );
  NANDN U4544 ( .A(n3872), .B(n3871), .Z(n3873) );
  NAND U4545 ( .A(n3874), .B(n3873), .Z(n3898) );
  XNOR U4546 ( .A(n3899), .B(n3898), .Z(n3884) );
  NANDN U4547 ( .A(n3876), .B(n3875), .Z(n3880) );
  NAND U4548 ( .A(n3878), .B(n3877), .Z(n3879) );
  NAND U4549 ( .A(n3880), .B(n3879), .Z(n3885) );
  XNOR U4550 ( .A(n3884), .B(n3885), .Z(n3886) );
  XOR U4551 ( .A(n3887), .B(n3886), .Z(n3903) );
  XNOR U4552 ( .A(sreg[1118]), .B(n3902), .Z(n3883) );
  XNOR U4553 ( .A(n3903), .B(n3883), .Z(c[1118]) );
  NANDN U4554 ( .A(n3885), .B(n3884), .Z(n3889) );
  NANDN U4555 ( .A(n3887), .B(n3886), .Z(n3888) );
  NAND U4556 ( .A(n3889), .B(n3888), .Z(n3908) );
  AND U4557 ( .A(b[2]), .B(a[97]), .Z(n3914) );
  AND U4558 ( .A(a[98]), .B(b[1]), .Z(n3912) );
  AND U4559 ( .A(a[96]), .B(b[3]), .Z(n3911) );
  XOR U4560 ( .A(n3912), .B(n3911), .Z(n3913) );
  XOR U4561 ( .A(n3914), .B(n3913), .Z(n3917) );
  NAND U4562 ( .A(b[0]), .B(a[99]), .Z(n3918) );
  XOR U4563 ( .A(n3917), .B(n3918), .Z(n3920) );
  OR U4564 ( .A(n3891), .B(n3890), .Z(n3895) );
  NANDN U4565 ( .A(n3893), .B(n3892), .Z(n3894) );
  NAND U4566 ( .A(n3895), .B(n3894), .Z(n3919) );
  XNOR U4567 ( .A(n3920), .B(n3919), .Z(n3905) );
  NANDN U4568 ( .A(n3897), .B(n3896), .Z(n3901) );
  OR U4569 ( .A(n3899), .B(n3898), .Z(n3900) );
  NAND U4570 ( .A(n3901), .B(n3900), .Z(n3906) );
  XNOR U4571 ( .A(n3905), .B(n3906), .Z(n3907) );
  XOR U4572 ( .A(n3908), .B(n3907), .Z(n3925) );
  XNOR U4573 ( .A(sreg[1119]), .B(n3924), .Z(n3904) );
  XOR U4574 ( .A(n3925), .B(n3904), .Z(c[1119]) );
  NANDN U4575 ( .A(n3906), .B(n3905), .Z(n3910) );
  NAND U4576 ( .A(n3908), .B(n3907), .Z(n3909) );
  AND U4577 ( .A(n3910), .B(n3909), .Z(n3931) );
  AND U4578 ( .A(b[2]), .B(a[98]), .Z(n3935) );
  AND U4579 ( .A(a[99]), .B(b[1]), .Z(n3933) );
  AND U4580 ( .A(a[97]), .B(b[3]), .Z(n3932) );
  XOR U4581 ( .A(n3933), .B(n3932), .Z(n3934) );
  XOR U4582 ( .A(n3935), .B(n3934), .Z(n3938) );
  NAND U4583 ( .A(b[0]), .B(a[100]), .Z(n3939) );
  XOR U4584 ( .A(n3938), .B(n3939), .Z(n3940) );
  OR U4585 ( .A(n3912), .B(n3911), .Z(n3916) );
  NANDN U4586 ( .A(n3914), .B(n3913), .Z(n3915) );
  AND U4587 ( .A(n3916), .B(n3915), .Z(n3941) );
  XOR U4588 ( .A(n3940), .B(n3941), .Z(n3929) );
  NANDN U4589 ( .A(n3918), .B(n3917), .Z(n3922) );
  OR U4590 ( .A(n3920), .B(n3919), .Z(n3921) );
  AND U4591 ( .A(n3922), .B(n3921), .Z(n3930) );
  XOR U4592 ( .A(n3929), .B(n3930), .Z(n3923) );
  XNOR U4593 ( .A(n3931), .B(n3923), .Z(n3928) );
  XNOR U4594 ( .A(sreg[1120]), .B(n3927), .Z(n3926) );
  XOR U4595 ( .A(n3928), .B(n3926), .Z(c[1120]) );
  AND U4596 ( .A(b[2]), .B(a[99]), .Z(n3951) );
  AND U4597 ( .A(a[100]), .B(b[1]), .Z(n3949) );
  AND U4598 ( .A(a[98]), .B(b[3]), .Z(n3948) );
  XOR U4599 ( .A(n3949), .B(n3948), .Z(n3950) );
  XOR U4600 ( .A(n3951), .B(n3950), .Z(n3954) );
  NAND U4601 ( .A(b[0]), .B(a[101]), .Z(n3955) );
  XOR U4602 ( .A(n3954), .B(n3955), .Z(n3957) );
  OR U4603 ( .A(n3933), .B(n3932), .Z(n3937) );
  NANDN U4604 ( .A(n3935), .B(n3934), .Z(n3936) );
  NAND U4605 ( .A(n3937), .B(n3936), .Z(n3956) );
  XNOR U4606 ( .A(n3957), .B(n3956), .Z(n3942) );
  XNOR U4607 ( .A(n3942), .B(n3943), .Z(n3945) );
  XOR U4608 ( .A(n3944), .B(n3945), .Z(n3960) );
  XOR U4609 ( .A(n3960), .B(sreg[1121]), .Z(n3961) );
  XOR U4610 ( .A(n3962), .B(n3961), .Z(c[1121]) );
  NANDN U4611 ( .A(n3943), .B(n3942), .Z(n3947) );
  NAND U4612 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U4613 ( .A(n3947), .B(n3946), .Z(n3971) );
  AND U4614 ( .A(b[2]), .B(a[100]), .Z(n3977) );
  AND U4615 ( .A(a[101]), .B(b[1]), .Z(n3975) );
  AND U4616 ( .A(a[99]), .B(b[3]), .Z(n3974) );
  XOR U4617 ( .A(n3975), .B(n3974), .Z(n3976) );
  XOR U4618 ( .A(n3977), .B(n3976), .Z(n3980) );
  NAND U4619 ( .A(b[0]), .B(a[102]), .Z(n3981) );
  XOR U4620 ( .A(n3980), .B(n3981), .Z(n3983) );
  OR U4621 ( .A(n3949), .B(n3948), .Z(n3953) );
  NANDN U4622 ( .A(n3951), .B(n3950), .Z(n3952) );
  NAND U4623 ( .A(n3953), .B(n3952), .Z(n3982) );
  XNOR U4624 ( .A(n3983), .B(n3982), .Z(n3968) );
  NANDN U4625 ( .A(n3955), .B(n3954), .Z(n3959) );
  OR U4626 ( .A(n3957), .B(n3956), .Z(n3958) );
  NAND U4627 ( .A(n3959), .B(n3958), .Z(n3969) );
  XNOR U4628 ( .A(n3968), .B(n3969), .Z(n3970) );
  XOR U4629 ( .A(n3971), .B(n3970), .Z(n3967) );
  NANDN U4630 ( .A(n3960), .B(sreg[1121]), .Z(n3964) );
  OR U4631 ( .A(n3962), .B(n3961), .Z(n3963) );
  NAND U4632 ( .A(n3964), .B(n3963), .Z(n3966) );
  XNOR U4633 ( .A(sreg[1122]), .B(n3966), .Z(n3965) );
  XOR U4634 ( .A(n3967), .B(n3965), .Z(c[1122]) );
  NANDN U4635 ( .A(n3969), .B(n3968), .Z(n3973) );
  NAND U4636 ( .A(n3971), .B(n3970), .Z(n3972) );
  NAND U4637 ( .A(n3973), .B(n3972), .Z(n3989) );
  AND U4638 ( .A(b[2]), .B(a[101]), .Z(n3995) );
  AND U4639 ( .A(a[102]), .B(b[1]), .Z(n3993) );
  AND U4640 ( .A(a[100]), .B(b[3]), .Z(n3992) );
  XOR U4641 ( .A(n3993), .B(n3992), .Z(n3994) );
  XOR U4642 ( .A(n3995), .B(n3994), .Z(n3998) );
  NAND U4643 ( .A(b[0]), .B(a[103]), .Z(n3999) );
  XOR U4644 ( .A(n3998), .B(n3999), .Z(n4001) );
  OR U4645 ( .A(n3975), .B(n3974), .Z(n3979) );
  NANDN U4646 ( .A(n3977), .B(n3976), .Z(n3978) );
  NAND U4647 ( .A(n3979), .B(n3978), .Z(n4000) );
  XNOR U4648 ( .A(n4001), .B(n4000), .Z(n3986) );
  NANDN U4649 ( .A(n3981), .B(n3980), .Z(n3985) );
  OR U4650 ( .A(n3983), .B(n3982), .Z(n3984) );
  NAND U4651 ( .A(n3985), .B(n3984), .Z(n3987) );
  XNOR U4652 ( .A(n3986), .B(n3987), .Z(n3988) );
  XNOR U4653 ( .A(n3989), .B(n3988), .Z(n4004) );
  XNOR U4654 ( .A(n4004), .B(sreg[1123]), .Z(n4005) );
  XOR U4655 ( .A(n4006), .B(n4005), .Z(c[1123]) );
  NANDN U4656 ( .A(n3987), .B(n3986), .Z(n3991) );
  NAND U4657 ( .A(n3989), .B(n3988), .Z(n3990) );
  NAND U4658 ( .A(n3991), .B(n3990), .Z(n4012) );
  AND U4659 ( .A(b[2]), .B(a[102]), .Z(n4018) );
  AND U4660 ( .A(a[103]), .B(b[1]), .Z(n4016) );
  AND U4661 ( .A(a[101]), .B(b[3]), .Z(n4015) );
  XOR U4662 ( .A(n4016), .B(n4015), .Z(n4017) );
  XOR U4663 ( .A(n4018), .B(n4017), .Z(n4021) );
  NAND U4664 ( .A(b[0]), .B(a[104]), .Z(n4022) );
  XOR U4665 ( .A(n4021), .B(n4022), .Z(n4024) );
  OR U4666 ( .A(n3993), .B(n3992), .Z(n3997) );
  NANDN U4667 ( .A(n3995), .B(n3994), .Z(n3996) );
  NAND U4668 ( .A(n3997), .B(n3996), .Z(n4023) );
  XNOR U4669 ( .A(n4024), .B(n4023), .Z(n4009) );
  NANDN U4670 ( .A(n3999), .B(n3998), .Z(n4003) );
  OR U4671 ( .A(n4001), .B(n4000), .Z(n4002) );
  NAND U4672 ( .A(n4003), .B(n4002), .Z(n4010) );
  XNOR U4673 ( .A(n4009), .B(n4010), .Z(n4011) );
  XNOR U4674 ( .A(n4012), .B(n4011), .Z(n4027) );
  XOR U4675 ( .A(sreg[1124]), .B(n4027), .Z(n4028) );
  NAND U4676 ( .A(n4004), .B(sreg[1123]), .Z(n4008) );
  OR U4677 ( .A(n4006), .B(n4005), .Z(n4007) );
  NAND U4678 ( .A(n4008), .B(n4007), .Z(n4029) );
  XOR U4679 ( .A(n4028), .B(n4029), .Z(c[1124]) );
  NANDN U4680 ( .A(n4010), .B(n4009), .Z(n4014) );
  NAND U4681 ( .A(n4012), .B(n4011), .Z(n4013) );
  NAND U4682 ( .A(n4014), .B(n4013), .Z(n4038) );
  AND U4683 ( .A(b[2]), .B(a[103]), .Z(n4044) );
  AND U4684 ( .A(a[104]), .B(b[1]), .Z(n4042) );
  AND U4685 ( .A(a[102]), .B(b[3]), .Z(n4041) );
  XOR U4686 ( .A(n4042), .B(n4041), .Z(n4043) );
  XOR U4687 ( .A(n4044), .B(n4043), .Z(n4047) );
  NAND U4688 ( .A(b[0]), .B(a[105]), .Z(n4048) );
  XOR U4689 ( .A(n4047), .B(n4048), .Z(n4050) );
  OR U4690 ( .A(n4016), .B(n4015), .Z(n4020) );
  NANDN U4691 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U4692 ( .A(n4020), .B(n4019), .Z(n4049) );
  XNOR U4693 ( .A(n4050), .B(n4049), .Z(n4035) );
  NANDN U4694 ( .A(n4022), .B(n4021), .Z(n4026) );
  OR U4695 ( .A(n4024), .B(n4023), .Z(n4025) );
  NAND U4696 ( .A(n4026), .B(n4025), .Z(n4036) );
  XNOR U4697 ( .A(n4035), .B(n4036), .Z(n4037) );
  XOR U4698 ( .A(n4038), .B(n4037), .Z(n4034) );
  OR U4699 ( .A(n4027), .B(sreg[1124]), .Z(n4031) );
  NANDN U4700 ( .A(n4029), .B(n4028), .Z(n4030) );
  AND U4701 ( .A(n4031), .B(n4030), .Z(n4033) );
  XNOR U4702 ( .A(sreg[1125]), .B(n4033), .Z(n4032) );
  XOR U4703 ( .A(n4034), .B(n4032), .Z(c[1125]) );
  NANDN U4704 ( .A(n4036), .B(n4035), .Z(n4040) );
  NAND U4705 ( .A(n4038), .B(n4037), .Z(n4039) );
  NAND U4706 ( .A(n4040), .B(n4039), .Z(n4056) );
  AND U4707 ( .A(b[2]), .B(a[104]), .Z(n4062) );
  AND U4708 ( .A(a[105]), .B(b[1]), .Z(n4060) );
  AND U4709 ( .A(a[103]), .B(b[3]), .Z(n4059) );
  XOR U4710 ( .A(n4060), .B(n4059), .Z(n4061) );
  XOR U4711 ( .A(n4062), .B(n4061), .Z(n4065) );
  NAND U4712 ( .A(b[0]), .B(a[106]), .Z(n4066) );
  XOR U4713 ( .A(n4065), .B(n4066), .Z(n4068) );
  OR U4714 ( .A(n4042), .B(n4041), .Z(n4046) );
  NANDN U4715 ( .A(n4044), .B(n4043), .Z(n4045) );
  NAND U4716 ( .A(n4046), .B(n4045), .Z(n4067) );
  XNOR U4717 ( .A(n4068), .B(n4067), .Z(n4053) );
  NANDN U4718 ( .A(n4048), .B(n4047), .Z(n4052) );
  OR U4719 ( .A(n4050), .B(n4049), .Z(n4051) );
  NAND U4720 ( .A(n4052), .B(n4051), .Z(n4054) );
  XNOR U4721 ( .A(n4053), .B(n4054), .Z(n4055) );
  XNOR U4722 ( .A(n4056), .B(n4055), .Z(n4071) );
  XNOR U4723 ( .A(n4071), .B(sreg[1126]), .Z(n4072) );
  XOR U4724 ( .A(n4073), .B(n4072), .Z(c[1126]) );
  NANDN U4725 ( .A(n4054), .B(n4053), .Z(n4058) );
  NAND U4726 ( .A(n4056), .B(n4055), .Z(n4057) );
  NAND U4727 ( .A(n4058), .B(n4057), .Z(n4082) );
  AND U4728 ( .A(b[2]), .B(a[105]), .Z(n4088) );
  AND U4729 ( .A(a[106]), .B(b[1]), .Z(n4086) );
  AND U4730 ( .A(a[104]), .B(b[3]), .Z(n4085) );
  XOR U4731 ( .A(n4086), .B(n4085), .Z(n4087) );
  XOR U4732 ( .A(n4088), .B(n4087), .Z(n4091) );
  NAND U4733 ( .A(b[0]), .B(a[107]), .Z(n4092) );
  XOR U4734 ( .A(n4091), .B(n4092), .Z(n4094) );
  OR U4735 ( .A(n4060), .B(n4059), .Z(n4064) );
  NANDN U4736 ( .A(n4062), .B(n4061), .Z(n4063) );
  NAND U4737 ( .A(n4064), .B(n4063), .Z(n4093) );
  XNOR U4738 ( .A(n4094), .B(n4093), .Z(n4079) );
  NANDN U4739 ( .A(n4066), .B(n4065), .Z(n4070) );
  OR U4740 ( .A(n4068), .B(n4067), .Z(n4069) );
  NAND U4741 ( .A(n4070), .B(n4069), .Z(n4080) );
  XNOR U4742 ( .A(n4079), .B(n4080), .Z(n4081) );
  XOR U4743 ( .A(n4082), .B(n4081), .Z(n4078) );
  NAND U4744 ( .A(n4071), .B(sreg[1126]), .Z(n4075) );
  OR U4745 ( .A(n4073), .B(n4072), .Z(n4074) );
  NAND U4746 ( .A(n4075), .B(n4074), .Z(n4077) );
  XNOR U4747 ( .A(sreg[1127]), .B(n4077), .Z(n4076) );
  XOR U4748 ( .A(n4078), .B(n4076), .Z(c[1127]) );
  NANDN U4749 ( .A(n4080), .B(n4079), .Z(n4084) );
  NAND U4750 ( .A(n4082), .B(n4081), .Z(n4083) );
  NAND U4751 ( .A(n4084), .B(n4083), .Z(n4100) );
  AND U4752 ( .A(b[2]), .B(a[106]), .Z(n4106) );
  AND U4753 ( .A(a[107]), .B(b[1]), .Z(n4104) );
  AND U4754 ( .A(a[105]), .B(b[3]), .Z(n4103) );
  XOR U4755 ( .A(n4104), .B(n4103), .Z(n4105) );
  XOR U4756 ( .A(n4106), .B(n4105), .Z(n4109) );
  NAND U4757 ( .A(b[0]), .B(a[108]), .Z(n4110) );
  XOR U4758 ( .A(n4109), .B(n4110), .Z(n4112) );
  OR U4759 ( .A(n4086), .B(n4085), .Z(n4090) );
  NANDN U4760 ( .A(n4088), .B(n4087), .Z(n4089) );
  NAND U4761 ( .A(n4090), .B(n4089), .Z(n4111) );
  XNOR U4762 ( .A(n4112), .B(n4111), .Z(n4097) );
  NANDN U4763 ( .A(n4092), .B(n4091), .Z(n4096) );
  OR U4764 ( .A(n4094), .B(n4093), .Z(n4095) );
  NAND U4765 ( .A(n4096), .B(n4095), .Z(n4098) );
  XNOR U4766 ( .A(n4097), .B(n4098), .Z(n4099) );
  XNOR U4767 ( .A(n4100), .B(n4099), .Z(n4115) );
  XNOR U4768 ( .A(n4115), .B(sreg[1128]), .Z(n4116) );
  XOR U4769 ( .A(n4117), .B(n4116), .Z(c[1128]) );
  NANDN U4770 ( .A(n4098), .B(n4097), .Z(n4102) );
  NAND U4771 ( .A(n4100), .B(n4099), .Z(n4101) );
  NAND U4772 ( .A(n4102), .B(n4101), .Z(n4124) );
  AND U4773 ( .A(b[2]), .B(a[107]), .Z(n4130) );
  AND U4774 ( .A(a[108]), .B(b[1]), .Z(n4128) );
  AND U4775 ( .A(a[106]), .B(b[3]), .Z(n4127) );
  XOR U4776 ( .A(n4128), .B(n4127), .Z(n4129) );
  XOR U4777 ( .A(n4130), .B(n4129), .Z(n4133) );
  NAND U4778 ( .A(b[0]), .B(a[109]), .Z(n4134) );
  XOR U4779 ( .A(n4133), .B(n4134), .Z(n4136) );
  OR U4780 ( .A(n4104), .B(n4103), .Z(n4108) );
  NANDN U4781 ( .A(n4106), .B(n4105), .Z(n4107) );
  NAND U4782 ( .A(n4108), .B(n4107), .Z(n4135) );
  XNOR U4783 ( .A(n4136), .B(n4135), .Z(n4121) );
  NANDN U4784 ( .A(n4110), .B(n4109), .Z(n4114) );
  OR U4785 ( .A(n4112), .B(n4111), .Z(n4113) );
  NAND U4786 ( .A(n4114), .B(n4113), .Z(n4122) );
  XNOR U4787 ( .A(n4121), .B(n4122), .Z(n4123) );
  XNOR U4788 ( .A(n4124), .B(n4123), .Z(n4140) );
  NAND U4789 ( .A(n4115), .B(sreg[1128]), .Z(n4119) );
  OR U4790 ( .A(n4117), .B(n4116), .Z(n4118) );
  AND U4791 ( .A(n4119), .B(n4118), .Z(n4139) );
  XNOR U4792 ( .A(n4139), .B(sreg[1129]), .Z(n4120) );
  XOR U4793 ( .A(n4140), .B(n4120), .Z(c[1129]) );
  NANDN U4794 ( .A(n4122), .B(n4121), .Z(n4126) );
  NAND U4795 ( .A(n4124), .B(n4123), .Z(n4125) );
  NAND U4796 ( .A(n4126), .B(n4125), .Z(n4147) );
  AND U4797 ( .A(b[2]), .B(a[108]), .Z(n4153) );
  AND U4798 ( .A(a[109]), .B(b[1]), .Z(n4151) );
  AND U4799 ( .A(a[107]), .B(b[3]), .Z(n4150) );
  XOR U4800 ( .A(n4151), .B(n4150), .Z(n4152) );
  XOR U4801 ( .A(n4153), .B(n4152), .Z(n4156) );
  NAND U4802 ( .A(b[0]), .B(a[110]), .Z(n4157) );
  XOR U4803 ( .A(n4156), .B(n4157), .Z(n4159) );
  OR U4804 ( .A(n4128), .B(n4127), .Z(n4132) );
  NANDN U4805 ( .A(n4130), .B(n4129), .Z(n4131) );
  NAND U4806 ( .A(n4132), .B(n4131), .Z(n4158) );
  XNOR U4807 ( .A(n4159), .B(n4158), .Z(n4144) );
  NANDN U4808 ( .A(n4134), .B(n4133), .Z(n4138) );
  OR U4809 ( .A(n4136), .B(n4135), .Z(n4137) );
  NAND U4810 ( .A(n4138), .B(n4137), .Z(n4145) );
  XNOR U4811 ( .A(n4144), .B(n4145), .Z(n4146) );
  XOR U4812 ( .A(n4147), .B(n4146), .Z(n4143) );
  XOR U4813 ( .A(sreg[1130]), .B(n4142), .Z(n4141) );
  XOR U4814 ( .A(n4143), .B(n4141), .Z(c[1130]) );
  NANDN U4815 ( .A(n4145), .B(n4144), .Z(n4149) );
  NAND U4816 ( .A(n4147), .B(n4146), .Z(n4148) );
  NAND U4817 ( .A(n4149), .B(n4148), .Z(n4165) );
  AND U4818 ( .A(b[2]), .B(a[109]), .Z(n4171) );
  AND U4819 ( .A(a[110]), .B(b[1]), .Z(n4169) );
  AND U4820 ( .A(a[108]), .B(b[3]), .Z(n4168) );
  XOR U4821 ( .A(n4169), .B(n4168), .Z(n4170) );
  XOR U4822 ( .A(n4171), .B(n4170), .Z(n4174) );
  NAND U4823 ( .A(b[0]), .B(a[111]), .Z(n4175) );
  XOR U4824 ( .A(n4174), .B(n4175), .Z(n4177) );
  OR U4825 ( .A(n4151), .B(n4150), .Z(n4155) );
  NANDN U4826 ( .A(n4153), .B(n4152), .Z(n4154) );
  NAND U4827 ( .A(n4155), .B(n4154), .Z(n4176) );
  XNOR U4828 ( .A(n4177), .B(n4176), .Z(n4162) );
  NANDN U4829 ( .A(n4157), .B(n4156), .Z(n4161) );
  OR U4830 ( .A(n4159), .B(n4158), .Z(n4160) );
  NAND U4831 ( .A(n4161), .B(n4160), .Z(n4163) );
  XNOR U4832 ( .A(n4162), .B(n4163), .Z(n4164) );
  XNOR U4833 ( .A(n4165), .B(n4164), .Z(n4180) );
  XNOR U4834 ( .A(n4180), .B(sreg[1131]), .Z(n4181) );
  XOR U4835 ( .A(n4182), .B(n4181), .Z(c[1131]) );
  NANDN U4836 ( .A(n4163), .B(n4162), .Z(n4167) );
  NAND U4837 ( .A(n4165), .B(n4164), .Z(n4166) );
  NAND U4838 ( .A(n4167), .B(n4166), .Z(n4188) );
  AND U4839 ( .A(b[2]), .B(a[110]), .Z(n4194) );
  AND U4840 ( .A(a[111]), .B(b[1]), .Z(n4192) );
  AND U4841 ( .A(a[109]), .B(b[3]), .Z(n4191) );
  XOR U4842 ( .A(n4192), .B(n4191), .Z(n4193) );
  XOR U4843 ( .A(n4194), .B(n4193), .Z(n4197) );
  NAND U4844 ( .A(b[0]), .B(a[112]), .Z(n4198) );
  XOR U4845 ( .A(n4197), .B(n4198), .Z(n4200) );
  OR U4846 ( .A(n4169), .B(n4168), .Z(n4173) );
  NANDN U4847 ( .A(n4171), .B(n4170), .Z(n4172) );
  NAND U4848 ( .A(n4173), .B(n4172), .Z(n4199) );
  XNOR U4849 ( .A(n4200), .B(n4199), .Z(n4185) );
  NANDN U4850 ( .A(n4175), .B(n4174), .Z(n4179) );
  OR U4851 ( .A(n4177), .B(n4176), .Z(n4178) );
  NAND U4852 ( .A(n4179), .B(n4178), .Z(n4186) );
  XNOR U4853 ( .A(n4185), .B(n4186), .Z(n4187) );
  XNOR U4854 ( .A(n4188), .B(n4187), .Z(n4203) );
  XNOR U4855 ( .A(n4203), .B(sreg[1132]), .Z(n4205) );
  NAND U4856 ( .A(n4180), .B(sreg[1131]), .Z(n4184) );
  OR U4857 ( .A(n4182), .B(n4181), .Z(n4183) );
  AND U4858 ( .A(n4184), .B(n4183), .Z(n4204) );
  XOR U4859 ( .A(n4205), .B(n4204), .Z(c[1132]) );
  NANDN U4860 ( .A(n4186), .B(n4185), .Z(n4190) );
  NAND U4861 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U4862 ( .A(n4190), .B(n4189), .Z(n4211) );
  AND U4863 ( .A(b[2]), .B(a[111]), .Z(n4217) );
  AND U4864 ( .A(a[112]), .B(b[1]), .Z(n4215) );
  AND U4865 ( .A(a[110]), .B(b[3]), .Z(n4214) );
  XOR U4866 ( .A(n4215), .B(n4214), .Z(n4216) );
  XOR U4867 ( .A(n4217), .B(n4216), .Z(n4220) );
  NAND U4868 ( .A(b[0]), .B(a[113]), .Z(n4221) );
  XOR U4869 ( .A(n4220), .B(n4221), .Z(n4223) );
  OR U4870 ( .A(n4192), .B(n4191), .Z(n4196) );
  NANDN U4871 ( .A(n4194), .B(n4193), .Z(n4195) );
  NAND U4872 ( .A(n4196), .B(n4195), .Z(n4222) );
  XNOR U4873 ( .A(n4223), .B(n4222), .Z(n4208) );
  NANDN U4874 ( .A(n4198), .B(n4197), .Z(n4202) );
  OR U4875 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U4876 ( .A(n4202), .B(n4201), .Z(n4209) );
  XNOR U4877 ( .A(n4208), .B(n4209), .Z(n4210) );
  XNOR U4878 ( .A(n4211), .B(n4210), .Z(n4226) );
  XOR U4879 ( .A(sreg[1133]), .B(n4226), .Z(n4227) );
  NAND U4880 ( .A(n4203), .B(sreg[1132]), .Z(n4207) );
  OR U4881 ( .A(n4205), .B(n4204), .Z(n4206) );
  NAND U4882 ( .A(n4207), .B(n4206), .Z(n4228) );
  XOR U4883 ( .A(n4227), .B(n4228), .Z(c[1133]) );
  NANDN U4884 ( .A(n4209), .B(n4208), .Z(n4213) );
  NAND U4885 ( .A(n4211), .B(n4210), .Z(n4212) );
  NAND U4886 ( .A(n4213), .B(n4212), .Z(n4234) );
  AND U4887 ( .A(b[2]), .B(a[112]), .Z(n4240) );
  AND U4888 ( .A(a[113]), .B(b[1]), .Z(n4238) );
  AND U4889 ( .A(a[111]), .B(b[3]), .Z(n4237) );
  XOR U4890 ( .A(n4238), .B(n4237), .Z(n4239) );
  XOR U4891 ( .A(n4240), .B(n4239), .Z(n4243) );
  NAND U4892 ( .A(b[0]), .B(a[114]), .Z(n4244) );
  XOR U4893 ( .A(n4243), .B(n4244), .Z(n4246) );
  OR U4894 ( .A(n4215), .B(n4214), .Z(n4219) );
  NANDN U4895 ( .A(n4217), .B(n4216), .Z(n4218) );
  NAND U4896 ( .A(n4219), .B(n4218), .Z(n4245) );
  XNOR U4897 ( .A(n4246), .B(n4245), .Z(n4231) );
  NANDN U4898 ( .A(n4221), .B(n4220), .Z(n4225) );
  OR U4899 ( .A(n4223), .B(n4222), .Z(n4224) );
  NAND U4900 ( .A(n4225), .B(n4224), .Z(n4232) );
  XNOR U4901 ( .A(n4231), .B(n4232), .Z(n4233) );
  XNOR U4902 ( .A(n4234), .B(n4233), .Z(n4249) );
  XNOR U4903 ( .A(n4249), .B(sreg[1134]), .Z(n4251) );
  OR U4904 ( .A(n4226), .B(sreg[1133]), .Z(n4230) );
  NANDN U4905 ( .A(n4228), .B(n4227), .Z(n4229) );
  NAND U4906 ( .A(n4230), .B(n4229), .Z(n4250) );
  XOR U4907 ( .A(n4251), .B(n4250), .Z(c[1134]) );
  NANDN U4908 ( .A(n4232), .B(n4231), .Z(n4236) );
  NAND U4909 ( .A(n4234), .B(n4233), .Z(n4235) );
  NAND U4910 ( .A(n4236), .B(n4235), .Z(n4257) );
  AND U4911 ( .A(b[2]), .B(a[113]), .Z(n4263) );
  AND U4912 ( .A(a[114]), .B(b[1]), .Z(n4261) );
  AND U4913 ( .A(a[112]), .B(b[3]), .Z(n4260) );
  XOR U4914 ( .A(n4261), .B(n4260), .Z(n4262) );
  XOR U4915 ( .A(n4263), .B(n4262), .Z(n4266) );
  NAND U4916 ( .A(b[0]), .B(a[115]), .Z(n4267) );
  XOR U4917 ( .A(n4266), .B(n4267), .Z(n4269) );
  OR U4918 ( .A(n4238), .B(n4237), .Z(n4242) );
  NANDN U4919 ( .A(n4240), .B(n4239), .Z(n4241) );
  NAND U4920 ( .A(n4242), .B(n4241), .Z(n4268) );
  XNOR U4921 ( .A(n4269), .B(n4268), .Z(n4254) );
  NANDN U4922 ( .A(n4244), .B(n4243), .Z(n4248) );
  OR U4923 ( .A(n4246), .B(n4245), .Z(n4247) );
  NAND U4924 ( .A(n4248), .B(n4247), .Z(n4255) );
  XNOR U4925 ( .A(n4254), .B(n4255), .Z(n4256) );
  XNOR U4926 ( .A(n4257), .B(n4256), .Z(n4272) );
  XNOR U4927 ( .A(n4272), .B(sreg[1135]), .Z(n4274) );
  NAND U4928 ( .A(n4249), .B(sreg[1134]), .Z(n4253) );
  OR U4929 ( .A(n4251), .B(n4250), .Z(n4252) );
  AND U4930 ( .A(n4253), .B(n4252), .Z(n4273) );
  XOR U4931 ( .A(n4274), .B(n4273), .Z(c[1135]) );
  NANDN U4932 ( .A(n4255), .B(n4254), .Z(n4259) );
  NAND U4933 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U4934 ( .A(n4259), .B(n4258), .Z(n4283) );
  AND U4935 ( .A(b[2]), .B(a[114]), .Z(n4295) );
  AND U4936 ( .A(a[115]), .B(b[1]), .Z(n4293) );
  AND U4937 ( .A(a[113]), .B(b[3]), .Z(n4292) );
  XOR U4938 ( .A(n4293), .B(n4292), .Z(n4294) );
  XOR U4939 ( .A(n4295), .B(n4294), .Z(n4286) );
  NAND U4940 ( .A(b[0]), .B(a[116]), .Z(n4287) );
  XOR U4941 ( .A(n4286), .B(n4287), .Z(n4289) );
  OR U4942 ( .A(n4261), .B(n4260), .Z(n4265) );
  NANDN U4943 ( .A(n4263), .B(n4262), .Z(n4264) );
  NAND U4944 ( .A(n4265), .B(n4264), .Z(n4288) );
  XNOR U4945 ( .A(n4289), .B(n4288), .Z(n4280) );
  NANDN U4946 ( .A(n4267), .B(n4266), .Z(n4271) );
  OR U4947 ( .A(n4269), .B(n4268), .Z(n4270) );
  NAND U4948 ( .A(n4271), .B(n4270), .Z(n4281) );
  XNOR U4949 ( .A(n4280), .B(n4281), .Z(n4282) );
  XOR U4950 ( .A(n4283), .B(n4282), .Z(n4279) );
  NAND U4951 ( .A(n4272), .B(sreg[1135]), .Z(n4276) );
  OR U4952 ( .A(n4274), .B(n4273), .Z(n4275) );
  NAND U4953 ( .A(n4276), .B(n4275), .Z(n4278) );
  XNOR U4954 ( .A(sreg[1136]), .B(n4278), .Z(n4277) );
  XOR U4955 ( .A(n4279), .B(n4277), .Z(c[1136]) );
  NANDN U4956 ( .A(n4281), .B(n4280), .Z(n4285) );
  NAND U4957 ( .A(n4283), .B(n4282), .Z(n4284) );
  NAND U4958 ( .A(n4285), .B(n4284), .Z(n4313) );
  NANDN U4959 ( .A(n4287), .B(n4286), .Z(n4291) );
  OR U4960 ( .A(n4289), .B(n4288), .Z(n4290) );
  NAND U4961 ( .A(n4291), .B(n4290), .Z(n4310) );
  AND U4962 ( .A(b[2]), .B(a[115]), .Z(n4301) );
  AND U4963 ( .A(a[116]), .B(b[1]), .Z(n4299) );
  AND U4964 ( .A(a[114]), .B(b[3]), .Z(n4298) );
  XOR U4965 ( .A(n4299), .B(n4298), .Z(n4300) );
  XOR U4966 ( .A(n4301), .B(n4300), .Z(n4304) );
  NAND U4967 ( .A(b[0]), .B(a[117]), .Z(n4305) );
  XNOR U4968 ( .A(n4304), .B(n4305), .Z(n4306) );
  OR U4969 ( .A(n4293), .B(n4292), .Z(n4297) );
  NANDN U4970 ( .A(n4295), .B(n4294), .Z(n4296) );
  AND U4971 ( .A(n4297), .B(n4296), .Z(n4307) );
  XNOR U4972 ( .A(n4306), .B(n4307), .Z(n4311) );
  XNOR U4973 ( .A(n4310), .B(n4311), .Z(n4312) );
  XNOR U4974 ( .A(n4313), .B(n4312), .Z(n4316) );
  XNOR U4975 ( .A(sreg[1137]), .B(n4316), .Z(n4317) );
  XOR U4976 ( .A(n4318), .B(n4317), .Z(c[1137]) );
  AND U4977 ( .A(b[2]), .B(a[116]), .Z(n4331) );
  AND U4978 ( .A(a[117]), .B(b[1]), .Z(n4329) );
  AND U4979 ( .A(a[115]), .B(b[3]), .Z(n4328) );
  XOR U4980 ( .A(n4329), .B(n4328), .Z(n4330) );
  XOR U4981 ( .A(n4331), .B(n4330), .Z(n4334) );
  NAND U4982 ( .A(b[0]), .B(a[118]), .Z(n4335) );
  XOR U4983 ( .A(n4334), .B(n4335), .Z(n4337) );
  OR U4984 ( .A(n4299), .B(n4298), .Z(n4303) );
  NANDN U4985 ( .A(n4301), .B(n4300), .Z(n4302) );
  NAND U4986 ( .A(n4303), .B(n4302), .Z(n4336) );
  XNOR U4987 ( .A(n4337), .B(n4336), .Z(n4322) );
  NANDN U4988 ( .A(n4305), .B(n4304), .Z(n4309) );
  NAND U4989 ( .A(n4307), .B(n4306), .Z(n4308) );
  NAND U4990 ( .A(n4309), .B(n4308), .Z(n4323) );
  XNOR U4991 ( .A(n4322), .B(n4323), .Z(n4324) );
  NANDN U4992 ( .A(n4311), .B(n4310), .Z(n4315) );
  NANDN U4993 ( .A(n4313), .B(n4312), .Z(n4314) );
  NAND U4994 ( .A(n4315), .B(n4314), .Z(n4325) );
  XOR U4995 ( .A(n4324), .B(n4325), .Z(n4341) );
  NAND U4996 ( .A(sreg[1137]), .B(n4316), .Z(n4320) );
  OR U4997 ( .A(n4318), .B(n4317), .Z(n4319) );
  NAND U4998 ( .A(n4320), .B(n4319), .Z(n4340) );
  XNOR U4999 ( .A(sreg[1138]), .B(n4340), .Z(n4321) );
  XNOR U5000 ( .A(n4341), .B(n4321), .Z(c[1138]) );
  NANDN U5001 ( .A(n4323), .B(n4322), .Z(n4327) );
  NANDN U5002 ( .A(n4325), .B(n4324), .Z(n4326) );
  NAND U5003 ( .A(n4327), .B(n4326), .Z(n4358) );
  AND U5004 ( .A(b[2]), .B(a[117]), .Z(n4352) );
  AND U5005 ( .A(a[118]), .B(b[1]), .Z(n4350) );
  AND U5006 ( .A(a[116]), .B(b[3]), .Z(n4349) );
  XOR U5007 ( .A(n4350), .B(n4349), .Z(n4351) );
  XOR U5008 ( .A(n4352), .B(n4351), .Z(n4343) );
  NAND U5009 ( .A(b[0]), .B(a[119]), .Z(n4344) );
  XOR U5010 ( .A(n4343), .B(n4344), .Z(n4346) );
  OR U5011 ( .A(n4329), .B(n4328), .Z(n4333) );
  NANDN U5012 ( .A(n4331), .B(n4330), .Z(n4332) );
  NAND U5013 ( .A(n4333), .B(n4332), .Z(n4345) );
  XNOR U5014 ( .A(n4346), .B(n4345), .Z(n4355) );
  NANDN U5015 ( .A(n4335), .B(n4334), .Z(n4339) );
  OR U5016 ( .A(n4337), .B(n4336), .Z(n4338) );
  NAND U5017 ( .A(n4339), .B(n4338), .Z(n4356) );
  XNOR U5018 ( .A(n4355), .B(n4356), .Z(n4357) );
  XOR U5019 ( .A(n4358), .B(n4357), .Z(n4362) );
  XNOR U5020 ( .A(sreg[1139]), .B(n4361), .Z(n4342) );
  XOR U5021 ( .A(n4362), .B(n4342), .Z(c[1139]) );
  NANDN U5022 ( .A(n4344), .B(n4343), .Z(n4348) );
  OR U5023 ( .A(n4346), .B(n4345), .Z(n4347) );
  NAND U5024 ( .A(n4348), .B(n4347), .Z(n4364) );
  AND U5025 ( .A(b[2]), .B(a[118]), .Z(n4373) );
  AND U5026 ( .A(a[119]), .B(b[1]), .Z(n4371) );
  AND U5027 ( .A(a[117]), .B(b[3]), .Z(n4370) );
  XOR U5028 ( .A(n4371), .B(n4370), .Z(n4372) );
  XOR U5029 ( .A(n4373), .B(n4372), .Z(n4376) );
  NAND U5030 ( .A(b[0]), .B(a[120]), .Z(n4377) );
  XNOR U5031 ( .A(n4376), .B(n4377), .Z(n4378) );
  OR U5032 ( .A(n4350), .B(n4349), .Z(n4354) );
  NANDN U5033 ( .A(n4352), .B(n4351), .Z(n4353) );
  AND U5034 ( .A(n4354), .B(n4353), .Z(n4379) );
  XNOR U5035 ( .A(n4378), .B(n4379), .Z(n4365) );
  XNOR U5036 ( .A(n4364), .B(n4365), .Z(n4366) );
  NANDN U5037 ( .A(n4356), .B(n4355), .Z(n4360) );
  NAND U5038 ( .A(n4358), .B(n4357), .Z(n4359) );
  AND U5039 ( .A(n4360), .B(n4359), .Z(n4367) );
  XNOR U5040 ( .A(n4366), .B(n4367), .Z(n4383) );
  XNOR U5041 ( .A(sreg[1140]), .B(n4382), .Z(n4363) );
  XOR U5042 ( .A(n4383), .B(n4363), .Z(c[1140]) );
  NANDN U5043 ( .A(n4365), .B(n4364), .Z(n4369) );
  NAND U5044 ( .A(n4367), .B(n4366), .Z(n4368) );
  NAND U5045 ( .A(n4369), .B(n4368), .Z(n4388) );
  AND U5046 ( .A(b[2]), .B(a[119]), .Z(n4394) );
  AND U5047 ( .A(a[120]), .B(b[1]), .Z(n4392) );
  AND U5048 ( .A(a[118]), .B(b[3]), .Z(n4391) );
  XOR U5049 ( .A(n4392), .B(n4391), .Z(n4393) );
  XOR U5050 ( .A(n4394), .B(n4393), .Z(n4397) );
  NAND U5051 ( .A(b[0]), .B(a[121]), .Z(n4398) );
  XOR U5052 ( .A(n4397), .B(n4398), .Z(n4400) );
  OR U5053 ( .A(n4371), .B(n4370), .Z(n4375) );
  NANDN U5054 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U5055 ( .A(n4375), .B(n4374), .Z(n4399) );
  XNOR U5056 ( .A(n4400), .B(n4399), .Z(n4385) );
  NANDN U5057 ( .A(n4377), .B(n4376), .Z(n4381) );
  NAND U5058 ( .A(n4379), .B(n4378), .Z(n4380) );
  NAND U5059 ( .A(n4381), .B(n4380), .Z(n4386) );
  XNOR U5060 ( .A(n4385), .B(n4386), .Z(n4387) );
  XOR U5061 ( .A(n4388), .B(n4387), .Z(n4404) );
  XNOR U5062 ( .A(sreg[1141]), .B(n4403), .Z(n4384) );
  XNOR U5063 ( .A(n4404), .B(n4384), .Z(c[1141]) );
  NANDN U5064 ( .A(n4386), .B(n4385), .Z(n4390) );
  NANDN U5065 ( .A(n4388), .B(n4387), .Z(n4389) );
  NAND U5066 ( .A(n4390), .B(n4389), .Z(n4409) );
  AND U5067 ( .A(b[2]), .B(a[120]), .Z(n4415) );
  AND U5068 ( .A(a[121]), .B(b[1]), .Z(n4413) );
  AND U5069 ( .A(a[119]), .B(b[3]), .Z(n4412) );
  XOR U5070 ( .A(n4413), .B(n4412), .Z(n4414) );
  XOR U5071 ( .A(n4415), .B(n4414), .Z(n4418) );
  NAND U5072 ( .A(b[0]), .B(a[122]), .Z(n4419) );
  XOR U5073 ( .A(n4418), .B(n4419), .Z(n4421) );
  OR U5074 ( .A(n4392), .B(n4391), .Z(n4396) );
  NANDN U5075 ( .A(n4394), .B(n4393), .Z(n4395) );
  NAND U5076 ( .A(n4396), .B(n4395), .Z(n4420) );
  XNOR U5077 ( .A(n4421), .B(n4420), .Z(n4406) );
  NANDN U5078 ( .A(n4398), .B(n4397), .Z(n4402) );
  OR U5079 ( .A(n4400), .B(n4399), .Z(n4401) );
  NAND U5080 ( .A(n4402), .B(n4401), .Z(n4407) );
  XNOR U5081 ( .A(n4406), .B(n4407), .Z(n4408) );
  XNOR U5082 ( .A(n4409), .B(n4408), .Z(n4425) );
  XOR U5083 ( .A(n4424), .B(sreg[1142]), .Z(n4405) );
  XOR U5084 ( .A(n4425), .B(n4405), .Z(c[1142]) );
  NANDN U5085 ( .A(n4407), .B(n4406), .Z(n4411) );
  NAND U5086 ( .A(n4409), .B(n4408), .Z(n4410) );
  NAND U5087 ( .A(n4411), .B(n4410), .Z(n4432) );
  AND U5088 ( .A(b[2]), .B(a[121]), .Z(n4438) );
  AND U5089 ( .A(a[122]), .B(b[1]), .Z(n4436) );
  AND U5090 ( .A(a[120]), .B(b[3]), .Z(n4435) );
  XOR U5091 ( .A(n4436), .B(n4435), .Z(n4437) );
  XOR U5092 ( .A(n4438), .B(n4437), .Z(n4441) );
  NAND U5093 ( .A(b[0]), .B(a[123]), .Z(n4442) );
  XOR U5094 ( .A(n4441), .B(n4442), .Z(n4444) );
  OR U5095 ( .A(n4413), .B(n4412), .Z(n4417) );
  NANDN U5096 ( .A(n4415), .B(n4414), .Z(n4416) );
  NAND U5097 ( .A(n4417), .B(n4416), .Z(n4443) );
  XNOR U5098 ( .A(n4444), .B(n4443), .Z(n4429) );
  NANDN U5099 ( .A(n4419), .B(n4418), .Z(n4423) );
  OR U5100 ( .A(n4421), .B(n4420), .Z(n4422) );
  NAND U5101 ( .A(n4423), .B(n4422), .Z(n4430) );
  XNOR U5102 ( .A(n4429), .B(n4430), .Z(n4431) );
  XNOR U5103 ( .A(n4432), .B(n4431), .Z(n4428) );
  XOR U5104 ( .A(n4427), .B(sreg[1143]), .Z(n4426) );
  XOR U5105 ( .A(n4428), .B(n4426), .Z(c[1143]) );
  NANDN U5106 ( .A(n4430), .B(n4429), .Z(n4434) );
  NAND U5107 ( .A(n4432), .B(n4431), .Z(n4433) );
  NAND U5108 ( .A(n4434), .B(n4433), .Z(n4455) );
  AND U5109 ( .A(b[2]), .B(a[122]), .Z(n4461) );
  AND U5110 ( .A(a[123]), .B(b[1]), .Z(n4459) );
  AND U5111 ( .A(a[121]), .B(b[3]), .Z(n4458) );
  XOR U5112 ( .A(n4459), .B(n4458), .Z(n4460) );
  XOR U5113 ( .A(n4461), .B(n4460), .Z(n4464) );
  NAND U5114 ( .A(b[0]), .B(a[124]), .Z(n4465) );
  XOR U5115 ( .A(n4464), .B(n4465), .Z(n4467) );
  OR U5116 ( .A(n4436), .B(n4435), .Z(n4440) );
  NANDN U5117 ( .A(n4438), .B(n4437), .Z(n4439) );
  NAND U5118 ( .A(n4440), .B(n4439), .Z(n4466) );
  XNOR U5119 ( .A(n4467), .B(n4466), .Z(n4452) );
  NANDN U5120 ( .A(n4442), .B(n4441), .Z(n4446) );
  OR U5121 ( .A(n4444), .B(n4443), .Z(n4445) );
  NAND U5122 ( .A(n4446), .B(n4445), .Z(n4453) );
  XNOR U5123 ( .A(n4452), .B(n4453), .Z(n4454) );
  XNOR U5124 ( .A(n4455), .B(n4454), .Z(n4447) );
  XNOR U5125 ( .A(n4447), .B(sreg[1144]), .Z(n4449) );
  XNOR U5126 ( .A(n4448), .B(n4449), .Z(c[1144]) );
  NAND U5127 ( .A(n4447), .B(sreg[1144]), .Z(n4451) );
  NANDN U5128 ( .A(n4449), .B(n4448), .Z(n4450) );
  AND U5129 ( .A(n4451), .B(n4450), .Z(n4490) );
  NANDN U5130 ( .A(n4453), .B(n4452), .Z(n4457) );
  NAND U5131 ( .A(n4455), .B(n4454), .Z(n4456) );
  NAND U5132 ( .A(n4457), .B(n4456), .Z(n4474) );
  AND U5133 ( .A(b[2]), .B(a[123]), .Z(n4480) );
  AND U5134 ( .A(a[124]), .B(b[1]), .Z(n4478) );
  AND U5135 ( .A(a[122]), .B(b[3]), .Z(n4477) );
  XOR U5136 ( .A(n4478), .B(n4477), .Z(n4479) );
  XOR U5137 ( .A(n4480), .B(n4479), .Z(n4483) );
  NAND U5138 ( .A(b[0]), .B(a[125]), .Z(n4484) );
  XOR U5139 ( .A(n4483), .B(n4484), .Z(n4486) );
  OR U5140 ( .A(n4459), .B(n4458), .Z(n4463) );
  NANDN U5141 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U5142 ( .A(n4463), .B(n4462), .Z(n4485) );
  XNOR U5143 ( .A(n4486), .B(n4485), .Z(n4471) );
  NANDN U5144 ( .A(n4465), .B(n4464), .Z(n4469) );
  OR U5145 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U5146 ( .A(n4469), .B(n4468), .Z(n4472) );
  XNOR U5147 ( .A(n4471), .B(n4472), .Z(n4473) );
  XNOR U5148 ( .A(n4474), .B(n4473), .Z(n4489) );
  XNOR U5149 ( .A(sreg[1145]), .B(n4489), .Z(n4470) );
  XOR U5150 ( .A(n4490), .B(n4470), .Z(c[1145]) );
  NANDN U5151 ( .A(n4472), .B(n4471), .Z(n4476) );
  NAND U5152 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U5153 ( .A(n4476), .B(n4475), .Z(n4497) );
  AND U5154 ( .A(b[2]), .B(a[124]), .Z(n4503) );
  AND U5155 ( .A(a[125]), .B(b[1]), .Z(n4501) );
  AND U5156 ( .A(a[123]), .B(b[3]), .Z(n4500) );
  XOR U5157 ( .A(n4501), .B(n4500), .Z(n4502) );
  XOR U5158 ( .A(n4503), .B(n4502), .Z(n4506) );
  NAND U5159 ( .A(b[0]), .B(a[126]), .Z(n4507) );
  XOR U5160 ( .A(n4506), .B(n4507), .Z(n4509) );
  OR U5161 ( .A(n4478), .B(n4477), .Z(n4482) );
  NANDN U5162 ( .A(n4480), .B(n4479), .Z(n4481) );
  NAND U5163 ( .A(n4482), .B(n4481), .Z(n4508) );
  XNOR U5164 ( .A(n4509), .B(n4508), .Z(n4494) );
  NANDN U5165 ( .A(n4484), .B(n4483), .Z(n4488) );
  OR U5166 ( .A(n4486), .B(n4485), .Z(n4487) );
  NAND U5167 ( .A(n4488), .B(n4487), .Z(n4495) );
  XNOR U5168 ( .A(n4494), .B(n4495), .Z(n4496) );
  XOR U5169 ( .A(n4497), .B(n4496), .Z(n4493) );
  XNOR U5170 ( .A(sreg[1146]), .B(n4492), .Z(n4491) );
  XOR U5171 ( .A(n4493), .B(n4491), .Z(c[1146]) );
  NANDN U5172 ( .A(n4495), .B(n4494), .Z(n4499) );
  NAND U5173 ( .A(n4497), .B(n4496), .Z(n4498) );
  NAND U5174 ( .A(n4499), .B(n4498), .Z(n4515) );
  AND U5175 ( .A(b[2]), .B(a[125]), .Z(n4521) );
  AND U5176 ( .A(a[126]), .B(b[1]), .Z(n4519) );
  AND U5177 ( .A(a[124]), .B(b[3]), .Z(n4518) );
  XOR U5178 ( .A(n4519), .B(n4518), .Z(n4520) );
  XOR U5179 ( .A(n4521), .B(n4520), .Z(n4524) );
  NAND U5180 ( .A(b[0]), .B(a[127]), .Z(n4525) );
  XOR U5181 ( .A(n4524), .B(n4525), .Z(n4527) );
  OR U5182 ( .A(n4501), .B(n4500), .Z(n4505) );
  NANDN U5183 ( .A(n4503), .B(n4502), .Z(n4504) );
  NAND U5184 ( .A(n4505), .B(n4504), .Z(n4526) );
  XNOR U5185 ( .A(n4527), .B(n4526), .Z(n4512) );
  NANDN U5186 ( .A(n4507), .B(n4506), .Z(n4511) );
  OR U5187 ( .A(n4509), .B(n4508), .Z(n4510) );
  NAND U5188 ( .A(n4511), .B(n4510), .Z(n4513) );
  XNOR U5189 ( .A(n4512), .B(n4513), .Z(n4514) );
  XNOR U5190 ( .A(n4515), .B(n4514), .Z(n4530) );
  XNOR U5191 ( .A(n4530), .B(sreg[1147]), .Z(n4531) );
  XOR U5192 ( .A(n4532), .B(n4531), .Z(c[1147]) );
  NANDN U5193 ( .A(n4513), .B(n4512), .Z(n4517) );
  NAND U5194 ( .A(n4515), .B(n4514), .Z(n4516) );
  NAND U5195 ( .A(n4517), .B(n4516), .Z(n4538) );
  AND U5196 ( .A(b[2]), .B(a[126]), .Z(n4544) );
  AND U5197 ( .A(a[127]), .B(b[1]), .Z(n4542) );
  AND U5198 ( .A(a[125]), .B(b[3]), .Z(n4541) );
  XOR U5199 ( .A(n4542), .B(n4541), .Z(n4543) );
  XOR U5200 ( .A(n4544), .B(n4543), .Z(n4547) );
  NAND U5201 ( .A(b[0]), .B(a[128]), .Z(n4548) );
  XOR U5202 ( .A(n4547), .B(n4548), .Z(n4550) );
  OR U5203 ( .A(n4519), .B(n4518), .Z(n4523) );
  NANDN U5204 ( .A(n4521), .B(n4520), .Z(n4522) );
  NAND U5205 ( .A(n4523), .B(n4522), .Z(n4549) );
  XNOR U5206 ( .A(n4550), .B(n4549), .Z(n4535) );
  NANDN U5207 ( .A(n4525), .B(n4524), .Z(n4529) );
  OR U5208 ( .A(n4527), .B(n4526), .Z(n4528) );
  NAND U5209 ( .A(n4529), .B(n4528), .Z(n4536) );
  XNOR U5210 ( .A(n4535), .B(n4536), .Z(n4537) );
  XNOR U5211 ( .A(n4538), .B(n4537), .Z(n4553) );
  XNOR U5212 ( .A(n4553), .B(sreg[1148]), .Z(n4555) );
  NAND U5213 ( .A(n4530), .B(sreg[1147]), .Z(n4534) );
  OR U5214 ( .A(n4532), .B(n4531), .Z(n4533) );
  AND U5215 ( .A(n4534), .B(n4533), .Z(n4554) );
  XOR U5216 ( .A(n4555), .B(n4554), .Z(c[1148]) );
  NANDN U5217 ( .A(n4536), .B(n4535), .Z(n4540) );
  NAND U5218 ( .A(n4538), .B(n4537), .Z(n4539) );
  NAND U5219 ( .A(n4540), .B(n4539), .Z(n4561) );
  AND U5220 ( .A(b[2]), .B(a[127]), .Z(n4567) );
  AND U5221 ( .A(a[128]), .B(b[1]), .Z(n4565) );
  AND U5222 ( .A(a[126]), .B(b[3]), .Z(n4564) );
  XOR U5223 ( .A(n4565), .B(n4564), .Z(n4566) );
  XOR U5224 ( .A(n4567), .B(n4566), .Z(n4570) );
  NAND U5225 ( .A(b[0]), .B(a[129]), .Z(n4571) );
  XOR U5226 ( .A(n4570), .B(n4571), .Z(n4573) );
  OR U5227 ( .A(n4542), .B(n4541), .Z(n4546) );
  NANDN U5228 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U5229 ( .A(n4546), .B(n4545), .Z(n4572) );
  XNOR U5230 ( .A(n4573), .B(n4572), .Z(n4558) );
  NANDN U5231 ( .A(n4548), .B(n4547), .Z(n4552) );
  OR U5232 ( .A(n4550), .B(n4549), .Z(n4551) );
  NAND U5233 ( .A(n4552), .B(n4551), .Z(n4559) );
  XNOR U5234 ( .A(n4558), .B(n4559), .Z(n4560) );
  XNOR U5235 ( .A(n4561), .B(n4560), .Z(n4576) );
  XOR U5236 ( .A(sreg[1149]), .B(n4576), .Z(n4577) );
  NAND U5237 ( .A(n4553), .B(sreg[1148]), .Z(n4557) );
  OR U5238 ( .A(n4555), .B(n4554), .Z(n4556) );
  NAND U5239 ( .A(n4557), .B(n4556), .Z(n4578) );
  XOR U5240 ( .A(n4577), .B(n4578), .Z(c[1149]) );
  NANDN U5241 ( .A(n4559), .B(n4558), .Z(n4563) );
  NAND U5242 ( .A(n4561), .B(n4560), .Z(n4562) );
  NAND U5243 ( .A(n4563), .B(n4562), .Z(n4587) );
  AND U5244 ( .A(b[2]), .B(a[128]), .Z(n4593) );
  AND U5245 ( .A(a[129]), .B(b[1]), .Z(n4591) );
  AND U5246 ( .A(a[127]), .B(b[3]), .Z(n4590) );
  XOR U5247 ( .A(n4591), .B(n4590), .Z(n4592) );
  XOR U5248 ( .A(n4593), .B(n4592), .Z(n4596) );
  NAND U5249 ( .A(b[0]), .B(a[130]), .Z(n4597) );
  XOR U5250 ( .A(n4596), .B(n4597), .Z(n4599) );
  OR U5251 ( .A(n4565), .B(n4564), .Z(n4569) );
  NANDN U5252 ( .A(n4567), .B(n4566), .Z(n4568) );
  NAND U5253 ( .A(n4569), .B(n4568), .Z(n4598) );
  XNOR U5254 ( .A(n4599), .B(n4598), .Z(n4584) );
  NANDN U5255 ( .A(n4571), .B(n4570), .Z(n4575) );
  OR U5256 ( .A(n4573), .B(n4572), .Z(n4574) );
  NAND U5257 ( .A(n4575), .B(n4574), .Z(n4585) );
  XNOR U5258 ( .A(n4584), .B(n4585), .Z(n4586) );
  XOR U5259 ( .A(n4587), .B(n4586), .Z(n4583) );
  OR U5260 ( .A(n4576), .B(sreg[1149]), .Z(n4580) );
  NANDN U5261 ( .A(n4578), .B(n4577), .Z(n4579) );
  AND U5262 ( .A(n4580), .B(n4579), .Z(n4582) );
  XNOR U5263 ( .A(sreg[1150]), .B(n4582), .Z(n4581) );
  XOR U5264 ( .A(n4583), .B(n4581), .Z(c[1150]) );
  NANDN U5265 ( .A(n4585), .B(n4584), .Z(n4589) );
  NAND U5266 ( .A(n4587), .B(n4586), .Z(n4588) );
  NAND U5267 ( .A(n4589), .B(n4588), .Z(n4605) );
  AND U5268 ( .A(b[2]), .B(a[129]), .Z(n4611) );
  AND U5269 ( .A(a[130]), .B(b[1]), .Z(n4609) );
  AND U5270 ( .A(a[128]), .B(b[3]), .Z(n4608) );
  XOR U5271 ( .A(n4609), .B(n4608), .Z(n4610) );
  XOR U5272 ( .A(n4611), .B(n4610), .Z(n4614) );
  NAND U5273 ( .A(b[0]), .B(a[131]), .Z(n4615) );
  XOR U5274 ( .A(n4614), .B(n4615), .Z(n4617) );
  OR U5275 ( .A(n4591), .B(n4590), .Z(n4595) );
  NANDN U5276 ( .A(n4593), .B(n4592), .Z(n4594) );
  NAND U5277 ( .A(n4595), .B(n4594), .Z(n4616) );
  XNOR U5278 ( .A(n4617), .B(n4616), .Z(n4602) );
  NANDN U5279 ( .A(n4597), .B(n4596), .Z(n4601) );
  OR U5280 ( .A(n4599), .B(n4598), .Z(n4600) );
  NAND U5281 ( .A(n4601), .B(n4600), .Z(n4603) );
  XNOR U5282 ( .A(n4602), .B(n4603), .Z(n4604) );
  XNOR U5283 ( .A(n4605), .B(n4604), .Z(n4620) );
  XNOR U5284 ( .A(n4620), .B(sreg[1151]), .Z(n4621) );
  XOR U5285 ( .A(n4622), .B(n4621), .Z(c[1151]) );
  NANDN U5286 ( .A(n4603), .B(n4602), .Z(n4607) );
  NAND U5287 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U5288 ( .A(n4607), .B(n4606), .Z(n4628) );
  AND U5289 ( .A(b[2]), .B(a[130]), .Z(n4640) );
  AND U5290 ( .A(a[131]), .B(b[1]), .Z(n4638) );
  AND U5291 ( .A(a[129]), .B(b[3]), .Z(n4637) );
  XOR U5292 ( .A(n4638), .B(n4637), .Z(n4639) );
  XOR U5293 ( .A(n4640), .B(n4639), .Z(n4631) );
  NAND U5294 ( .A(b[0]), .B(a[132]), .Z(n4632) );
  XOR U5295 ( .A(n4631), .B(n4632), .Z(n4634) );
  OR U5296 ( .A(n4609), .B(n4608), .Z(n4613) );
  NANDN U5297 ( .A(n4611), .B(n4610), .Z(n4612) );
  NAND U5298 ( .A(n4613), .B(n4612), .Z(n4633) );
  XNOR U5299 ( .A(n4634), .B(n4633), .Z(n4625) );
  NANDN U5300 ( .A(n4615), .B(n4614), .Z(n4619) );
  OR U5301 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U5302 ( .A(n4619), .B(n4618), .Z(n4626) );
  XNOR U5303 ( .A(n4625), .B(n4626), .Z(n4627) );
  XNOR U5304 ( .A(n4628), .B(n4627), .Z(n4643) );
  XNOR U5305 ( .A(n4643), .B(sreg[1152]), .Z(n4645) );
  NAND U5306 ( .A(n4620), .B(sreg[1151]), .Z(n4624) );
  OR U5307 ( .A(n4622), .B(n4621), .Z(n4623) );
  AND U5308 ( .A(n4624), .B(n4623), .Z(n4644) );
  XOR U5309 ( .A(n4645), .B(n4644), .Z(c[1152]) );
  NANDN U5310 ( .A(n4626), .B(n4625), .Z(n4630) );
  NAND U5311 ( .A(n4628), .B(n4627), .Z(n4629) );
  NAND U5312 ( .A(n4630), .B(n4629), .Z(n4663) );
  NANDN U5313 ( .A(n4632), .B(n4631), .Z(n4636) );
  OR U5314 ( .A(n4634), .B(n4633), .Z(n4635) );
  NAND U5315 ( .A(n4636), .B(n4635), .Z(n4660) );
  AND U5316 ( .A(b[2]), .B(a[131]), .Z(n4651) );
  AND U5317 ( .A(a[132]), .B(b[1]), .Z(n4649) );
  AND U5318 ( .A(a[130]), .B(b[3]), .Z(n4648) );
  XOR U5319 ( .A(n4649), .B(n4648), .Z(n4650) );
  XOR U5320 ( .A(n4651), .B(n4650), .Z(n4654) );
  NAND U5321 ( .A(b[0]), .B(a[133]), .Z(n4655) );
  XNOR U5322 ( .A(n4654), .B(n4655), .Z(n4656) );
  OR U5323 ( .A(n4638), .B(n4637), .Z(n4642) );
  NANDN U5324 ( .A(n4640), .B(n4639), .Z(n4641) );
  AND U5325 ( .A(n4642), .B(n4641), .Z(n4657) );
  XNOR U5326 ( .A(n4656), .B(n4657), .Z(n4661) );
  XNOR U5327 ( .A(n4660), .B(n4661), .Z(n4662) );
  XNOR U5328 ( .A(n4663), .B(n4662), .Z(n4666) );
  XNOR U5329 ( .A(sreg[1153]), .B(n4666), .Z(n4668) );
  NAND U5330 ( .A(n4643), .B(sreg[1152]), .Z(n4647) );
  OR U5331 ( .A(n4645), .B(n4644), .Z(n4646) );
  AND U5332 ( .A(n4647), .B(n4646), .Z(n4667) );
  XOR U5333 ( .A(n4668), .B(n4667), .Z(c[1153]) );
  AND U5334 ( .A(b[2]), .B(a[132]), .Z(n4680) );
  AND U5335 ( .A(a[133]), .B(b[1]), .Z(n4678) );
  AND U5336 ( .A(a[131]), .B(b[3]), .Z(n4677) );
  XOR U5337 ( .A(n4678), .B(n4677), .Z(n4679) );
  XOR U5338 ( .A(n4680), .B(n4679), .Z(n4683) );
  NAND U5339 ( .A(b[0]), .B(a[134]), .Z(n4684) );
  XOR U5340 ( .A(n4683), .B(n4684), .Z(n4686) );
  OR U5341 ( .A(n4649), .B(n4648), .Z(n4653) );
  NANDN U5342 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U5343 ( .A(n4653), .B(n4652), .Z(n4685) );
  XNOR U5344 ( .A(n4686), .B(n4685), .Z(n4671) );
  NANDN U5345 ( .A(n4655), .B(n4654), .Z(n4659) );
  NAND U5346 ( .A(n4657), .B(n4656), .Z(n4658) );
  NAND U5347 ( .A(n4659), .B(n4658), .Z(n4672) );
  XNOR U5348 ( .A(n4671), .B(n4672), .Z(n4673) );
  NANDN U5349 ( .A(n4661), .B(n4660), .Z(n4665) );
  NANDN U5350 ( .A(n4663), .B(n4662), .Z(n4664) );
  NAND U5351 ( .A(n4665), .B(n4664), .Z(n4674) );
  XOR U5352 ( .A(n4673), .B(n4674), .Z(n4689) );
  XNOR U5353 ( .A(n4689), .B(sreg[1154]), .Z(n4691) );
  NAND U5354 ( .A(sreg[1153]), .B(n4666), .Z(n4670) );
  OR U5355 ( .A(n4668), .B(n4667), .Z(n4669) );
  AND U5356 ( .A(n4670), .B(n4669), .Z(n4690) );
  XOR U5357 ( .A(n4691), .B(n4690), .Z(c[1154]) );
  NANDN U5358 ( .A(n4672), .B(n4671), .Z(n4676) );
  NANDN U5359 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U5360 ( .A(n4676), .B(n4675), .Z(n4712) );
  AND U5361 ( .A(b[2]), .B(a[133]), .Z(n4706) );
  AND U5362 ( .A(a[134]), .B(b[1]), .Z(n4704) );
  AND U5363 ( .A(a[132]), .B(b[3]), .Z(n4703) );
  XOR U5364 ( .A(n4704), .B(n4703), .Z(n4705) );
  XOR U5365 ( .A(n4706), .B(n4705), .Z(n4697) );
  NAND U5366 ( .A(b[0]), .B(a[135]), .Z(n4698) );
  XOR U5367 ( .A(n4697), .B(n4698), .Z(n4700) );
  OR U5368 ( .A(n4678), .B(n4677), .Z(n4682) );
  NANDN U5369 ( .A(n4680), .B(n4679), .Z(n4681) );
  NAND U5370 ( .A(n4682), .B(n4681), .Z(n4699) );
  XNOR U5371 ( .A(n4700), .B(n4699), .Z(n4709) );
  NANDN U5372 ( .A(n4684), .B(n4683), .Z(n4688) );
  OR U5373 ( .A(n4686), .B(n4685), .Z(n4687) );
  NAND U5374 ( .A(n4688), .B(n4687), .Z(n4710) );
  XNOR U5375 ( .A(n4709), .B(n4710), .Z(n4711) );
  XOR U5376 ( .A(n4712), .B(n4711), .Z(n4696) );
  NAND U5377 ( .A(n4689), .B(sreg[1154]), .Z(n4693) );
  OR U5378 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U5379 ( .A(n4693), .B(n4692), .Z(n4695) );
  XNOR U5380 ( .A(sreg[1155]), .B(n4695), .Z(n4694) );
  XOR U5381 ( .A(n4696), .B(n4694), .Z(c[1155]) );
  NANDN U5382 ( .A(n4698), .B(n4697), .Z(n4702) );
  OR U5383 ( .A(n4700), .B(n4699), .Z(n4701) );
  NAND U5384 ( .A(n4702), .B(n4701), .Z(n4715) );
  AND U5385 ( .A(b[2]), .B(a[134]), .Z(n4730) );
  AND U5386 ( .A(a[135]), .B(b[1]), .Z(n4728) );
  AND U5387 ( .A(a[133]), .B(b[3]), .Z(n4727) );
  XOR U5388 ( .A(n4728), .B(n4727), .Z(n4729) );
  XOR U5389 ( .A(n4730), .B(n4729), .Z(n4721) );
  NAND U5390 ( .A(b[0]), .B(a[136]), .Z(n4722) );
  XNOR U5391 ( .A(n4721), .B(n4722), .Z(n4723) );
  OR U5392 ( .A(n4704), .B(n4703), .Z(n4708) );
  NANDN U5393 ( .A(n4706), .B(n4705), .Z(n4707) );
  AND U5394 ( .A(n4708), .B(n4707), .Z(n4724) );
  XNOR U5395 ( .A(n4723), .B(n4724), .Z(n4716) );
  XNOR U5396 ( .A(n4715), .B(n4716), .Z(n4717) );
  NANDN U5397 ( .A(n4710), .B(n4709), .Z(n4714) );
  NAND U5398 ( .A(n4712), .B(n4711), .Z(n4713) );
  NAND U5399 ( .A(n4714), .B(n4713), .Z(n4718) );
  XOR U5400 ( .A(n4717), .B(n4718), .Z(n4733) );
  XNOR U5401 ( .A(sreg[1156]), .B(n4733), .Z(n4734) );
  XNOR U5402 ( .A(n4735), .B(n4734), .Z(c[1156]) );
  NANDN U5403 ( .A(n4716), .B(n4715), .Z(n4720) );
  NANDN U5404 ( .A(n4718), .B(n4717), .Z(n4719) );
  NAND U5405 ( .A(n4720), .B(n4719), .Z(n4756) );
  NANDN U5406 ( .A(n4722), .B(n4721), .Z(n4726) );
  NAND U5407 ( .A(n4724), .B(n4723), .Z(n4725) );
  NAND U5408 ( .A(n4726), .B(n4725), .Z(n4753) );
  AND U5409 ( .A(b[2]), .B(a[135]), .Z(n4744) );
  AND U5410 ( .A(a[136]), .B(b[1]), .Z(n4742) );
  AND U5411 ( .A(a[134]), .B(b[3]), .Z(n4741) );
  XOR U5412 ( .A(n4742), .B(n4741), .Z(n4743) );
  XOR U5413 ( .A(n4744), .B(n4743), .Z(n4747) );
  NAND U5414 ( .A(b[0]), .B(a[137]), .Z(n4748) );
  XNOR U5415 ( .A(n4747), .B(n4748), .Z(n4749) );
  OR U5416 ( .A(n4728), .B(n4727), .Z(n4732) );
  NANDN U5417 ( .A(n4730), .B(n4729), .Z(n4731) );
  AND U5418 ( .A(n4732), .B(n4731), .Z(n4750) );
  XNOR U5419 ( .A(n4749), .B(n4750), .Z(n4754) );
  XNOR U5420 ( .A(n4753), .B(n4754), .Z(n4755) );
  XOR U5421 ( .A(n4756), .B(n4755), .Z(n4740) );
  NANDN U5422 ( .A(sreg[1156]), .B(n4733), .Z(n4737) );
  NAND U5423 ( .A(n4735), .B(n4734), .Z(n4736) );
  AND U5424 ( .A(n4737), .B(n4736), .Z(n4739) );
  XOR U5425 ( .A(sreg[1157]), .B(n4739), .Z(n4738) );
  XOR U5426 ( .A(n4740), .B(n4738), .Z(c[1157]) );
  AND U5427 ( .A(b[2]), .B(a[136]), .Z(n4773) );
  AND U5428 ( .A(a[137]), .B(b[1]), .Z(n4771) );
  AND U5429 ( .A(a[135]), .B(b[3]), .Z(n4770) );
  XOR U5430 ( .A(n4771), .B(n4770), .Z(n4772) );
  XOR U5431 ( .A(n4773), .B(n4772), .Z(n4764) );
  NAND U5432 ( .A(b[0]), .B(a[138]), .Z(n4765) );
  XOR U5433 ( .A(n4764), .B(n4765), .Z(n4767) );
  OR U5434 ( .A(n4742), .B(n4741), .Z(n4746) );
  NANDN U5435 ( .A(n4744), .B(n4743), .Z(n4745) );
  NAND U5436 ( .A(n4746), .B(n4745), .Z(n4766) );
  XNOR U5437 ( .A(n4767), .B(n4766), .Z(n4776) );
  NANDN U5438 ( .A(n4748), .B(n4747), .Z(n4752) );
  NAND U5439 ( .A(n4750), .B(n4749), .Z(n4751) );
  NAND U5440 ( .A(n4752), .B(n4751), .Z(n4777) );
  XNOR U5441 ( .A(n4776), .B(n4777), .Z(n4778) );
  NANDN U5442 ( .A(n4754), .B(n4753), .Z(n4758) );
  NAND U5443 ( .A(n4756), .B(n4755), .Z(n4757) );
  NAND U5444 ( .A(n4758), .B(n4757), .Z(n4779) );
  XOR U5445 ( .A(n4778), .B(n4779), .Z(n4759) );
  XNOR U5446 ( .A(n4759), .B(sreg[1158]), .Z(n4761) );
  XNOR U5447 ( .A(n4760), .B(n4761), .Z(c[1158]) );
  NAND U5448 ( .A(n4759), .B(sreg[1158]), .Z(n4763) );
  NANDN U5449 ( .A(n4761), .B(n4760), .Z(n4762) );
  NAND U5450 ( .A(n4763), .B(n4762), .Z(n4783) );
  NANDN U5451 ( .A(n4765), .B(n4764), .Z(n4769) );
  OR U5452 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U5453 ( .A(n4769), .B(n4768), .Z(n4785) );
  AND U5454 ( .A(b[2]), .B(a[137]), .Z(n4800) );
  AND U5455 ( .A(a[138]), .B(b[1]), .Z(n4798) );
  AND U5456 ( .A(a[136]), .B(b[3]), .Z(n4797) );
  XOR U5457 ( .A(n4798), .B(n4797), .Z(n4799) );
  XOR U5458 ( .A(n4800), .B(n4799), .Z(n4791) );
  NAND U5459 ( .A(b[0]), .B(a[139]), .Z(n4792) );
  XNOR U5460 ( .A(n4791), .B(n4792), .Z(n4793) );
  OR U5461 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U5462 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U5463 ( .A(n4775), .B(n4774), .Z(n4794) );
  XNOR U5464 ( .A(n4793), .B(n4794), .Z(n4786) );
  XNOR U5465 ( .A(n4785), .B(n4786), .Z(n4787) );
  NANDN U5466 ( .A(n4777), .B(n4776), .Z(n4781) );
  NANDN U5467 ( .A(n4779), .B(n4778), .Z(n4780) );
  AND U5468 ( .A(n4781), .B(n4780), .Z(n4788) );
  XNOR U5469 ( .A(n4787), .B(n4788), .Z(n4784) );
  XOR U5470 ( .A(sreg[1159]), .B(n4784), .Z(n4782) );
  XNOR U5471 ( .A(n4783), .B(n4782), .Z(c[1159]) );
  NANDN U5472 ( .A(n4786), .B(n4785), .Z(n4790) );
  NAND U5473 ( .A(n4788), .B(n4787), .Z(n4789) );
  NAND U5474 ( .A(n4790), .B(n4789), .Z(n4818) );
  NANDN U5475 ( .A(n4792), .B(n4791), .Z(n4796) );
  NAND U5476 ( .A(n4794), .B(n4793), .Z(n4795) );
  NAND U5477 ( .A(n4796), .B(n4795), .Z(n4815) );
  AND U5478 ( .A(b[2]), .B(a[138]), .Z(n4806) );
  AND U5479 ( .A(a[139]), .B(b[1]), .Z(n4804) );
  AND U5480 ( .A(a[137]), .B(b[3]), .Z(n4803) );
  XOR U5481 ( .A(n4804), .B(n4803), .Z(n4805) );
  XOR U5482 ( .A(n4806), .B(n4805), .Z(n4809) );
  NAND U5483 ( .A(b[0]), .B(a[140]), .Z(n4810) );
  XNOR U5484 ( .A(n4809), .B(n4810), .Z(n4811) );
  OR U5485 ( .A(n4798), .B(n4797), .Z(n4802) );
  NANDN U5486 ( .A(n4800), .B(n4799), .Z(n4801) );
  AND U5487 ( .A(n4802), .B(n4801), .Z(n4812) );
  XNOR U5488 ( .A(n4811), .B(n4812), .Z(n4816) );
  XNOR U5489 ( .A(n4815), .B(n4816), .Z(n4817) );
  XOR U5490 ( .A(n4818), .B(n4817), .Z(n4821) );
  XNOR U5491 ( .A(sreg[1160]), .B(n4821), .Z(n4822) );
  XOR U5492 ( .A(n4823), .B(n4822), .Z(c[1160]) );
  AND U5493 ( .A(b[2]), .B(a[139]), .Z(n4835) );
  AND U5494 ( .A(a[140]), .B(b[1]), .Z(n4833) );
  AND U5495 ( .A(a[138]), .B(b[3]), .Z(n4832) );
  XOR U5496 ( .A(n4833), .B(n4832), .Z(n4834) );
  XOR U5497 ( .A(n4835), .B(n4834), .Z(n4826) );
  NAND U5498 ( .A(b[0]), .B(a[141]), .Z(n4827) );
  XOR U5499 ( .A(n4826), .B(n4827), .Z(n4829) );
  OR U5500 ( .A(n4804), .B(n4803), .Z(n4808) );
  NANDN U5501 ( .A(n4806), .B(n4805), .Z(n4807) );
  NAND U5502 ( .A(n4808), .B(n4807), .Z(n4828) );
  XNOR U5503 ( .A(n4829), .B(n4828), .Z(n4838) );
  NANDN U5504 ( .A(n4810), .B(n4809), .Z(n4814) );
  NAND U5505 ( .A(n4812), .B(n4811), .Z(n4813) );
  NAND U5506 ( .A(n4814), .B(n4813), .Z(n4839) );
  XNOR U5507 ( .A(n4838), .B(n4839), .Z(n4840) );
  NANDN U5508 ( .A(n4816), .B(n4815), .Z(n4820) );
  NAND U5509 ( .A(n4818), .B(n4817), .Z(n4819) );
  NAND U5510 ( .A(n4820), .B(n4819), .Z(n4841) );
  XOR U5511 ( .A(n4840), .B(n4841), .Z(n4844) );
  XNOR U5512 ( .A(n4844), .B(sreg[1161]), .Z(n4846) );
  NAND U5513 ( .A(sreg[1160]), .B(n4821), .Z(n4825) );
  OR U5514 ( .A(n4823), .B(n4822), .Z(n4824) );
  AND U5515 ( .A(n4825), .B(n4824), .Z(n4845) );
  XOR U5516 ( .A(n4846), .B(n4845), .Z(c[1161]) );
  NANDN U5517 ( .A(n4827), .B(n4826), .Z(n4831) );
  OR U5518 ( .A(n4829), .B(n4828), .Z(n4830) );
  NAND U5519 ( .A(n4831), .B(n4830), .Z(n4852) );
  AND U5520 ( .A(b[2]), .B(a[140]), .Z(n4861) );
  AND U5521 ( .A(a[141]), .B(b[1]), .Z(n4859) );
  AND U5522 ( .A(a[139]), .B(b[3]), .Z(n4858) );
  XOR U5523 ( .A(n4859), .B(n4858), .Z(n4860) );
  XOR U5524 ( .A(n4861), .B(n4860), .Z(n4864) );
  NAND U5525 ( .A(b[0]), .B(a[142]), .Z(n4865) );
  XNOR U5526 ( .A(n4864), .B(n4865), .Z(n4866) );
  OR U5527 ( .A(n4833), .B(n4832), .Z(n4837) );
  NANDN U5528 ( .A(n4835), .B(n4834), .Z(n4836) );
  AND U5529 ( .A(n4837), .B(n4836), .Z(n4867) );
  XNOR U5530 ( .A(n4866), .B(n4867), .Z(n4853) );
  XNOR U5531 ( .A(n4852), .B(n4853), .Z(n4854) );
  NANDN U5532 ( .A(n4839), .B(n4838), .Z(n4843) );
  NANDN U5533 ( .A(n4841), .B(n4840), .Z(n4842) );
  NAND U5534 ( .A(n4843), .B(n4842), .Z(n4855) );
  XOR U5535 ( .A(n4854), .B(n4855), .Z(n4851) );
  NAND U5536 ( .A(n4844), .B(sreg[1161]), .Z(n4848) );
  OR U5537 ( .A(n4846), .B(n4845), .Z(n4847) );
  AND U5538 ( .A(n4848), .B(n4847), .Z(n4850) );
  XNOR U5539 ( .A(n4850), .B(sreg[1162]), .Z(n4849) );
  XNOR U5540 ( .A(n4851), .B(n4849), .Z(c[1162]) );
  NANDN U5541 ( .A(n4853), .B(n4852), .Z(n4857) );
  NANDN U5542 ( .A(n4855), .B(n4854), .Z(n4856) );
  NAND U5543 ( .A(n4857), .B(n4856), .Z(n4885) );
  AND U5544 ( .A(b[2]), .B(a[141]), .Z(n4879) );
  AND U5545 ( .A(a[142]), .B(b[1]), .Z(n4877) );
  AND U5546 ( .A(a[140]), .B(b[3]), .Z(n4876) );
  XOR U5547 ( .A(n4877), .B(n4876), .Z(n4878) );
  XOR U5548 ( .A(n4879), .B(n4878), .Z(n4870) );
  NAND U5549 ( .A(b[0]), .B(a[143]), .Z(n4871) );
  XOR U5550 ( .A(n4870), .B(n4871), .Z(n4873) );
  OR U5551 ( .A(n4859), .B(n4858), .Z(n4863) );
  NANDN U5552 ( .A(n4861), .B(n4860), .Z(n4862) );
  NAND U5553 ( .A(n4863), .B(n4862), .Z(n4872) );
  XNOR U5554 ( .A(n4873), .B(n4872), .Z(n4882) );
  NANDN U5555 ( .A(n4865), .B(n4864), .Z(n4869) );
  NAND U5556 ( .A(n4867), .B(n4866), .Z(n4868) );
  NAND U5557 ( .A(n4869), .B(n4868), .Z(n4883) );
  XNOR U5558 ( .A(n4882), .B(n4883), .Z(n4884) );
  XOR U5559 ( .A(n4885), .B(n4884), .Z(n4888) );
  XNOR U5560 ( .A(n4888), .B(sreg[1163]), .Z(n4890) );
  XNOR U5561 ( .A(n4889), .B(n4890), .Z(c[1163]) );
  NANDN U5562 ( .A(n4871), .B(n4870), .Z(n4875) );
  OR U5563 ( .A(n4873), .B(n4872), .Z(n4874) );
  NAND U5564 ( .A(n4875), .B(n4874), .Z(n4893) );
  AND U5565 ( .A(b[2]), .B(a[142]), .Z(n4908) );
  AND U5566 ( .A(a[143]), .B(b[1]), .Z(n4906) );
  AND U5567 ( .A(a[141]), .B(b[3]), .Z(n4905) );
  XOR U5568 ( .A(n4906), .B(n4905), .Z(n4907) );
  XOR U5569 ( .A(n4908), .B(n4907), .Z(n4899) );
  NAND U5570 ( .A(b[0]), .B(a[144]), .Z(n4900) );
  XNOR U5571 ( .A(n4899), .B(n4900), .Z(n4901) );
  OR U5572 ( .A(n4877), .B(n4876), .Z(n4881) );
  NANDN U5573 ( .A(n4879), .B(n4878), .Z(n4880) );
  AND U5574 ( .A(n4881), .B(n4880), .Z(n4902) );
  XNOR U5575 ( .A(n4901), .B(n4902), .Z(n4894) );
  XNOR U5576 ( .A(n4893), .B(n4894), .Z(n4895) );
  NANDN U5577 ( .A(n4883), .B(n4882), .Z(n4887) );
  NANDN U5578 ( .A(n4885), .B(n4884), .Z(n4886) );
  AND U5579 ( .A(n4887), .B(n4886), .Z(n4896) );
  XOR U5580 ( .A(n4895), .B(n4896), .Z(n4911) );
  XNOR U5581 ( .A(sreg[1164]), .B(n4911), .Z(n4913) );
  NAND U5582 ( .A(n4888), .B(sreg[1163]), .Z(n4892) );
  NANDN U5583 ( .A(n4890), .B(n4889), .Z(n4891) );
  AND U5584 ( .A(n4892), .B(n4891), .Z(n4912) );
  XOR U5585 ( .A(n4913), .B(n4912), .Z(c[1164]) );
  NANDN U5586 ( .A(n4894), .B(n4893), .Z(n4898) );
  NAND U5587 ( .A(n4896), .B(n4895), .Z(n4897) );
  NAND U5588 ( .A(n4898), .B(n4897), .Z(n4919) );
  NANDN U5589 ( .A(n4900), .B(n4899), .Z(n4904) );
  NAND U5590 ( .A(n4902), .B(n4901), .Z(n4903) );
  NAND U5591 ( .A(n4904), .B(n4903), .Z(n4916) );
  AND U5592 ( .A(b[2]), .B(a[143]), .Z(n4925) );
  AND U5593 ( .A(a[144]), .B(b[1]), .Z(n4923) );
  AND U5594 ( .A(a[142]), .B(b[3]), .Z(n4922) );
  XOR U5595 ( .A(n4923), .B(n4922), .Z(n4924) );
  XOR U5596 ( .A(n4925), .B(n4924), .Z(n4928) );
  NAND U5597 ( .A(b[0]), .B(a[145]), .Z(n4929) );
  XNOR U5598 ( .A(n4928), .B(n4929), .Z(n4930) );
  OR U5599 ( .A(n4906), .B(n4905), .Z(n4910) );
  NANDN U5600 ( .A(n4908), .B(n4907), .Z(n4909) );
  AND U5601 ( .A(n4910), .B(n4909), .Z(n4931) );
  XNOR U5602 ( .A(n4930), .B(n4931), .Z(n4917) );
  XNOR U5603 ( .A(n4916), .B(n4917), .Z(n4918) );
  XOR U5604 ( .A(n4919), .B(n4918), .Z(n4934) );
  XOR U5605 ( .A(sreg[1165]), .B(n4934), .Z(n4935) );
  NAND U5606 ( .A(sreg[1164]), .B(n4911), .Z(n4915) );
  OR U5607 ( .A(n4913), .B(n4912), .Z(n4914) );
  NAND U5608 ( .A(n4915), .B(n4914), .Z(n4936) );
  XOR U5609 ( .A(n4935), .B(n4936), .Z(c[1165]) );
  NANDN U5610 ( .A(n4917), .B(n4916), .Z(n4921) );
  NAND U5611 ( .A(n4919), .B(n4918), .Z(n4920) );
  NAND U5612 ( .A(n4921), .B(n4920), .Z(n4943) );
  AND U5613 ( .A(b[2]), .B(a[144]), .Z(n4949) );
  AND U5614 ( .A(a[145]), .B(b[1]), .Z(n4947) );
  AND U5615 ( .A(a[143]), .B(b[3]), .Z(n4946) );
  XOR U5616 ( .A(n4947), .B(n4946), .Z(n4948) );
  XOR U5617 ( .A(n4949), .B(n4948), .Z(n4952) );
  NAND U5618 ( .A(b[0]), .B(a[146]), .Z(n4953) );
  XOR U5619 ( .A(n4952), .B(n4953), .Z(n4955) );
  OR U5620 ( .A(n4923), .B(n4922), .Z(n4927) );
  NANDN U5621 ( .A(n4925), .B(n4924), .Z(n4926) );
  NAND U5622 ( .A(n4927), .B(n4926), .Z(n4954) );
  XNOR U5623 ( .A(n4955), .B(n4954), .Z(n4940) );
  NANDN U5624 ( .A(n4929), .B(n4928), .Z(n4933) );
  NAND U5625 ( .A(n4931), .B(n4930), .Z(n4932) );
  NAND U5626 ( .A(n4933), .B(n4932), .Z(n4941) );
  XNOR U5627 ( .A(n4940), .B(n4941), .Z(n4942) );
  XOR U5628 ( .A(n4943), .B(n4942), .Z(n4959) );
  OR U5629 ( .A(n4934), .B(sreg[1165]), .Z(n4938) );
  NANDN U5630 ( .A(n4936), .B(n4935), .Z(n4937) );
  AND U5631 ( .A(n4938), .B(n4937), .Z(n4958) );
  XNOR U5632 ( .A(sreg[1166]), .B(n4958), .Z(n4939) );
  XNOR U5633 ( .A(n4959), .B(n4939), .Z(c[1166]) );
  NANDN U5634 ( .A(n4941), .B(n4940), .Z(n4945) );
  NANDN U5635 ( .A(n4943), .B(n4942), .Z(n4944) );
  NAND U5636 ( .A(n4945), .B(n4944), .Z(n4966) );
  AND U5637 ( .A(b[2]), .B(a[145]), .Z(n4972) );
  AND U5638 ( .A(a[146]), .B(b[1]), .Z(n4970) );
  AND U5639 ( .A(a[144]), .B(b[3]), .Z(n4969) );
  XOR U5640 ( .A(n4970), .B(n4969), .Z(n4971) );
  XOR U5641 ( .A(n4972), .B(n4971), .Z(n4975) );
  NAND U5642 ( .A(b[0]), .B(a[147]), .Z(n4976) );
  XOR U5643 ( .A(n4975), .B(n4976), .Z(n4978) );
  OR U5644 ( .A(n4947), .B(n4946), .Z(n4951) );
  NANDN U5645 ( .A(n4949), .B(n4948), .Z(n4950) );
  NAND U5646 ( .A(n4951), .B(n4950), .Z(n4977) );
  XNOR U5647 ( .A(n4978), .B(n4977), .Z(n4963) );
  NANDN U5648 ( .A(n4953), .B(n4952), .Z(n4957) );
  OR U5649 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U5650 ( .A(n4957), .B(n4956), .Z(n4964) );
  XNOR U5651 ( .A(n4963), .B(n4964), .Z(n4965) );
  XNOR U5652 ( .A(n4966), .B(n4965), .Z(n4962) );
  XOR U5653 ( .A(n4961), .B(sreg[1167]), .Z(n4960) );
  XOR U5654 ( .A(n4962), .B(n4960), .Z(c[1167]) );
  NANDN U5655 ( .A(n4964), .B(n4963), .Z(n4968) );
  NAND U5656 ( .A(n4966), .B(n4965), .Z(n4967) );
  NAND U5657 ( .A(n4968), .B(n4967), .Z(n4984) );
  AND U5658 ( .A(b[2]), .B(a[146]), .Z(n4990) );
  AND U5659 ( .A(a[147]), .B(b[1]), .Z(n4988) );
  AND U5660 ( .A(a[145]), .B(b[3]), .Z(n4987) );
  XOR U5661 ( .A(n4988), .B(n4987), .Z(n4989) );
  XOR U5662 ( .A(n4990), .B(n4989), .Z(n4993) );
  NAND U5663 ( .A(b[0]), .B(a[148]), .Z(n4994) );
  XOR U5664 ( .A(n4993), .B(n4994), .Z(n4996) );
  OR U5665 ( .A(n4970), .B(n4969), .Z(n4974) );
  NANDN U5666 ( .A(n4972), .B(n4971), .Z(n4973) );
  NAND U5667 ( .A(n4974), .B(n4973), .Z(n4995) );
  XNOR U5668 ( .A(n4996), .B(n4995), .Z(n4981) );
  NANDN U5669 ( .A(n4976), .B(n4975), .Z(n4980) );
  OR U5670 ( .A(n4978), .B(n4977), .Z(n4979) );
  NAND U5671 ( .A(n4980), .B(n4979), .Z(n4982) );
  XNOR U5672 ( .A(n4981), .B(n4982), .Z(n4983) );
  XNOR U5673 ( .A(n4984), .B(n4983), .Z(n4999) );
  XNOR U5674 ( .A(n4999), .B(sreg[1168]), .Z(n5001) );
  XNOR U5675 ( .A(n5000), .B(n5001), .Z(c[1168]) );
  NANDN U5676 ( .A(n4982), .B(n4981), .Z(n4986) );
  NAND U5677 ( .A(n4984), .B(n4983), .Z(n4985) );
  NAND U5678 ( .A(n4986), .B(n4985), .Z(n5007) );
  AND U5679 ( .A(b[2]), .B(a[147]), .Z(n5013) );
  AND U5680 ( .A(a[148]), .B(b[1]), .Z(n5011) );
  AND U5681 ( .A(a[146]), .B(b[3]), .Z(n5010) );
  XOR U5682 ( .A(n5011), .B(n5010), .Z(n5012) );
  XOR U5683 ( .A(n5013), .B(n5012), .Z(n5016) );
  NAND U5684 ( .A(b[0]), .B(a[149]), .Z(n5017) );
  XOR U5685 ( .A(n5016), .B(n5017), .Z(n5019) );
  OR U5686 ( .A(n4988), .B(n4987), .Z(n4992) );
  NANDN U5687 ( .A(n4990), .B(n4989), .Z(n4991) );
  NAND U5688 ( .A(n4992), .B(n4991), .Z(n5018) );
  XNOR U5689 ( .A(n5019), .B(n5018), .Z(n5004) );
  NANDN U5690 ( .A(n4994), .B(n4993), .Z(n4998) );
  OR U5691 ( .A(n4996), .B(n4995), .Z(n4997) );
  NAND U5692 ( .A(n4998), .B(n4997), .Z(n5005) );
  XNOR U5693 ( .A(n5004), .B(n5005), .Z(n5006) );
  XNOR U5694 ( .A(n5007), .B(n5006), .Z(n5022) );
  XNOR U5695 ( .A(n5022), .B(sreg[1169]), .Z(n5024) );
  NAND U5696 ( .A(n4999), .B(sreg[1168]), .Z(n5003) );
  NANDN U5697 ( .A(n5001), .B(n5000), .Z(n5002) );
  AND U5698 ( .A(n5003), .B(n5002), .Z(n5023) );
  XOR U5699 ( .A(n5024), .B(n5023), .Z(c[1169]) );
  NANDN U5700 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U5701 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U5702 ( .A(n5009), .B(n5008), .Z(n5033) );
  AND U5703 ( .A(b[2]), .B(a[148]), .Z(n5039) );
  AND U5704 ( .A(a[149]), .B(b[1]), .Z(n5037) );
  AND U5705 ( .A(a[147]), .B(b[3]), .Z(n5036) );
  XOR U5706 ( .A(n5037), .B(n5036), .Z(n5038) );
  XOR U5707 ( .A(n5039), .B(n5038), .Z(n5042) );
  NAND U5708 ( .A(b[0]), .B(a[150]), .Z(n5043) );
  XOR U5709 ( .A(n5042), .B(n5043), .Z(n5045) );
  OR U5710 ( .A(n5011), .B(n5010), .Z(n5015) );
  NANDN U5711 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U5712 ( .A(n5015), .B(n5014), .Z(n5044) );
  XNOR U5713 ( .A(n5045), .B(n5044), .Z(n5030) );
  NANDN U5714 ( .A(n5017), .B(n5016), .Z(n5021) );
  OR U5715 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U5716 ( .A(n5021), .B(n5020), .Z(n5031) );
  XNOR U5717 ( .A(n5030), .B(n5031), .Z(n5032) );
  XNOR U5718 ( .A(n5033), .B(n5032), .Z(n5029) );
  NAND U5719 ( .A(n5022), .B(sreg[1169]), .Z(n5026) );
  OR U5720 ( .A(n5024), .B(n5023), .Z(n5025) );
  AND U5721 ( .A(n5026), .B(n5025), .Z(n5028) );
  XNOR U5722 ( .A(n5028), .B(sreg[1170]), .Z(n5027) );
  XOR U5723 ( .A(n5029), .B(n5027), .Z(c[1170]) );
  NANDN U5724 ( .A(n5031), .B(n5030), .Z(n5035) );
  NAND U5725 ( .A(n5033), .B(n5032), .Z(n5034) );
  NAND U5726 ( .A(n5035), .B(n5034), .Z(n5051) );
  AND U5727 ( .A(b[2]), .B(a[149]), .Z(n5057) );
  AND U5728 ( .A(a[150]), .B(b[1]), .Z(n5055) );
  AND U5729 ( .A(a[148]), .B(b[3]), .Z(n5054) );
  XOR U5730 ( .A(n5055), .B(n5054), .Z(n5056) );
  XOR U5731 ( .A(n5057), .B(n5056), .Z(n5060) );
  NAND U5732 ( .A(b[0]), .B(a[151]), .Z(n5061) );
  XOR U5733 ( .A(n5060), .B(n5061), .Z(n5063) );
  OR U5734 ( .A(n5037), .B(n5036), .Z(n5041) );
  NANDN U5735 ( .A(n5039), .B(n5038), .Z(n5040) );
  NAND U5736 ( .A(n5041), .B(n5040), .Z(n5062) );
  XNOR U5737 ( .A(n5063), .B(n5062), .Z(n5048) );
  NANDN U5738 ( .A(n5043), .B(n5042), .Z(n5047) );
  OR U5739 ( .A(n5045), .B(n5044), .Z(n5046) );
  NAND U5740 ( .A(n5047), .B(n5046), .Z(n5049) );
  XNOR U5741 ( .A(n5048), .B(n5049), .Z(n5050) );
  XNOR U5742 ( .A(n5051), .B(n5050), .Z(n5066) );
  XNOR U5743 ( .A(n5066), .B(sreg[1171]), .Z(n5068) );
  XNOR U5744 ( .A(n5067), .B(n5068), .Z(c[1171]) );
  NANDN U5745 ( .A(n5049), .B(n5048), .Z(n5053) );
  NAND U5746 ( .A(n5051), .B(n5050), .Z(n5052) );
  NAND U5747 ( .A(n5053), .B(n5052), .Z(n5075) );
  AND U5748 ( .A(b[2]), .B(a[150]), .Z(n5081) );
  AND U5749 ( .A(a[151]), .B(b[1]), .Z(n5079) );
  AND U5750 ( .A(a[149]), .B(b[3]), .Z(n5078) );
  XOR U5751 ( .A(n5079), .B(n5078), .Z(n5080) );
  XOR U5752 ( .A(n5081), .B(n5080), .Z(n5084) );
  NAND U5753 ( .A(b[0]), .B(a[152]), .Z(n5085) );
  XOR U5754 ( .A(n5084), .B(n5085), .Z(n5087) );
  OR U5755 ( .A(n5055), .B(n5054), .Z(n5059) );
  NANDN U5756 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U5757 ( .A(n5059), .B(n5058), .Z(n5086) );
  XNOR U5758 ( .A(n5087), .B(n5086), .Z(n5072) );
  NANDN U5759 ( .A(n5061), .B(n5060), .Z(n5065) );
  OR U5760 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U5761 ( .A(n5065), .B(n5064), .Z(n5073) );
  XNOR U5762 ( .A(n5072), .B(n5073), .Z(n5074) );
  XNOR U5763 ( .A(n5075), .B(n5074), .Z(n5091) );
  NAND U5764 ( .A(n5066), .B(sreg[1171]), .Z(n5070) );
  NANDN U5765 ( .A(n5068), .B(n5067), .Z(n5069) );
  AND U5766 ( .A(n5070), .B(n5069), .Z(n5090) );
  XNOR U5767 ( .A(n5090), .B(sreg[1172]), .Z(n5071) );
  XOR U5768 ( .A(n5091), .B(n5071), .Z(c[1172]) );
  NANDN U5769 ( .A(n5073), .B(n5072), .Z(n5077) );
  NAND U5770 ( .A(n5075), .B(n5074), .Z(n5076) );
  NAND U5771 ( .A(n5077), .B(n5076), .Z(n5098) );
  AND U5772 ( .A(b[2]), .B(a[151]), .Z(n5104) );
  AND U5773 ( .A(a[152]), .B(b[1]), .Z(n5102) );
  AND U5774 ( .A(a[150]), .B(b[3]), .Z(n5101) );
  XOR U5775 ( .A(n5102), .B(n5101), .Z(n5103) );
  XOR U5776 ( .A(n5104), .B(n5103), .Z(n5107) );
  NAND U5777 ( .A(b[0]), .B(a[153]), .Z(n5108) );
  XOR U5778 ( .A(n5107), .B(n5108), .Z(n5110) );
  OR U5779 ( .A(n5079), .B(n5078), .Z(n5083) );
  NANDN U5780 ( .A(n5081), .B(n5080), .Z(n5082) );
  NAND U5781 ( .A(n5083), .B(n5082), .Z(n5109) );
  XNOR U5782 ( .A(n5110), .B(n5109), .Z(n5095) );
  NANDN U5783 ( .A(n5085), .B(n5084), .Z(n5089) );
  OR U5784 ( .A(n5087), .B(n5086), .Z(n5088) );
  NAND U5785 ( .A(n5089), .B(n5088), .Z(n5096) );
  XNOR U5786 ( .A(n5095), .B(n5096), .Z(n5097) );
  XNOR U5787 ( .A(n5098), .B(n5097), .Z(n5094) );
  XOR U5788 ( .A(n5093), .B(sreg[1173]), .Z(n5092) );
  XOR U5789 ( .A(n5094), .B(n5092), .Z(c[1173]) );
  NANDN U5790 ( .A(n5096), .B(n5095), .Z(n5100) );
  NAND U5791 ( .A(n5098), .B(n5097), .Z(n5099) );
  NAND U5792 ( .A(n5100), .B(n5099), .Z(n5121) );
  AND U5793 ( .A(b[2]), .B(a[152]), .Z(n5127) );
  AND U5794 ( .A(a[153]), .B(b[1]), .Z(n5125) );
  AND U5795 ( .A(a[151]), .B(b[3]), .Z(n5124) );
  XOR U5796 ( .A(n5125), .B(n5124), .Z(n5126) );
  XOR U5797 ( .A(n5127), .B(n5126), .Z(n5130) );
  NAND U5798 ( .A(b[0]), .B(a[154]), .Z(n5131) );
  XOR U5799 ( .A(n5130), .B(n5131), .Z(n5133) );
  OR U5800 ( .A(n5102), .B(n5101), .Z(n5106) );
  NANDN U5801 ( .A(n5104), .B(n5103), .Z(n5105) );
  NAND U5802 ( .A(n5106), .B(n5105), .Z(n5132) );
  XNOR U5803 ( .A(n5133), .B(n5132), .Z(n5118) );
  NANDN U5804 ( .A(n5108), .B(n5107), .Z(n5112) );
  OR U5805 ( .A(n5110), .B(n5109), .Z(n5111) );
  NAND U5806 ( .A(n5112), .B(n5111), .Z(n5119) );
  XNOR U5807 ( .A(n5118), .B(n5119), .Z(n5120) );
  XNOR U5808 ( .A(n5121), .B(n5120), .Z(n5113) );
  XOR U5809 ( .A(sreg[1174]), .B(n5113), .Z(n5114) );
  XOR U5810 ( .A(n5115), .B(n5114), .Z(c[1174]) );
  OR U5811 ( .A(n5113), .B(sreg[1174]), .Z(n5117) );
  NANDN U5812 ( .A(n5115), .B(n5114), .Z(n5116) );
  NAND U5813 ( .A(n5117), .B(n5116), .Z(n5138) );
  NANDN U5814 ( .A(n5119), .B(n5118), .Z(n5123) );
  NAND U5815 ( .A(n5121), .B(n5120), .Z(n5122) );
  NAND U5816 ( .A(n5123), .B(n5122), .Z(n5144) );
  AND U5817 ( .A(b[2]), .B(a[153]), .Z(n5150) );
  AND U5818 ( .A(a[154]), .B(b[1]), .Z(n5148) );
  AND U5819 ( .A(a[152]), .B(b[3]), .Z(n5147) );
  XOR U5820 ( .A(n5148), .B(n5147), .Z(n5149) );
  XOR U5821 ( .A(n5150), .B(n5149), .Z(n5153) );
  NAND U5822 ( .A(b[0]), .B(a[155]), .Z(n5154) );
  XOR U5823 ( .A(n5153), .B(n5154), .Z(n5156) );
  OR U5824 ( .A(n5125), .B(n5124), .Z(n5129) );
  NANDN U5825 ( .A(n5127), .B(n5126), .Z(n5128) );
  NAND U5826 ( .A(n5129), .B(n5128), .Z(n5155) );
  XNOR U5827 ( .A(n5156), .B(n5155), .Z(n5141) );
  NANDN U5828 ( .A(n5131), .B(n5130), .Z(n5135) );
  OR U5829 ( .A(n5133), .B(n5132), .Z(n5134) );
  NAND U5830 ( .A(n5135), .B(n5134), .Z(n5142) );
  XNOR U5831 ( .A(n5141), .B(n5142), .Z(n5143) );
  XNOR U5832 ( .A(n5144), .B(n5143), .Z(n5136) );
  XNOR U5833 ( .A(n5136), .B(sreg[1175]), .Z(n5137) );
  XOR U5834 ( .A(n5138), .B(n5137), .Z(c[1175]) );
  NAND U5835 ( .A(n5136), .B(sreg[1175]), .Z(n5140) );
  OR U5836 ( .A(n5138), .B(n5137), .Z(n5139) );
  AND U5837 ( .A(n5140), .B(n5139), .Z(n5179) );
  NANDN U5838 ( .A(n5142), .B(n5141), .Z(n5146) );
  NAND U5839 ( .A(n5144), .B(n5143), .Z(n5145) );
  NAND U5840 ( .A(n5146), .B(n5145), .Z(n5163) );
  AND U5841 ( .A(b[2]), .B(a[154]), .Z(n5169) );
  AND U5842 ( .A(a[155]), .B(b[1]), .Z(n5167) );
  AND U5843 ( .A(a[153]), .B(b[3]), .Z(n5166) );
  XOR U5844 ( .A(n5167), .B(n5166), .Z(n5168) );
  XOR U5845 ( .A(n5169), .B(n5168), .Z(n5172) );
  NAND U5846 ( .A(b[0]), .B(a[156]), .Z(n5173) );
  XOR U5847 ( .A(n5172), .B(n5173), .Z(n5175) );
  OR U5848 ( .A(n5148), .B(n5147), .Z(n5152) );
  NANDN U5849 ( .A(n5150), .B(n5149), .Z(n5151) );
  NAND U5850 ( .A(n5152), .B(n5151), .Z(n5174) );
  XNOR U5851 ( .A(n5175), .B(n5174), .Z(n5160) );
  NANDN U5852 ( .A(n5154), .B(n5153), .Z(n5158) );
  OR U5853 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U5854 ( .A(n5158), .B(n5157), .Z(n5161) );
  XNOR U5855 ( .A(n5160), .B(n5161), .Z(n5162) );
  XNOR U5856 ( .A(n5163), .B(n5162), .Z(n5178) );
  XNOR U5857 ( .A(sreg[1176]), .B(n5178), .Z(n5159) );
  XOR U5858 ( .A(n5179), .B(n5159), .Z(c[1176]) );
  NANDN U5859 ( .A(n5161), .B(n5160), .Z(n5165) );
  NAND U5860 ( .A(n5163), .B(n5162), .Z(n5164) );
  NAND U5861 ( .A(n5165), .B(n5164), .Z(n5186) );
  AND U5862 ( .A(b[2]), .B(a[155]), .Z(n5192) );
  AND U5863 ( .A(a[156]), .B(b[1]), .Z(n5190) );
  AND U5864 ( .A(a[154]), .B(b[3]), .Z(n5189) );
  XOR U5865 ( .A(n5190), .B(n5189), .Z(n5191) );
  XOR U5866 ( .A(n5192), .B(n5191), .Z(n5195) );
  NAND U5867 ( .A(b[0]), .B(a[157]), .Z(n5196) );
  XOR U5868 ( .A(n5195), .B(n5196), .Z(n5198) );
  OR U5869 ( .A(n5167), .B(n5166), .Z(n5171) );
  NANDN U5870 ( .A(n5169), .B(n5168), .Z(n5170) );
  NAND U5871 ( .A(n5171), .B(n5170), .Z(n5197) );
  XNOR U5872 ( .A(n5198), .B(n5197), .Z(n5183) );
  NANDN U5873 ( .A(n5173), .B(n5172), .Z(n5177) );
  OR U5874 ( .A(n5175), .B(n5174), .Z(n5176) );
  NAND U5875 ( .A(n5177), .B(n5176), .Z(n5184) );
  XNOR U5876 ( .A(n5183), .B(n5184), .Z(n5185) );
  XNOR U5877 ( .A(n5186), .B(n5185), .Z(n5182) );
  XOR U5878 ( .A(n5181), .B(sreg[1177]), .Z(n5180) );
  XOR U5879 ( .A(n5182), .B(n5180), .Z(c[1177]) );
  NANDN U5880 ( .A(n5184), .B(n5183), .Z(n5188) );
  NAND U5881 ( .A(n5186), .B(n5185), .Z(n5187) );
  NAND U5882 ( .A(n5188), .B(n5187), .Z(n5204) );
  AND U5883 ( .A(b[2]), .B(a[156]), .Z(n5210) );
  AND U5884 ( .A(a[157]), .B(b[1]), .Z(n5208) );
  AND U5885 ( .A(a[155]), .B(b[3]), .Z(n5207) );
  XOR U5886 ( .A(n5208), .B(n5207), .Z(n5209) );
  XOR U5887 ( .A(n5210), .B(n5209), .Z(n5213) );
  NAND U5888 ( .A(b[0]), .B(a[158]), .Z(n5214) );
  XOR U5889 ( .A(n5213), .B(n5214), .Z(n5216) );
  OR U5890 ( .A(n5190), .B(n5189), .Z(n5194) );
  NANDN U5891 ( .A(n5192), .B(n5191), .Z(n5193) );
  NAND U5892 ( .A(n5194), .B(n5193), .Z(n5215) );
  XNOR U5893 ( .A(n5216), .B(n5215), .Z(n5201) );
  NANDN U5894 ( .A(n5196), .B(n5195), .Z(n5200) );
  OR U5895 ( .A(n5198), .B(n5197), .Z(n5199) );
  NAND U5896 ( .A(n5200), .B(n5199), .Z(n5202) );
  XNOR U5897 ( .A(n5201), .B(n5202), .Z(n5203) );
  XNOR U5898 ( .A(n5204), .B(n5203), .Z(n5219) );
  XNOR U5899 ( .A(n5219), .B(sreg[1178]), .Z(n5221) );
  XNOR U5900 ( .A(n5220), .B(n5221), .Z(c[1178]) );
  NANDN U5901 ( .A(n5202), .B(n5201), .Z(n5206) );
  NAND U5902 ( .A(n5204), .B(n5203), .Z(n5205) );
  NAND U5903 ( .A(n5206), .B(n5205), .Z(n5227) );
  AND U5904 ( .A(b[2]), .B(a[157]), .Z(n5233) );
  AND U5905 ( .A(a[158]), .B(b[1]), .Z(n5231) );
  AND U5906 ( .A(a[156]), .B(b[3]), .Z(n5230) );
  XOR U5907 ( .A(n5231), .B(n5230), .Z(n5232) );
  XOR U5908 ( .A(n5233), .B(n5232), .Z(n5236) );
  NAND U5909 ( .A(b[0]), .B(a[159]), .Z(n5237) );
  XOR U5910 ( .A(n5236), .B(n5237), .Z(n5239) );
  OR U5911 ( .A(n5208), .B(n5207), .Z(n5212) );
  NANDN U5912 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U5913 ( .A(n5212), .B(n5211), .Z(n5238) );
  XNOR U5914 ( .A(n5239), .B(n5238), .Z(n5224) );
  NANDN U5915 ( .A(n5214), .B(n5213), .Z(n5218) );
  OR U5916 ( .A(n5216), .B(n5215), .Z(n5217) );
  NAND U5917 ( .A(n5218), .B(n5217), .Z(n5225) );
  XNOR U5918 ( .A(n5224), .B(n5225), .Z(n5226) );
  XNOR U5919 ( .A(n5227), .B(n5226), .Z(n5242) );
  XOR U5920 ( .A(sreg[1179]), .B(n5242), .Z(n5243) );
  NAND U5921 ( .A(n5219), .B(sreg[1178]), .Z(n5223) );
  NANDN U5922 ( .A(n5221), .B(n5220), .Z(n5222) );
  NAND U5923 ( .A(n5223), .B(n5222), .Z(n5244) );
  XOR U5924 ( .A(n5243), .B(n5244), .Z(c[1179]) );
  NANDN U5925 ( .A(n5225), .B(n5224), .Z(n5229) );
  NAND U5926 ( .A(n5227), .B(n5226), .Z(n5228) );
  NAND U5927 ( .A(n5229), .B(n5228), .Z(n5253) );
  AND U5928 ( .A(b[2]), .B(a[158]), .Z(n5259) );
  AND U5929 ( .A(a[159]), .B(b[1]), .Z(n5257) );
  AND U5930 ( .A(a[157]), .B(b[3]), .Z(n5256) );
  XOR U5931 ( .A(n5257), .B(n5256), .Z(n5258) );
  XOR U5932 ( .A(n5259), .B(n5258), .Z(n5262) );
  NAND U5933 ( .A(b[0]), .B(a[160]), .Z(n5263) );
  XOR U5934 ( .A(n5262), .B(n5263), .Z(n5265) );
  OR U5935 ( .A(n5231), .B(n5230), .Z(n5235) );
  NANDN U5936 ( .A(n5233), .B(n5232), .Z(n5234) );
  NAND U5937 ( .A(n5235), .B(n5234), .Z(n5264) );
  XNOR U5938 ( .A(n5265), .B(n5264), .Z(n5250) );
  NANDN U5939 ( .A(n5237), .B(n5236), .Z(n5241) );
  OR U5940 ( .A(n5239), .B(n5238), .Z(n5240) );
  NAND U5941 ( .A(n5241), .B(n5240), .Z(n5251) );
  XNOR U5942 ( .A(n5250), .B(n5251), .Z(n5252) );
  XOR U5943 ( .A(n5253), .B(n5252), .Z(n5249) );
  OR U5944 ( .A(n5242), .B(sreg[1179]), .Z(n5246) );
  NANDN U5945 ( .A(n5244), .B(n5243), .Z(n5245) );
  AND U5946 ( .A(n5246), .B(n5245), .Z(n5248) );
  XNOR U5947 ( .A(sreg[1180]), .B(n5248), .Z(n5247) );
  XOR U5948 ( .A(n5249), .B(n5247), .Z(c[1180]) );
  NANDN U5949 ( .A(n5251), .B(n5250), .Z(n5255) );
  NAND U5950 ( .A(n5253), .B(n5252), .Z(n5254) );
  NAND U5951 ( .A(n5255), .B(n5254), .Z(n5271) );
  AND U5952 ( .A(b[2]), .B(a[159]), .Z(n5277) );
  AND U5953 ( .A(a[160]), .B(b[1]), .Z(n5275) );
  AND U5954 ( .A(a[158]), .B(b[3]), .Z(n5274) );
  XOR U5955 ( .A(n5275), .B(n5274), .Z(n5276) );
  XOR U5956 ( .A(n5277), .B(n5276), .Z(n5280) );
  NAND U5957 ( .A(b[0]), .B(a[161]), .Z(n5281) );
  XOR U5958 ( .A(n5280), .B(n5281), .Z(n5283) );
  OR U5959 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U5960 ( .A(n5259), .B(n5258), .Z(n5260) );
  NAND U5961 ( .A(n5261), .B(n5260), .Z(n5282) );
  XNOR U5962 ( .A(n5283), .B(n5282), .Z(n5268) );
  NANDN U5963 ( .A(n5263), .B(n5262), .Z(n5267) );
  OR U5964 ( .A(n5265), .B(n5264), .Z(n5266) );
  NAND U5965 ( .A(n5267), .B(n5266), .Z(n5269) );
  XNOR U5966 ( .A(n5268), .B(n5269), .Z(n5270) );
  XNOR U5967 ( .A(n5271), .B(n5270), .Z(n5286) );
  XNOR U5968 ( .A(n5286), .B(sreg[1181]), .Z(n5287) );
  XOR U5969 ( .A(n5288), .B(n5287), .Z(c[1181]) );
  NANDN U5970 ( .A(n5269), .B(n5268), .Z(n5273) );
  NAND U5971 ( .A(n5271), .B(n5270), .Z(n5272) );
  NAND U5972 ( .A(n5273), .B(n5272), .Z(n5297) );
  AND U5973 ( .A(b[2]), .B(a[160]), .Z(n5303) );
  AND U5974 ( .A(a[161]), .B(b[1]), .Z(n5301) );
  AND U5975 ( .A(a[159]), .B(b[3]), .Z(n5300) );
  XOR U5976 ( .A(n5301), .B(n5300), .Z(n5302) );
  XOR U5977 ( .A(n5303), .B(n5302), .Z(n5306) );
  NAND U5978 ( .A(b[0]), .B(a[162]), .Z(n5307) );
  XOR U5979 ( .A(n5306), .B(n5307), .Z(n5309) );
  OR U5980 ( .A(n5275), .B(n5274), .Z(n5279) );
  NANDN U5981 ( .A(n5277), .B(n5276), .Z(n5278) );
  NAND U5982 ( .A(n5279), .B(n5278), .Z(n5308) );
  XNOR U5983 ( .A(n5309), .B(n5308), .Z(n5294) );
  NANDN U5984 ( .A(n5281), .B(n5280), .Z(n5285) );
  OR U5985 ( .A(n5283), .B(n5282), .Z(n5284) );
  NAND U5986 ( .A(n5285), .B(n5284), .Z(n5295) );
  XNOR U5987 ( .A(n5294), .B(n5295), .Z(n5296) );
  XOR U5988 ( .A(n5297), .B(n5296), .Z(n5293) );
  NAND U5989 ( .A(n5286), .B(sreg[1181]), .Z(n5290) );
  OR U5990 ( .A(n5288), .B(n5287), .Z(n5289) );
  NAND U5991 ( .A(n5290), .B(n5289), .Z(n5292) );
  XNOR U5992 ( .A(sreg[1182]), .B(n5292), .Z(n5291) );
  XOR U5993 ( .A(n5293), .B(n5291), .Z(c[1182]) );
  NANDN U5994 ( .A(n5295), .B(n5294), .Z(n5299) );
  NAND U5995 ( .A(n5297), .B(n5296), .Z(n5298) );
  NAND U5996 ( .A(n5299), .B(n5298), .Z(n5315) );
  AND U5997 ( .A(b[2]), .B(a[161]), .Z(n5321) );
  AND U5998 ( .A(a[162]), .B(b[1]), .Z(n5319) );
  AND U5999 ( .A(a[160]), .B(b[3]), .Z(n5318) );
  XOR U6000 ( .A(n5319), .B(n5318), .Z(n5320) );
  XOR U6001 ( .A(n5321), .B(n5320), .Z(n5324) );
  NAND U6002 ( .A(b[0]), .B(a[163]), .Z(n5325) );
  XOR U6003 ( .A(n5324), .B(n5325), .Z(n5327) );
  OR U6004 ( .A(n5301), .B(n5300), .Z(n5305) );
  NANDN U6005 ( .A(n5303), .B(n5302), .Z(n5304) );
  NAND U6006 ( .A(n5305), .B(n5304), .Z(n5326) );
  XNOR U6007 ( .A(n5327), .B(n5326), .Z(n5312) );
  NANDN U6008 ( .A(n5307), .B(n5306), .Z(n5311) );
  OR U6009 ( .A(n5309), .B(n5308), .Z(n5310) );
  NAND U6010 ( .A(n5311), .B(n5310), .Z(n5313) );
  XNOR U6011 ( .A(n5312), .B(n5313), .Z(n5314) );
  XNOR U6012 ( .A(n5315), .B(n5314), .Z(n5330) );
  XNOR U6013 ( .A(n5330), .B(sreg[1183]), .Z(n5331) );
  XOR U6014 ( .A(n5332), .B(n5331), .Z(c[1183]) );
  NANDN U6015 ( .A(n5313), .B(n5312), .Z(n5317) );
  NAND U6016 ( .A(n5315), .B(n5314), .Z(n5316) );
  NAND U6017 ( .A(n5317), .B(n5316), .Z(n5343) );
  AND U6018 ( .A(b[2]), .B(a[162]), .Z(n5349) );
  AND U6019 ( .A(a[163]), .B(b[1]), .Z(n5347) );
  AND U6020 ( .A(a[161]), .B(b[3]), .Z(n5346) );
  XOR U6021 ( .A(n5347), .B(n5346), .Z(n5348) );
  XOR U6022 ( .A(n5349), .B(n5348), .Z(n5352) );
  NAND U6023 ( .A(b[0]), .B(a[164]), .Z(n5353) );
  XOR U6024 ( .A(n5352), .B(n5353), .Z(n5355) );
  OR U6025 ( .A(n5319), .B(n5318), .Z(n5323) );
  NANDN U6026 ( .A(n5321), .B(n5320), .Z(n5322) );
  NAND U6027 ( .A(n5323), .B(n5322), .Z(n5354) );
  XNOR U6028 ( .A(n5355), .B(n5354), .Z(n5340) );
  NANDN U6029 ( .A(n5325), .B(n5324), .Z(n5329) );
  OR U6030 ( .A(n5327), .B(n5326), .Z(n5328) );
  NAND U6031 ( .A(n5329), .B(n5328), .Z(n5341) );
  XNOR U6032 ( .A(n5340), .B(n5341), .Z(n5342) );
  XNOR U6033 ( .A(n5343), .B(n5342), .Z(n5335) );
  XOR U6034 ( .A(sreg[1184]), .B(n5335), .Z(n5336) );
  NAND U6035 ( .A(n5330), .B(sreg[1183]), .Z(n5334) );
  OR U6036 ( .A(n5332), .B(n5331), .Z(n5333) );
  NAND U6037 ( .A(n5334), .B(n5333), .Z(n5337) );
  XOR U6038 ( .A(n5336), .B(n5337), .Z(c[1184]) );
  OR U6039 ( .A(n5335), .B(sreg[1184]), .Z(n5339) );
  NANDN U6040 ( .A(n5337), .B(n5336), .Z(n5338) );
  AND U6041 ( .A(n5339), .B(n5338), .Z(n5377) );
  NANDN U6042 ( .A(n5341), .B(n5340), .Z(n5345) );
  NAND U6043 ( .A(n5343), .B(n5342), .Z(n5344) );
  NAND U6044 ( .A(n5345), .B(n5344), .Z(n5362) );
  AND U6045 ( .A(b[2]), .B(a[163]), .Z(n5368) );
  AND U6046 ( .A(a[164]), .B(b[1]), .Z(n5366) );
  AND U6047 ( .A(a[162]), .B(b[3]), .Z(n5365) );
  XOR U6048 ( .A(n5366), .B(n5365), .Z(n5367) );
  XOR U6049 ( .A(n5368), .B(n5367), .Z(n5371) );
  NAND U6050 ( .A(b[0]), .B(a[165]), .Z(n5372) );
  XOR U6051 ( .A(n5371), .B(n5372), .Z(n5374) );
  OR U6052 ( .A(n5347), .B(n5346), .Z(n5351) );
  NANDN U6053 ( .A(n5349), .B(n5348), .Z(n5350) );
  NAND U6054 ( .A(n5351), .B(n5350), .Z(n5373) );
  XNOR U6055 ( .A(n5374), .B(n5373), .Z(n5359) );
  NANDN U6056 ( .A(n5353), .B(n5352), .Z(n5357) );
  OR U6057 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U6058 ( .A(n5357), .B(n5356), .Z(n5360) );
  XNOR U6059 ( .A(n5359), .B(n5360), .Z(n5361) );
  XNOR U6060 ( .A(n5362), .B(n5361), .Z(n5378) );
  XOR U6061 ( .A(sreg[1185]), .B(n5378), .Z(n5358) );
  XOR U6062 ( .A(n5377), .B(n5358), .Z(c[1185]) );
  NANDN U6063 ( .A(n5360), .B(n5359), .Z(n5364) );
  NAND U6064 ( .A(n5362), .B(n5361), .Z(n5363) );
  NAND U6065 ( .A(n5364), .B(n5363), .Z(n5385) );
  AND U6066 ( .A(b[2]), .B(a[164]), .Z(n5391) );
  AND U6067 ( .A(a[165]), .B(b[1]), .Z(n5389) );
  AND U6068 ( .A(a[163]), .B(b[3]), .Z(n5388) );
  XOR U6069 ( .A(n5389), .B(n5388), .Z(n5390) );
  XOR U6070 ( .A(n5391), .B(n5390), .Z(n5394) );
  NAND U6071 ( .A(b[0]), .B(a[166]), .Z(n5395) );
  XOR U6072 ( .A(n5394), .B(n5395), .Z(n5397) );
  OR U6073 ( .A(n5366), .B(n5365), .Z(n5370) );
  NANDN U6074 ( .A(n5368), .B(n5367), .Z(n5369) );
  NAND U6075 ( .A(n5370), .B(n5369), .Z(n5396) );
  XNOR U6076 ( .A(n5397), .B(n5396), .Z(n5382) );
  NANDN U6077 ( .A(n5372), .B(n5371), .Z(n5376) );
  OR U6078 ( .A(n5374), .B(n5373), .Z(n5375) );
  NAND U6079 ( .A(n5376), .B(n5375), .Z(n5383) );
  XNOR U6080 ( .A(n5382), .B(n5383), .Z(n5384) );
  XNOR U6081 ( .A(n5385), .B(n5384), .Z(n5381) );
  XOR U6082 ( .A(n5380), .B(sreg[1186]), .Z(n5379) );
  XOR U6083 ( .A(n5381), .B(n5379), .Z(c[1186]) );
  NANDN U6084 ( .A(n5383), .B(n5382), .Z(n5387) );
  NAND U6085 ( .A(n5385), .B(n5384), .Z(n5386) );
  NAND U6086 ( .A(n5387), .B(n5386), .Z(n5403) );
  AND U6087 ( .A(b[2]), .B(a[165]), .Z(n5409) );
  AND U6088 ( .A(a[166]), .B(b[1]), .Z(n5407) );
  AND U6089 ( .A(a[164]), .B(b[3]), .Z(n5406) );
  XOR U6090 ( .A(n5407), .B(n5406), .Z(n5408) );
  XOR U6091 ( .A(n5409), .B(n5408), .Z(n5412) );
  NAND U6092 ( .A(b[0]), .B(a[167]), .Z(n5413) );
  XOR U6093 ( .A(n5412), .B(n5413), .Z(n5415) );
  OR U6094 ( .A(n5389), .B(n5388), .Z(n5393) );
  NANDN U6095 ( .A(n5391), .B(n5390), .Z(n5392) );
  NAND U6096 ( .A(n5393), .B(n5392), .Z(n5414) );
  XNOR U6097 ( .A(n5415), .B(n5414), .Z(n5400) );
  NANDN U6098 ( .A(n5395), .B(n5394), .Z(n5399) );
  OR U6099 ( .A(n5397), .B(n5396), .Z(n5398) );
  NAND U6100 ( .A(n5399), .B(n5398), .Z(n5401) );
  XNOR U6101 ( .A(n5400), .B(n5401), .Z(n5402) );
  XNOR U6102 ( .A(n5403), .B(n5402), .Z(n5418) );
  XNOR U6103 ( .A(n5418), .B(sreg[1187]), .Z(n5420) );
  XNOR U6104 ( .A(n5419), .B(n5420), .Z(c[1187]) );
  NANDN U6105 ( .A(n5401), .B(n5400), .Z(n5405) );
  NAND U6106 ( .A(n5403), .B(n5402), .Z(n5404) );
  NAND U6107 ( .A(n5405), .B(n5404), .Z(n5426) );
  AND U6108 ( .A(b[2]), .B(a[166]), .Z(n5432) );
  AND U6109 ( .A(a[167]), .B(b[1]), .Z(n5430) );
  AND U6110 ( .A(a[165]), .B(b[3]), .Z(n5429) );
  XOR U6111 ( .A(n5430), .B(n5429), .Z(n5431) );
  XOR U6112 ( .A(n5432), .B(n5431), .Z(n5435) );
  NAND U6113 ( .A(b[0]), .B(a[168]), .Z(n5436) );
  XOR U6114 ( .A(n5435), .B(n5436), .Z(n5438) );
  OR U6115 ( .A(n5407), .B(n5406), .Z(n5411) );
  NANDN U6116 ( .A(n5409), .B(n5408), .Z(n5410) );
  NAND U6117 ( .A(n5411), .B(n5410), .Z(n5437) );
  XNOR U6118 ( .A(n5438), .B(n5437), .Z(n5423) );
  NANDN U6119 ( .A(n5413), .B(n5412), .Z(n5417) );
  OR U6120 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U6121 ( .A(n5417), .B(n5416), .Z(n5424) );
  XNOR U6122 ( .A(n5423), .B(n5424), .Z(n5425) );
  XNOR U6123 ( .A(n5426), .B(n5425), .Z(n5441) );
  XNOR U6124 ( .A(n5441), .B(sreg[1188]), .Z(n5443) );
  NAND U6125 ( .A(n5418), .B(sreg[1187]), .Z(n5422) );
  NANDN U6126 ( .A(n5420), .B(n5419), .Z(n5421) );
  AND U6127 ( .A(n5422), .B(n5421), .Z(n5442) );
  XOR U6128 ( .A(n5443), .B(n5442), .Z(c[1188]) );
  NANDN U6129 ( .A(n5424), .B(n5423), .Z(n5428) );
  NAND U6130 ( .A(n5426), .B(n5425), .Z(n5427) );
  NAND U6131 ( .A(n5428), .B(n5427), .Z(n5452) );
  AND U6132 ( .A(b[2]), .B(a[167]), .Z(n5458) );
  AND U6133 ( .A(a[168]), .B(b[1]), .Z(n5456) );
  AND U6134 ( .A(a[166]), .B(b[3]), .Z(n5455) );
  XOR U6135 ( .A(n5456), .B(n5455), .Z(n5457) );
  XOR U6136 ( .A(n5458), .B(n5457), .Z(n5461) );
  NAND U6137 ( .A(b[0]), .B(a[169]), .Z(n5462) );
  XOR U6138 ( .A(n5461), .B(n5462), .Z(n5464) );
  OR U6139 ( .A(n5430), .B(n5429), .Z(n5434) );
  NANDN U6140 ( .A(n5432), .B(n5431), .Z(n5433) );
  NAND U6141 ( .A(n5434), .B(n5433), .Z(n5463) );
  XNOR U6142 ( .A(n5464), .B(n5463), .Z(n5449) );
  NANDN U6143 ( .A(n5436), .B(n5435), .Z(n5440) );
  OR U6144 ( .A(n5438), .B(n5437), .Z(n5439) );
  NAND U6145 ( .A(n5440), .B(n5439), .Z(n5450) );
  XNOR U6146 ( .A(n5449), .B(n5450), .Z(n5451) );
  XNOR U6147 ( .A(n5452), .B(n5451), .Z(n5448) );
  NAND U6148 ( .A(n5441), .B(sreg[1188]), .Z(n5445) );
  OR U6149 ( .A(n5443), .B(n5442), .Z(n5444) );
  AND U6150 ( .A(n5445), .B(n5444), .Z(n5447) );
  XNOR U6151 ( .A(n5447), .B(sreg[1189]), .Z(n5446) );
  XOR U6152 ( .A(n5448), .B(n5446), .Z(c[1189]) );
  NANDN U6153 ( .A(n5450), .B(n5449), .Z(n5454) );
  NAND U6154 ( .A(n5452), .B(n5451), .Z(n5453) );
  NAND U6155 ( .A(n5454), .B(n5453), .Z(n5470) );
  AND U6156 ( .A(b[2]), .B(a[168]), .Z(n5476) );
  AND U6157 ( .A(a[169]), .B(b[1]), .Z(n5474) );
  AND U6158 ( .A(a[167]), .B(b[3]), .Z(n5473) );
  XOR U6159 ( .A(n5474), .B(n5473), .Z(n5475) );
  XOR U6160 ( .A(n5476), .B(n5475), .Z(n5479) );
  NAND U6161 ( .A(b[0]), .B(a[170]), .Z(n5480) );
  XOR U6162 ( .A(n5479), .B(n5480), .Z(n5482) );
  OR U6163 ( .A(n5456), .B(n5455), .Z(n5460) );
  NANDN U6164 ( .A(n5458), .B(n5457), .Z(n5459) );
  NAND U6165 ( .A(n5460), .B(n5459), .Z(n5481) );
  XNOR U6166 ( .A(n5482), .B(n5481), .Z(n5467) );
  NANDN U6167 ( .A(n5462), .B(n5461), .Z(n5466) );
  OR U6168 ( .A(n5464), .B(n5463), .Z(n5465) );
  NAND U6169 ( .A(n5466), .B(n5465), .Z(n5468) );
  XNOR U6170 ( .A(n5467), .B(n5468), .Z(n5469) );
  XOR U6171 ( .A(n5470), .B(n5469), .Z(n5485) );
  XOR U6172 ( .A(sreg[1190]), .B(n5485), .Z(n5487) );
  XNOR U6173 ( .A(n5486), .B(n5487), .Z(c[1190]) );
  NANDN U6174 ( .A(n5468), .B(n5467), .Z(n5472) );
  NAND U6175 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U6176 ( .A(n5472), .B(n5471), .Z(n5493) );
  AND U6177 ( .A(b[2]), .B(a[169]), .Z(n5499) );
  AND U6178 ( .A(a[170]), .B(b[1]), .Z(n5497) );
  AND U6179 ( .A(a[168]), .B(b[3]), .Z(n5496) );
  XOR U6180 ( .A(n5497), .B(n5496), .Z(n5498) );
  XOR U6181 ( .A(n5499), .B(n5498), .Z(n5502) );
  NAND U6182 ( .A(b[0]), .B(a[171]), .Z(n5503) );
  XOR U6183 ( .A(n5502), .B(n5503), .Z(n5505) );
  OR U6184 ( .A(n5474), .B(n5473), .Z(n5478) );
  NANDN U6185 ( .A(n5476), .B(n5475), .Z(n5477) );
  NAND U6186 ( .A(n5478), .B(n5477), .Z(n5504) );
  XNOR U6187 ( .A(n5505), .B(n5504), .Z(n5490) );
  NANDN U6188 ( .A(n5480), .B(n5479), .Z(n5484) );
  OR U6189 ( .A(n5482), .B(n5481), .Z(n5483) );
  NAND U6190 ( .A(n5484), .B(n5483), .Z(n5491) );
  XNOR U6191 ( .A(n5490), .B(n5491), .Z(n5492) );
  XNOR U6192 ( .A(n5493), .B(n5492), .Z(n5508) );
  XOR U6193 ( .A(sreg[1191]), .B(n5508), .Z(n5509) );
  NANDN U6194 ( .A(n5485), .B(sreg[1190]), .Z(n5489) );
  NANDN U6195 ( .A(n5487), .B(n5486), .Z(n5488) );
  NAND U6196 ( .A(n5489), .B(n5488), .Z(n5510) );
  XOR U6197 ( .A(n5509), .B(n5510), .Z(c[1191]) );
  NANDN U6198 ( .A(n5491), .B(n5490), .Z(n5495) );
  NAND U6199 ( .A(n5493), .B(n5492), .Z(n5494) );
  NAND U6200 ( .A(n5495), .B(n5494), .Z(n5516) );
  AND U6201 ( .A(b[2]), .B(a[170]), .Z(n5522) );
  AND U6202 ( .A(a[171]), .B(b[1]), .Z(n5520) );
  AND U6203 ( .A(a[169]), .B(b[3]), .Z(n5519) );
  XOR U6204 ( .A(n5520), .B(n5519), .Z(n5521) );
  XOR U6205 ( .A(n5522), .B(n5521), .Z(n5525) );
  NAND U6206 ( .A(b[0]), .B(a[172]), .Z(n5526) );
  XOR U6207 ( .A(n5525), .B(n5526), .Z(n5528) );
  OR U6208 ( .A(n5497), .B(n5496), .Z(n5501) );
  NANDN U6209 ( .A(n5499), .B(n5498), .Z(n5500) );
  NAND U6210 ( .A(n5501), .B(n5500), .Z(n5527) );
  XNOR U6211 ( .A(n5528), .B(n5527), .Z(n5513) );
  NANDN U6212 ( .A(n5503), .B(n5502), .Z(n5507) );
  OR U6213 ( .A(n5505), .B(n5504), .Z(n5506) );
  NAND U6214 ( .A(n5507), .B(n5506), .Z(n5514) );
  XNOR U6215 ( .A(n5513), .B(n5514), .Z(n5515) );
  XNOR U6216 ( .A(n5516), .B(n5515), .Z(n5531) );
  XOR U6217 ( .A(sreg[1192]), .B(n5531), .Z(n5532) );
  OR U6218 ( .A(n5508), .B(sreg[1191]), .Z(n5512) );
  NANDN U6219 ( .A(n5510), .B(n5509), .Z(n5511) );
  AND U6220 ( .A(n5512), .B(n5511), .Z(n5533) );
  XOR U6221 ( .A(n5532), .B(n5533), .Z(c[1192]) );
  NANDN U6222 ( .A(n5514), .B(n5513), .Z(n5518) );
  NAND U6223 ( .A(n5516), .B(n5515), .Z(n5517) );
  NAND U6224 ( .A(n5518), .B(n5517), .Z(n5542) );
  AND U6225 ( .A(b[2]), .B(a[171]), .Z(n5554) );
  AND U6226 ( .A(a[172]), .B(b[1]), .Z(n5552) );
  AND U6227 ( .A(a[170]), .B(b[3]), .Z(n5551) );
  XOR U6228 ( .A(n5552), .B(n5551), .Z(n5553) );
  XOR U6229 ( .A(n5554), .B(n5553), .Z(n5545) );
  NAND U6230 ( .A(b[0]), .B(a[173]), .Z(n5546) );
  XOR U6231 ( .A(n5545), .B(n5546), .Z(n5548) );
  OR U6232 ( .A(n5520), .B(n5519), .Z(n5524) );
  NANDN U6233 ( .A(n5522), .B(n5521), .Z(n5523) );
  NAND U6234 ( .A(n5524), .B(n5523), .Z(n5547) );
  XNOR U6235 ( .A(n5548), .B(n5547), .Z(n5539) );
  NANDN U6236 ( .A(n5526), .B(n5525), .Z(n5530) );
  OR U6237 ( .A(n5528), .B(n5527), .Z(n5529) );
  NAND U6238 ( .A(n5530), .B(n5529), .Z(n5540) );
  XNOR U6239 ( .A(n5539), .B(n5540), .Z(n5541) );
  XOR U6240 ( .A(n5542), .B(n5541), .Z(n5538) );
  OR U6241 ( .A(n5531), .B(sreg[1192]), .Z(n5535) );
  NANDN U6242 ( .A(n5533), .B(n5532), .Z(n5534) );
  AND U6243 ( .A(n5535), .B(n5534), .Z(n5537) );
  XNOR U6244 ( .A(sreg[1193]), .B(n5537), .Z(n5536) );
  XOR U6245 ( .A(n5538), .B(n5536), .Z(c[1193]) );
  NANDN U6246 ( .A(n5540), .B(n5539), .Z(n5544) );
  NAND U6247 ( .A(n5542), .B(n5541), .Z(n5543) );
  NAND U6248 ( .A(n5544), .B(n5543), .Z(n5577) );
  NANDN U6249 ( .A(n5546), .B(n5545), .Z(n5550) );
  OR U6250 ( .A(n5548), .B(n5547), .Z(n5549) );
  NAND U6251 ( .A(n5550), .B(n5549), .Z(n5574) );
  AND U6252 ( .A(b[2]), .B(a[172]), .Z(n5565) );
  AND U6253 ( .A(a[173]), .B(b[1]), .Z(n5563) );
  AND U6254 ( .A(a[171]), .B(b[3]), .Z(n5562) );
  XOR U6255 ( .A(n5563), .B(n5562), .Z(n5564) );
  XOR U6256 ( .A(n5565), .B(n5564), .Z(n5568) );
  NAND U6257 ( .A(b[0]), .B(a[174]), .Z(n5569) );
  XNOR U6258 ( .A(n5568), .B(n5569), .Z(n5570) );
  OR U6259 ( .A(n5552), .B(n5551), .Z(n5556) );
  NANDN U6260 ( .A(n5554), .B(n5553), .Z(n5555) );
  AND U6261 ( .A(n5556), .B(n5555), .Z(n5571) );
  XNOR U6262 ( .A(n5570), .B(n5571), .Z(n5575) );
  XNOR U6263 ( .A(n5574), .B(n5575), .Z(n5576) );
  XOR U6264 ( .A(n5577), .B(n5576), .Z(n5557) );
  XNOR U6265 ( .A(sreg[1194]), .B(n5557), .Z(n5558) );
  XNOR U6266 ( .A(n5559), .B(n5558), .Z(c[1194]) );
  NANDN U6267 ( .A(sreg[1194]), .B(n5557), .Z(n5561) );
  NAND U6268 ( .A(n5559), .B(n5558), .Z(n5560) );
  AND U6269 ( .A(n5561), .B(n5560), .Z(n5599) );
  AND U6270 ( .A(b[2]), .B(a[173]), .Z(n5590) );
  AND U6271 ( .A(a[174]), .B(b[1]), .Z(n5588) );
  AND U6272 ( .A(a[172]), .B(b[3]), .Z(n5587) );
  XOR U6273 ( .A(n5588), .B(n5587), .Z(n5589) );
  XOR U6274 ( .A(n5590), .B(n5589), .Z(n5593) );
  NAND U6275 ( .A(b[0]), .B(a[175]), .Z(n5594) );
  XOR U6276 ( .A(n5593), .B(n5594), .Z(n5596) );
  OR U6277 ( .A(n5563), .B(n5562), .Z(n5567) );
  NANDN U6278 ( .A(n5565), .B(n5564), .Z(n5566) );
  NAND U6279 ( .A(n5567), .B(n5566), .Z(n5595) );
  XNOR U6280 ( .A(n5596), .B(n5595), .Z(n5581) );
  NANDN U6281 ( .A(n5569), .B(n5568), .Z(n5573) );
  NAND U6282 ( .A(n5571), .B(n5570), .Z(n5572) );
  NAND U6283 ( .A(n5573), .B(n5572), .Z(n5582) );
  XNOR U6284 ( .A(n5581), .B(n5582), .Z(n5583) );
  NANDN U6285 ( .A(n5575), .B(n5574), .Z(n5579) );
  NANDN U6286 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U6287 ( .A(n5579), .B(n5578), .Z(n5584) );
  XNOR U6288 ( .A(n5583), .B(n5584), .Z(n5600) );
  XOR U6289 ( .A(sreg[1195]), .B(n5600), .Z(n5580) );
  XOR U6290 ( .A(n5599), .B(n5580), .Z(c[1195]) );
  NANDN U6291 ( .A(n5582), .B(n5581), .Z(n5586) );
  NAND U6292 ( .A(n5584), .B(n5583), .Z(n5585) );
  NAND U6293 ( .A(n5586), .B(n5585), .Z(n5617) );
  AND U6294 ( .A(b[2]), .B(a[174]), .Z(n5611) );
  AND U6295 ( .A(a[175]), .B(b[1]), .Z(n5609) );
  AND U6296 ( .A(a[173]), .B(b[3]), .Z(n5608) );
  XOR U6297 ( .A(n5609), .B(n5608), .Z(n5610) );
  XOR U6298 ( .A(n5611), .B(n5610), .Z(n5602) );
  NAND U6299 ( .A(b[0]), .B(a[176]), .Z(n5603) );
  XOR U6300 ( .A(n5602), .B(n5603), .Z(n5605) );
  OR U6301 ( .A(n5588), .B(n5587), .Z(n5592) );
  NANDN U6302 ( .A(n5590), .B(n5589), .Z(n5591) );
  NAND U6303 ( .A(n5592), .B(n5591), .Z(n5604) );
  XNOR U6304 ( .A(n5605), .B(n5604), .Z(n5614) );
  NANDN U6305 ( .A(n5594), .B(n5593), .Z(n5598) );
  OR U6306 ( .A(n5596), .B(n5595), .Z(n5597) );
  NAND U6307 ( .A(n5598), .B(n5597), .Z(n5615) );
  XNOR U6308 ( .A(n5614), .B(n5615), .Z(n5616) );
  XOR U6309 ( .A(n5617), .B(n5616), .Z(n5621) );
  XOR U6310 ( .A(sreg[1196]), .B(n5620), .Z(n5601) );
  XOR U6311 ( .A(n5621), .B(n5601), .Z(c[1196]) );
  NANDN U6312 ( .A(n5603), .B(n5602), .Z(n5607) );
  OR U6313 ( .A(n5605), .B(n5604), .Z(n5606) );
  NAND U6314 ( .A(n5607), .B(n5606), .Z(n5623) );
  AND U6315 ( .A(b[2]), .B(a[175]), .Z(n5638) );
  AND U6316 ( .A(a[176]), .B(b[1]), .Z(n5636) );
  AND U6317 ( .A(a[174]), .B(b[3]), .Z(n5635) );
  XOR U6318 ( .A(n5636), .B(n5635), .Z(n5637) );
  XOR U6319 ( .A(n5638), .B(n5637), .Z(n5629) );
  NAND U6320 ( .A(b[0]), .B(a[177]), .Z(n5630) );
  XNOR U6321 ( .A(n5629), .B(n5630), .Z(n5631) );
  OR U6322 ( .A(n5609), .B(n5608), .Z(n5613) );
  NANDN U6323 ( .A(n5611), .B(n5610), .Z(n5612) );
  AND U6324 ( .A(n5613), .B(n5612), .Z(n5632) );
  XNOR U6325 ( .A(n5631), .B(n5632), .Z(n5624) );
  XNOR U6326 ( .A(n5623), .B(n5624), .Z(n5625) );
  NANDN U6327 ( .A(n5615), .B(n5614), .Z(n5619) );
  NAND U6328 ( .A(n5617), .B(n5616), .Z(n5618) );
  NAND U6329 ( .A(n5619), .B(n5618), .Z(n5626) );
  XOR U6330 ( .A(n5625), .B(n5626), .Z(n5643) );
  XOR U6331 ( .A(n5642), .B(sreg[1197]), .Z(n5622) );
  XNOR U6332 ( .A(n5643), .B(n5622), .Z(c[1197]) );
  NANDN U6333 ( .A(n5624), .B(n5623), .Z(n5628) );
  NANDN U6334 ( .A(n5626), .B(n5625), .Z(n5627) );
  NAND U6335 ( .A(n5628), .B(n5627), .Z(n5649) );
  NANDN U6336 ( .A(n5630), .B(n5629), .Z(n5634) );
  NAND U6337 ( .A(n5632), .B(n5631), .Z(n5633) );
  AND U6338 ( .A(n5634), .B(n5633), .Z(n5648) );
  AND U6339 ( .A(b[2]), .B(a[176]), .Z(n5653) );
  AND U6340 ( .A(a[177]), .B(b[1]), .Z(n5651) );
  AND U6341 ( .A(a[175]), .B(b[3]), .Z(n5650) );
  XOR U6342 ( .A(n5651), .B(n5650), .Z(n5652) );
  XOR U6343 ( .A(n5653), .B(n5652), .Z(n5656) );
  NAND U6344 ( .A(b[0]), .B(a[178]), .Z(n5657) );
  XOR U6345 ( .A(n5656), .B(n5657), .Z(n5659) );
  OR U6346 ( .A(n5636), .B(n5635), .Z(n5640) );
  NANDN U6347 ( .A(n5638), .B(n5637), .Z(n5639) );
  NAND U6348 ( .A(n5640), .B(n5639), .Z(n5658) );
  XOR U6349 ( .A(n5659), .B(n5658), .Z(n5647) );
  XNOR U6350 ( .A(n5648), .B(n5647), .Z(n5641) );
  XOR U6351 ( .A(n5649), .B(n5641), .Z(n5646) );
  XOR U6352 ( .A(sreg[1198]), .B(n5645), .Z(n5644) );
  XNOR U6353 ( .A(n5646), .B(n5644), .Z(c[1198]) );
  AND U6354 ( .A(b[2]), .B(a[177]), .Z(n5676) );
  AND U6355 ( .A(a[178]), .B(b[1]), .Z(n5674) );
  AND U6356 ( .A(a[176]), .B(b[3]), .Z(n5673) );
  XOR U6357 ( .A(n5674), .B(n5673), .Z(n5675) );
  XOR U6358 ( .A(n5676), .B(n5675), .Z(n5667) );
  NAND U6359 ( .A(b[0]), .B(a[179]), .Z(n5668) );
  XOR U6360 ( .A(n5667), .B(n5668), .Z(n5670) );
  OR U6361 ( .A(n5651), .B(n5650), .Z(n5655) );
  NANDN U6362 ( .A(n5653), .B(n5652), .Z(n5654) );
  NAND U6363 ( .A(n5655), .B(n5654), .Z(n5669) );
  XNOR U6364 ( .A(n5670), .B(n5669), .Z(n5679) );
  NANDN U6365 ( .A(n5657), .B(n5656), .Z(n5661) );
  OR U6366 ( .A(n5659), .B(n5658), .Z(n5660) );
  NAND U6367 ( .A(n5661), .B(n5660), .Z(n5680) );
  XNOR U6368 ( .A(n5679), .B(n5680), .Z(n5681) );
  XOR U6369 ( .A(n5682), .B(n5681), .Z(n5662) );
  XNOR U6370 ( .A(n5662), .B(sreg[1199]), .Z(n5663) );
  XOR U6371 ( .A(n5664), .B(n5663), .Z(c[1199]) );
  NAND U6372 ( .A(n5662), .B(sreg[1199]), .Z(n5666) );
  OR U6373 ( .A(n5664), .B(n5663), .Z(n5665) );
  NAND U6374 ( .A(n5666), .B(n5665), .Z(n5686) );
  NANDN U6375 ( .A(n5668), .B(n5667), .Z(n5672) );
  OR U6376 ( .A(n5670), .B(n5669), .Z(n5671) );
  NAND U6377 ( .A(n5672), .B(n5671), .Z(n5688) );
  AND U6378 ( .A(b[2]), .B(a[178]), .Z(n5697) );
  AND U6379 ( .A(a[179]), .B(b[1]), .Z(n5695) );
  AND U6380 ( .A(a[177]), .B(b[3]), .Z(n5694) );
  XOR U6381 ( .A(n5695), .B(n5694), .Z(n5696) );
  XOR U6382 ( .A(n5697), .B(n5696), .Z(n5700) );
  NAND U6383 ( .A(b[0]), .B(a[180]), .Z(n5701) );
  XNOR U6384 ( .A(n5700), .B(n5701), .Z(n5702) );
  OR U6385 ( .A(n5674), .B(n5673), .Z(n5678) );
  NANDN U6386 ( .A(n5676), .B(n5675), .Z(n5677) );
  AND U6387 ( .A(n5678), .B(n5677), .Z(n5703) );
  XNOR U6388 ( .A(n5702), .B(n5703), .Z(n5689) );
  XNOR U6389 ( .A(n5688), .B(n5689), .Z(n5690) );
  NANDN U6390 ( .A(n5680), .B(n5679), .Z(n5684) );
  NANDN U6391 ( .A(n5682), .B(n5681), .Z(n5683) );
  AND U6392 ( .A(n5684), .B(n5683), .Z(n5691) );
  XNOR U6393 ( .A(n5690), .B(n5691), .Z(n5687) );
  XOR U6394 ( .A(sreg[1200]), .B(n5687), .Z(n5685) );
  XNOR U6395 ( .A(n5686), .B(n5685), .Z(c[1200]) );
  NANDN U6396 ( .A(n5689), .B(n5688), .Z(n5693) );
  NAND U6397 ( .A(n5691), .B(n5690), .Z(n5692) );
  NAND U6398 ( .A(n5693), .B(n5692), .Z(n5709) );
  AND U6399 ( .A(b[2]), .B(a[179]), .Z(n5713) );
  AND U6400 ( .A(a[180]), .B(b[1]), .Z(n5711) );
  AND U6401 ( .A(a[178]), .B(b[3]), .Z(n5710) );
  XOR U6402 ( .A(n5711), .B(n5710), .Z(n5712) );
  XOR U6403 ( .A(n5713), .B(n5712), .Z(n5716) );
  NAND U6404 ( .A(b[0]), .B(a[181]), .Z(n5717) );
  XOR U6405 ( .A(n5716), .B(n5717), .Z(n5718) );
  OR U6406 ( .A(n5695), .B(n5694), .Z(n5699) );
  NANDN U6407 ( .A(n5697), .B(n5696), .Z(n5698) );
  AND U6408 ( .A(n5699), .B(n5698), .Z(n5719) );
  XOR U6409 ( .A(n5718), .B(n5719), .Z(n5707) );
  NANDN U6410 ( .A(n5701), .B(n5700), .Z(n5705) );
  NAND U6411 ( .A(n5703), .B(n5702), .Z(n5704) );
  AND U6412 ( .A(n5705), .B(n5704), .Z(n5708) );
  XOR U6413 ( .A(n5707), .B(n5708), .Z(n5706) );
  XOR U6414 ( .A(n5709), .B(n5706), .Z(n5720) );
  XNOR U6415 ( .A(n5720), .B(sreg[1201]), .Z(n5721) );
  XOR U6416 ( .A(n5722), .B(n5721), .Z(c[1201]) );
  AND U6417 ( .A(b[2]), .B(a[180]), .Z(n5737) );
  AND U6418 ( .A(a[181]), .B(b[1]), .Z(n5735) );
  AND U6419 ( .A(a[179]), .B(b[3]), .Z(n5734) );
  XOR U6420 ( .A(n5735), .B(n5734), .Z(n5736) );
  XOR U6421 ( .A(n5737), .B(n5736), .Z(n5740) );
  NAND U6422 ( .A(b[0]), .B(a[182]), .Z(n5741) );
  XOR U6423 ( .A(n5740), .B(n5741), .Z(n5743) );
  OR U6424 ( .A(n5711), .B(n5710), .Z(n5715) );
  NANDN U6425 ( .A(n5713), .B(n5712), .Z(n5714) );
  NAND U6426 ( .A(n5715), .B(n5714), .Z(n5742) );
  XNOR U6427 ( .A(n5743), .B(n5742), .Z(n5728) );
  XNOR U6428 ( .A(n5728), .B(n5729), .Z(n5731) );
  XOR U6429 ( .A(n5730), .B(n5731), .Z(n5727) );
  NAND U6430 ( .A(n5720), .B(sreg[1201]), .Z(n5724) );
  OR U6431 ( .A(n5722), .B(n5721), .Z(n5723) );
  AND U6432 ( .A(n5724), .B(n5723), .Z(n5726) );
  XNOR U6433 ( .A(n5726), .B(sreg[1202]), .Z(n5725) );
  XNOR U6434 ( .A(n5727), .B(n5725), .Z(c[1202]) );
  NANDN U6435 ( .A(n5729), .B(n5728), .Z(n5733) );
  NAND U6436 ( .A(n5731), .B(n5730), .Z(n5732) );
  NAND U6437 ( .A(n5733), .B(n5732), .Z(n5754) );
  AND U6438 ( .A(b[2]), .B(a[181]), .Z(n5760) );
  AND U6439 ( .A(a[182]), .B(b[1]), .Z(n5758) );
  AND U6440 ( .A(a[180]), .B(b[3]), .Z(n5757) );
  XOR U6441 ( .A(n5758), .B(n5757), .Z(n5759) );
  XOR U6442 ( .A(n5760), .B(n5759), .Z(n5763) );
  NAND U6443 ( .A(b[0]), .B(a[183]), .Z(n5764) );
  XOR U6444 ( .A(n5763), .B(n5764), .Z(n5766) );
  OR U6445 ( .A(n5735), .B(n5734), .Z(n5739) );
  NANDN U6446 ( .A(n5737), .B(n5736), .Z(n5738) );
  NAND U6447 ( .A(n5739), .B(n5738), .Z(n5765) );
  XNOR U6448 ( .A(n5766), .B(n5765), .Z(n5751) );
  NANDN U6449 ( .A(n5741), .B(n5740), .Z(n5745) );
  OR U6450 ( .A(n5743), .B(n5742), .Z(n5744) );
  NAND U6451 ( .A(n5745), .B(n5744), .Z(n5752) );
  XNOR U6452 ( .A(n5751), .B(n5752), .Z(n5753) );
  XNOR U6453 ( .A(n5754), .B(n5753), .Z(n5746) );
  XOR U6454 ( .A(sreg[1203]), .B(n5746), .Z(n5747) );
  XOR U6455 ( .A(n5748), .B(n5747), .Z(c[1203]) );
  OR U6456 ( .A(n5746), .B(sreg[1203]), .Z(n5750) );
  NANDN U6457 ( .A(n5748), .B(n5747), .Z(n5749) );
  AND U6458 ( .A(n5750), .B(n5749), .Z(n5770) );
  NANDN U6459 ( .A(n5752), .B(n5751), .Z(n5756) );
  NAND U6460 ( .A(n5754), .B(n5753), .Z(n5755) );
  NAND U6461 ( .A(n5756), .B(n5755), .Z(n5775) );
  AND U6462 ( .A(b[2]), .B(a[182]), .Z(n5781) );
  AND U6463 ( .A(a[183]), .B(b[1]), .Z(n5779) );
  AND U6464 ( .A(a[181]), .B(b[3]), .Z(n5778) );
  XOR U6465 ( .A(n5779), .B(n5778), .Z(n5780) );
  XOR U6466 ( .A(n5781), .B(n5780), .Z(n5784) );
  NAND U6467 ( .A(b[0]), .B(a[184]), .Z(n5785) );
  XOR U6468 ( .A(n5784), .B(n5785), .Z(n5787) );
  OR U6469 ( .A(n5758), .B(n5757), .Z(n5762) );
  NANDN U6470 ( .A(n5760), .B(n5759), .Z(n5761) );
  NAND U6471 ( .A(n5762), .B(n5761), .Z(n5786) );
  XNOR U6472 ( .A(n5787), .B(n5786), .Z(n5772) );
  NANDN U6473 ( .A(n5764), .B(n5763), .Z(n5768) );
  OR U6474 ( .A(n5766), .B(n5765), .Z(n5767) );
  NAND U6475 ( .A(n5768), .B(n5767), .Z(n5773) );
  XNOR U6476 ( .A(n5772), .B(n5773), .Z(n5774) );
  XNOR U6477 ( .A(n5775), .B(n5774), .Z(n5771) );
  XOR U6478 ( .A(sreg[1204]), .B(n5771), .Z(n5769) );
  XOR U6479 ( .A(n5770), .B(n5769), .Z(c[1204]) );
  NANDN U6480 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U6481 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U6482 ( .A(n5777), .B(n5776), .Z(n5793) );
  AND U6483 ( .A(b[2]), .B(a[183]), .Z(n5799) );
  AND U6484 ( .A(a[184]), .B(b[1]), .Z(n5797) );
  AND U6485 ( .A(a[182]), .B(b[3]), .Z(n5796) );
  XOR U6486 ( .A(n5797), .B(n5796), .Z(n5798) );
  XOR U6487 ( .A(n5799), .B(n5798), .Z(n5802) );
  NAND U6488 ( .A(b[0]), .B(a[185]), .Z(n5803) );
  XOR U6489 ( .A(n5802), .B(n5803), .Z(n5805) );
  OR U6490 ( .A(n5779), .B(n5778), .Z(n5783) );
  NANDN U6491 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U6492 ( .A(n5783), .B(n5782), .Z(n5804) );
  XNOR U6493 ( .A(n5805), .B(n5804), .Z(n5790) );
  NANDN U6494 ( .A(n5785), .B(n5784), .Z(n5789) );
  OR U6495 ( .A(n5787), .B(n5786), .Z(n5788) );
  NAND U6496 ( .A(n5789), .B(n5788), .Z(n5791) );
  XNOR U6497 ( .A(n5790), .B(n5791), .Z(n5792) );
  XNOR U6498 ( .A(n5793), .B(n5792), .Z(n5808) );
  XNOR U6499 ( .A(n5808), .B(sreg[1205]), .Z(n5810) );
  XNOR U6500 ( .A(n5809), .B(n5810), .Z(c[1205]) );
  NANDN U6501 ( .A(n5791), .B(n5790), .Z(n5795) );
  NAND U6502 ( .A(n5793), .B(n5792), .Z(n5794) );
  NAND U6503 ( .A(n5795), .B(n5794), .Z(n5816) );
  AND U6504 ( .A(b[2]), .B(a[184]), .Z(n5822) );
  AND U6505 ( .A(a[185]), .B(b[1]), .Z(n5820) );
  AND U6506 ( .A(a[183]), .B(b[3]), .Z(n5819) );
  XOR U6507 ( .A(n5820), .B(n5819), .Z(n5821) );
  XOR U6508 ( .A(n5822), .B(n5821), .Z(n5825) );
  NAND U6509 ( .A(b[0]), .B(a[186]), .Z(n5826) );
  XOR U6510 ( .A(n5825), .B(n5826), .Z(n5828) );
  OR U6511 ( .A(n5797), .B(n5796), .Z(n5801) );
  NANDN U6512 ( .A(n5799), .B(n5798), .Z(n5800) );
  NAND U6513 ( .A(n5801), .B(n5800), .Z(n5827) );
  XNOR U6514 ( .A(n5828), .B(n5827), .Z(n5813) );
  NANDN U6515 ( .A(n5803), .B(n5802), .Z(n5807) );
  OR U6516 ( .A(n5805), .B(n5804), .Z(n5806) );
  NAND U6517 ( .A(n5807), .B(n5806), .Z(n5814) );
  XNOR U6518 ( .A(n5813), .B(n5814), .Z(n5815) );
  XNOR U6519 ( .A(n5816), .B(n5815), .Z(n5831) );
  XNOR U6520 ( .A(n5831), .B(sreg[1206]), .Z(n5833) );
  NAND U6521 ( .A(n5808), .B(sreg[1205]), .Z(n5812) );
  NANDN U6522 ( .A(n5810), .B(n5809), .Z(n5811) );
  AND U6523 ( .A(n5812), .B(n5811), .Z(n5832) );
  XOR U6524 ( .A(n5833), .B(n5832), .Z(c[1206]) );
  NANDN U6525 ( .A(n5814), .B(n5813), .Z(n5818) );
  NAND U6526 ( .A(n5816), .B(n5815), .Z(n5817) );
  NAND U6527 ( .A(n5818), .B(n5817), .Z(n5839) );
  AND U6528 ( .A(b[2]), .B(a[185]), .Z(n5845) );
  AND U6529 ( .A(a[186]), .B(b[1]), .Z(n5843) );
  AND U6530 ( .A(a[184]), .B(b[3]), .Z(n5842) );
  XOR U6531 ( .A(n5843), .B(n5842), .Z(n5844) );
  XOR U6532 ( .A(n5845), .B(n5844), .Z(n5848) );
  NAND U6533 ( .A(b[0]), .B(a[187]), .Z(n5849) );
  XOR U6534 ( .A(n5848), .B(n5849), .Z(n5851) );
  OR U6535 ( .A(n5820), .B(n5819), .Z(n5824) );
  NANDN U6536 ( .A(n5822), .B(n5821), .Z(n5823) );
  NAND U6537 ( .A(n5824), .B(n5823), .Z(n5850) );
  XNOR U6538 ( .A(n5851), .B(n5850), .Z(n5836) );
  NANDN U6539 ( .A(n5826), .B(n5825), .Z(n5830) );
  OR U6540 ( .A(n5828), .B(n5827), .Z(n5829) );
  NAND U6541 ( .A(n5830), .B(n5829), .Z(n5837) );
  XNOR U6542 ( .A(n5836), .B(n5837), .Z(n5838) );
  XNOR U6543 ( .A(n5839), .B(n5838), .Z(n5854) );
  XOR U6544 ( .A(sreg[1207]), .B(n5854), .Z(n5855) );
  NAND U6545 ( .A(n5831), .B(sreg[1206]), .Z(n5835) );
  OR U6546 ( .A(n5833), .B(n5832), .Z(n5834) );
  NAND U6547 ( .A(n5835), .B(n5834), .Z(n5856) );
  XOR U6548 ( .A(n5855), .B(n5856), .Z(c[1207]) );
  NANDN U6549 ( .A(n5837), .B(n5836), .Z(n5841) );
  NAND U6550 ( .A(n5839), .B(n5838), .Z(n5840) );
  NAND U6551 ( .A(n5841), .B(n5840), .Z(n5865) );
  AND U6552 ( .A(b[2]), .B(a[186]), .Z(n5871) );
  AND U6553 ( .A(a[187]), .B(b[1]), .Z(n5869) );
  AND U6554 ( .A(a[185]), .B(b[3]), .Z(n5868) );
  XOR U6555 ( .A(n5869), .B(n5868), .Z(n5870) );
  XOR U6556 ( .A(n5871), .B(n5870), .Z(n5874) );
  NAND U6557 ( .A(b[0]), .B(a[188]), .Z(n5875) );
  XOR U6558 ( .A(n5874), .B(n5875), .Z(n5877) );
  OR U6559 ( .A(n5843), .B(n5842), .Z(n5847) );
  NANDN U6560 ( .A(n5845), .B(n5844), .Z(n5846) );
  NAND U6561 ( .A(n5847), .B(n5846), .Z(n5876) );
  XNOR U6562 ( .A(n5877), .B(n5876), .Z(n5862) );
  NANDN U6563 ( .A(n5849), .B(n5848), .Z(n5853) );
  OR U6564 ( .A(n5851), .B(n5850), .Z(n5852) );
  NAND U6565 ( .A(n5853), .B(n5852), .Z(n5863) );
  XNOR U6566 ( .A(n5862), .B(n5863), .Z(n5864) );
  XOR U6567 ( .A(n5865), .B(n5864), .Z(n5861) );
  OR U6568 ( .A(n5854), .B(sreg[1207]), .Z(n5858) );
  NANDN U6569 ( .A(n5856), .B(n5855), .Z(n5857) );
  AND U6570 ( .A(n5858), .B(n5857), .Z(n5860) );
  XNOR U6571 ( .A(sreg[1208]), .B(n5860), .Z(n5859) );
  XOR U6572 ( .A(n5861), .B(n5859), .Z(c[1208]) );
  NANDN U6573 ( .A(n5863), .B(n5862), .Z(n5867) );
  NAND U6574 ( .A(n5865), .B(n5864), .Z(n5866) );
  NAND U6575 ( .A(n5867), .B(n5866), .Z(n5883) );
  AND U6576 ( .A(b[2]), .B(a[187]), .Z(n5889) );
  AND U6577 ( .A(a[188]), .B(b[1]), .Z(n5887) );
  AND U6578 ( .A(a[186]), .B(b[3]), .Z(n5886) );
  XOR U6579 ( .A(n5887), .B(n5886), .Z(n5888) );
  XOR U6580 ( .A(n5889), .B(n5888), .Z(n5892) );
  NAND U6581 ( .A(b[0]), .B(a[189]), .Z(n5893) );
  XOR U6582 ( .A(n5892), .B(n5893), .Z(n5895) );
  OR U6583 ( .A(n5869), .B(n5868), .Z(n5873) );
  NANDN U6584 ( .A(n5871), .B(n5870), .Z(n5872) );
  NAND U6585 ( .A(n5873), .B(n5872), .Z(n5894) );
  XNOR U6586 ( .A(n5895), .B(n5894), .Z(n5880) );
  NANDN U6587 ( .A(n5875), .B(n5874), .Z(n5879) );
  OR U6588 ( .A(n5877), .B(n5876), .Z(n5878) );
  NAND U6589 ( .A(n5879), .B(n5878), .Z(n5881) );
  XNOR U6590 ( .A(n5880), .B(n5881), .Z(n5882) );
  XNOR U6591 ( .A(n5883), .B(n5882), .Z(n5898) );
  XNOR U6592 ( .A(n5898), .B(sreg[1209]), .Z(n5899) );
  XOR U6593 ( .A(n5900), .B(n5899), .Z(c[1209]) );
  NANDN U6594 ( .A(n5881), .B(n5880), .Z(n5885) );
  NAND U6595 ( .A(n5883), .B(n5882), .Z(n5884) );
  NAND U6596 ( .A(n5885), .B(n5884), .Z(n5906) );
  AND U6597 ( .A(b[2]), .B(a[188]), .Z(n5912) );
  AND U6598 ( .A(a[189]), .B(b[1]), .Z(n5910) );
  AND U6599 ( .A(a[187]), .B(b[3]), .Z(n5909) );
  XOR U6600 ( .A(n5910), .B(n5909), .Z(n5911) );
  XOR U6601 ( .A(n5912), .B(n5911), .Z(n5915) );
  NAND U6602 ( .A(b[0]), .B(a[190]), .Z(n5916) );
  XOR U6603 ( .A(n5915), .B(n5916), .Z(n5918) );
  OR U6604 ( .A(n5887), .B(n5886), .Z(n5891) );
  NANDN U6605 ( .A(n5889), .B(n5888), .Z(n5890) );
  NAND U6606 ( .A(n5891), .B(n5890), .Z(n5917) );
  XNOR U6607 ( .A(n5918), .B(n5917), .Z(n5903) );
  NANDN U6608 ( .A(n5893), .B(n5892), .Z(n5897) );
  OR U6609 ( .A(n5895), .B(n5894), .Z(n5896) );
  NAND U6610 ( .A(n5897), .B(n5896), .Z(n5904) );
  XNOR U6611 ( .A(n5903), .B(n5904), .Z(n5905) );
  XNOR U6612 ( .A(n5906), .B(n5905), .Z(n5921) );
  XOR U6613 ( .A(sreg[1210]), .B(n5921), .Z(n5922) );
  NAND U6614 ( .A(n5898), .B(sreg[1209]), .Z(n5902) );
  OR U6615 ( .A(n5900), .B(n5899), .Z(n5901) );
  NAND U6616 ( .A(n5902), .B(n5901), .Z(n5923) );
  XOR U6617 ( .A(n5922), .B(n5923), .Z(c[1210]) );
  NANDN U6618 ( .A(n5904), .B(n5903), .Z(n5908) );
  NAND U6619 ( .A(n5906), .B(n5905), .Z(n5907) );
  NAND U6620 ( .A(n5908), .B(n5907), .Z(n5932) );
  AND U6621 ( .A(b[2]), .B(a[189]), .Z(n5938) );
  AND U6622 ( .A(a[190]), .B(b[1]), .Z(n5936) );
  AND U6623 ( .A(a[188]), .B(b[3]), .Z(n5935) );
  XOR U6624 ( .A(n5936), .B(n5935), .Z(n5937) );
  XOR U6625 ( .A(n5938), .B(n5937), .Z(n5941) );
  NAND U6626 ( .A(b[0]), .B(a[191]), .Z(n5942) );
  XOR U6627 ( .A(n5941), .B(n5942), .Z(n5944) );
  OR U6628 ( .A(n5910), .B(n5909), .Z(n5914) );
  NANDN U6629 ( .A(n5912), .B(n5911), .Z(n5913) );
  NAND U6630 ( .A(n5914), .B(n5913), .Z(n5943) );
  XNOR U6631 ( .A(n5944), .B(n5943), .Z(n5929) );
  NANDN U6632 ( .A(n5916), .B(n5915), .Z(n5920) );
  OR U6633 ( .A(n5918), .B(n5917), .Z(n5919) );
  NAND U6634 ( .A(n5920), .B(n5919), .Z(n5930) );
  XNOR U6635 ( .A(n5929), .B(n5930), .Z(n5931) );
  XOR U6636 ( .A(n5932), .B(n5931), .Z(n5928) );
  OR U6637 ( .A(n5921), .B(sreg[1210]), .Z(n5925) );
  NANDN U6638 ( .A(n5923), .B(n5922), .Z(n5924) );
  AND U6639 ( .A(n5925), .B(n5924), .Z(n5927) );
  XNOR U6640 ( .A(sreg[1211]), .B(n5927), .Z(n5926) );
  XOR U6641 ( .A(n5928), .B(n5926), .Z(c[1211]) );
  NANDN U6642 ( .A(n5930), .B(n5929), .Z(n5934) );
  NAND U6643 ( .A(n5932), .B(n5931), .Z(n5933) );
  NAND U6644 ( .A(n5934), .B(n5933), .Z(n5950) );
  AND U6645 ( .A(b[2]), .B(a[190]), .Z(n5956) );
  AND U6646 ( .A(a[191]), .B(b[1]), .Z(n5954) );
  AND U6647 ( .A(a[189]), .B(b[3]), .Z(n5953) );
  XOR U6648 ( .A(n5954), .B(n5953), .Z(n5955) );
  XOR U6649 ( .A(n5956), .B(n5955), .Z(n5959) );
  NAND U6650 ( .A(b[0]), .B(a[192]), .Z(n5960) );
  XOR U6651 ( .A(n5959), .B(n5960), .Z(n5962) );
  OR U6652 ( .A(n5936), .B(n5935), .Z(n5940) );
  NANDN U6653 ( .A(n5938), .B(n5937), .Z(n5939) );
  NAND U6654 ( .A(n5940), .B(n5939), .Z(n5961) );
  XNOR U6655 ( .A(n5962), .B(n5961), .Z(n5947) );
  NANDN U6656 ( .A(n5942), .B(n5941), .Z(n5946) );
  OR U6657 ( .A(n5944), .B(n5943), .Z(n5945) );
  NAND U6658 ( .A(n5946), .B(n5945), .Z(n5948) );
  XNOR U6659 ( .A(n5947), .B(n5948), .Z(n5949) );
  XNOR U6660 ( .A(n5950), .B(n5949), .Z(n5965) );
  XNOR U6661 ( .A(n5965), .B(sreg[1212]), .Z(n5966) );
  XOR U6662 ( .A(n5967), .B(n5966), .Z(c[1212]) );
  NANDN U6663 ( .A(n5948), .B(n5947), .Z(n5952) );
  NAND U6664 ( .A(n5950), .B(n5949), .Z(n5951) );
  NAND U6665 ( .A(n5952), .B(n5951), .Z(n5974) );
  AND U6666 ( .A(b[2]), .B(a[191]), .Z(n5980) );
  AND U6667 ( .A(a[192]), .B(b[1]), .Z(n5978) );
  AND U6668 ( .A(a[190]), .B(b[3]), .Z(n5977) );
  XOR U6669 ( .A(n5978), .B(n5977), .Z(n5979) );
  XOR U6670 ( .A(n5980), .B(n5979), .Z(n5983) );
  NAND U6671 ( .A(b[0]), .B(a[193]), .Z(n5984) );
  XOR U6672 ( .A(n5983), .B(n5984), .Z(n5986) );
  OR U6673 ( .A(n5954), .B(n5953), .Z(n5958) );
  NANDN U6674 ( .A(n5956), .B(n5955), .Z(n5957) );
  NAND U6675 ( .A(n5958), .B(n5957), .Z(n5985) );
  XNOR U6676 ( .A(n5986), .B(n5985), .Z(n5971) );
  NANDN U6677 ( .A(n5960), .B(n5959), .Z(n5964) );
  OR U6678 ( .A(n5962), .B(n5961), .Z(n5963) );
  NAND U6679 ( .A(n5964), .B(n5963), .Z(n5972) );
  XNOR U6680 ( .A(n5971), .B(n5972), .Z(n5973) );
  XOR U6681 ( .A(n5974), .B(n5973), .Z(n5990) );
  NAND U6682 ( .A(n5965), .B(sreg[1212]), .Z(n5969) );
  OR U6683 ( .A(n5967), .B(n5966), .Z(n5968) );
  NAND U6684 ( .A(n5969), .B(n5968), .Z(n5989) );
  XNOR U6685 ( .A(sreg[1213]), .B(n5989), .Z(n5970) );
  XOR U6686 ( .A(n5990), .B(n5970), .Z(c[1213]) );
  NANDN U6687 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U6688 ( .A(n5974), .B(n5973), .Z(n5975) );
  NAND U6689 ( .A(n5976), .B(n5975), .Z(n5995) );
  AND U6690 ( .A(b[2]), .B(a[192]), .Z(n6001) );
  AND U6691 ( .A(a[193]), .B(b[1]), .Z(n5999) );
  AND U6692 ( .A(a[191]), .B(b[3]), .Z(n5998) );
  XOR U6693 ( .A(n5999), .B(n5998), .Z(n6000) );
  XOR U6694 ( .A(n6001), .B(n6000), .Z(n6004) );
  NAND U6695 ( .A(b[0]), .B(a[194]), .Z(n6005) );
  XOR U6696 ( .A(n6004), .B(n6005), .Z(n6007) );
  OR U6697 ( .A(n5978), .B(n5977), .Z(n5982) );
  NANDN U6698 ( .A(n5980), .B(n5979), .Z(n5981) );
  NAND U6699 ( .A(n5982), .B(n5981), .Z(n6006) );
  XNOR U6700 ( .A(n6007), .B(n6006), .Z(n5992) );
  NANDN U6701 ( .A(n5984), .B(n5983), .Z(n5988) );
  OR U6702 ( .A(n5986), .B(n5985), .Z(n5987) );
  NAND U6703 ( .A(n5988), .B(n5987), .Z(n5993) );
  XNOR U6704 ( .A(n5992), .B(n5993), .Z(n5994) );
  XOR U6705 ( .A(n5995), .B(n5994), .Z(n6011) );
  XNOR U6706 ( .A(sreg[1214]), .B(n6010), .Z(n5991) );
  XOR U6707 ( .A(n6011), .B(n5991), .Z(c[1214]) );
  NANDN U6708 ( .A(n5993), .B(n5992), .Z(n5997) );
  NAND U6709 ( .A(n5995), .B(n5994), .Z(n5996) );
  NAND U6710 ( .A(n5997), .B(n5996), .Z(n6016) );
  AND U6711 ( .A(b[2]), .B(a[193]), .Z(n6022) );
  AND U6712 ( .A(a[194]), .B(b[1]), .Z(n6020) );
  AND U6713 ( .A(a[192]), .B(b[3]), .Z(n6019) );
  XOR U6714 ( .A(n6020), .B(n6019), .Z(n6021) );
  XOR U6715 ( .A(n6022), .B(n6021), .Z(n6025) );
  NAND U6716 ( .A(b[0]), .B(a[195]), .Z(n6026) );
  XOR U6717 ( .A(n6025), .B(n6026), .Z(n6028) );
  OR U6718 ( .A(n5999), .B(n5998), .Z(n6003) );
  NANDN U6719 ( .A(n6001), .B(n6000), .Z(n6002) );
  NAND U6720 ( .A(n6003), .B(n6002), .Z(n6027) );
  XNOR U6721 ( .A(n6028), .B(n6027), .Z(n6013) );
  NANDN U6722 ( .A(n6005), .B(n6004), .Z(n6009) );
  OR U6723 ( .A(n6007), .B(n6006), .Z(n6008) );
  NAND U6724 ( .A(n6009), .B(n6008), .Z(n6014) );
  XNOR U6725 ( .A(n6013), .B(n6014), .Z(n6015) );
  XOR U6726 ( .A(n6016), .B(n6015), .Z(n6032) );
  XNOR U6727 ( .A(sreg[1215]), .B(n6031), .Z(n6012) );
  XOR U6728 ( .A(n6032), .B(n6012), .Z(c[1215]) );
  NANDN U6729 ( .A(n6014), .B(n6013), .Z(n6018) );
  NAND U6730 ( .A(n6016), .B(n6015), .Z(n6017) );
  NAND U6731 ( .A(n6018), .B(n6017), .Z(n6039) );
  AND U6732 ( .A(b[2]), .B(a[194]), .Z(n6051) );
  AND U6733 ( .A(a[195]), .B(b[1]), .Z(n6049) );
  AND U6734 ( .A(a[193]), .B(b[3]), .Z(n6048) );
  XOR U6735 ( .A(n6049), .B(n6048), .Z(n6050) );
  XOR U6736 ( .A(n6051), .B(n6050), .Z(n6042) );
  NAND U6737 ( .A(b[0]), .B(a[196]), .Z(n6043) );
  XOR U6738 ( .A(n6042), .B(n6043), .Z(n6045) );
  OR U6739 ( .A(n6020), .B(n6019), .Z(n6024) );
  NANDN U6740 ( .A(n6022), .B(n6021), .Z(n6023) );
  NAND U6741 ( .A(n6024), .B(n6023), .Z(n6044) );
  XNOR U6742 ( .A(n6045), .B(n6044), .Z(n6036) );
  NANDN U6743 ( .A(n6026), .B(n6025), .Z(n6030) );
  OR U6744 ( .A(n6028), .B(n6027), .Z(n6029) );
  NAND U6745 ( .A(n6030), .B(n6029), .Z(n6037) );
  XNOR U6746 ( .A(n6036), .B(n6037), .Z(n6038) );
  XNOR U6747 ( .A(n6039), .B(n6038), .Z(n6035) );
  XOR U6748 ( .A(n6034), .B(sreg[1216]), .Z(n6033) );
  XOR U6749 ( .A(n6035), .B(n6033), .Z(c[1216]) );
  NANDN U6750 ( .A(n6037), .B(n6036), .Z(n6041) );
  NAND U6751 ( .A(n6039), .B(n6038), .Z(n6040) );
  NAND U6752 ( .A(n6041), .B(n6040), .Z(n6069) );
  NANDN U6753 ( .A(n6043), .B(n6042), .Z(n6047) );
  OR U6754 ( .A(n6045), .B(n6044), .Z(n6046) );
  NAND U6755 ( .A(n6047), .B(n6046), .Z(n6066) );
  AND U6756 ( .A(b[2]), .B(a[195]), .Z(n6057) );
  AND U6757 ( .A(a[196]), .B(b[1]), .Z(n6055) );
  AND U6758 ( .A(a[194]), .B(b[3]), .Z(n6054) );
  XOR U6759 ( .A(n6055), .B(n6054), .Z(n6056) );
  XOR U6760 ( .A(n6057), .B(n6056), .Z(n6060) );
  NAND U6761 ( .A(b[0]), .B(a[197]), .Z(n6061) );
  XNOR U6762 ( .A(n6060), .B(n6061), .Z(n6062) );
  OR U6763 ( .A(n6049), .B(n6048), .Z(n6053) );
  NANDN U6764 ( .A(n6051), .B(n6050), .Z(n6052) );
  AND U6765 ( .A(n6053), .B(n6052), .Z(n6063) );
  XNOR U6766 ( .A(n6062), .B(n6063), .Z(n6067) );
  XNOR U6767 ( .A(n6066), .B(n6067), .Z(n6068) );
  XNOR U6768 ( .A(n6069), .B(n6068), .Z(n6072) );
  XNOR U6769 ( .A(sreg[1217]), .B(n6072), .Z(n6074) );
  XNOR U6770 ( .A(n6073), .B(n6074), .Z(c[1217]) );
  AND U6771 ( .A(b[2]), .B(a[196]), .Z(n6089) );
  AND U6772 ( .A(a[197]), .B(b[1]), .Z(n6087) );
  AND U6773 ( .A(a[195]), .B(b[3]), .Z(n6086) );
  XOR U6774 ( .A(n6087), .B(n6086), .Z(n6088) );
  XOR U6775 ( .A(n6089), .B(n6088), .Z(n6092) );
  NAND U6776 ( .A(b[0]), .B(a[198]), .Z(n6093) );
  XOR U6777 ( .A(n6092), .B(n6093), .Z(n6095) );
  OR U6778 ( .A(n6055), .B(n6054), .Z(n6059) );
  NANDN U6779 ( .A(n6057), .B(n6056), .Z(n6058) );
  NAND U6780 ( .A(n6059), .B(n6058), .Z(n6094) );
  XNOR U6781 ( .A(n6095), .B(n6094), .Z(n6080) );
  NANDN U6782 ( .A(n6061), .B(n6060), .Z(n6065) );
  NAND U6783 ( .A(n6063), .B(n6062), .Z(n6064) );
  NAND U6784 ( .A(n6065), .B(n6064), .Z(n6081) );
  XNOR U6785 ( .A(n6080), .B(n6081), .Z(n6082) );
  NANDN U6786 ( .A(n6067), .B(n6066), .Z(n6071) );
  NANDN U6787 ( .A(n6069), .B(n6068), .Z(n6070) );
  NAND U6788 ( .A(n6071), .B(n6070), .Z(n6083) );
  XOR U6789 ( .A(n6082), .B(n6083), .Z(n6079) );
  NAND U6790 ( .A(sreg[1217]), .B(n6072), .Z(n6076) );
  NANDN U6791 ( .A(n6074), .B(n6073), .Z(n6075) );
  NAND U6792 ( .A(n6076), .B(n6075), .Z(n6078) );
  XNOR U6793 ( .A(sreg[1218]), .B(n6078), .Z(n6077) );
  XNOR U6794 ( .A(n6079), .B(n6077), .Z(c[1218]) );
  NANDN U6795 ( .A(n6081), .B(n6080), .Z(n6085) );
  NANDN U6796 ( .A(n6083), .B(n6082), .Z(n6084) );
  NAND U6797 ( .A(n6085), .B(n6084), .Z(n6113) );
  AND U6798 ( .A(b[2]), .B(a[197]), .Z(n6107) );
  AND U6799 ( .A(a[198]), .B(b[1]), .Z(n6105) );
  AND U6800 ( .A(a[196]), .B(b[3]), .Z(n6104) );
  XOR U6801 ( .A(n6105), .B(n6104), .Z(n6106) );
  XOR U6802 ( .A(n6107), .B(n6106), .Z(n6098) );
  NAND U6803 ( .A(b[0]), .B(a[199]), .Z(n6099) );
  XOR U6804 ( .A(n6098), .B(n6099), .Z(n6101) );
  OR U6805 ( .A(n6087), .B(n6086), .Z(n6091) );
  NANDN U6806 ( .A(n6089), .B(n6088), .Z(n6090) );
  NAND U6807 ( .A(n6091), .B(n6090), .Z(n6100) );
  XNOR U6808 ( .A(n6101), .B(n6100), .Z(n6110) );
  NANDN U6809 ( .A(n6093), .B(n6092), .Z(n6097) );
  OR U6810 ( .A(n6095), .B(n6094), .Z(n6096) );
  NAND U6811 ( .A(n6097), .B(n6096), .Z(n6111) );
  XNOR U6812 ( .A(n6110), .B(n6111), .Z(n6112) );
  XNOR U6813 ( .A(n6113), .B(n6112), .Z(n6116) );
  XNOR U6814 ( .A(n6116), .B(sreg[1219]), .Z(n6117) );
  XOR U6815 ( .A(n6118), .B(n6117), .Z(c[1219]) );
  NANDN U6816 ( .A(n6099), .B(n6098), .Z(n6103) );
  OR U6817 ( .A(n6101), .B(n6100), .Z(n6102) );
  NAND U6818 ( .A(n6103), .B(n6102), .Z(n6136) );
  AND U6819 ( .A(b[2]), .B(a[198]), .Z(n6127) );
  AND U6820 ( .A(a[199]), .B(b[1]), .Z(n6125) );
  AND U6821 ( .A(a[197]), .B(b[3]), .Z(n6124) );
  XOR U6822 ( .A(n6125), .B(n6124), .Z(n6126) );
  XOR U6823 ( .A(n6127), .B(n6126), .Z(n6130) );
  NAND U6824 ( .A(b[0]), .B(a[200]), .Z(n6131) );
  XNOR U6825 ( .A(n6130), .B(n6131), .Z(n6132) );
  OR U6826 ( .A(n6105), .B(n6104), .Z(n6109) );
  NANDN U6827 ( .A(n6107), .B(n6106), .Z(n6108) );
  AND U6828 ( .A(n6109), .B(n6108), .Z(n6133) );
  XNOR U6829 ( .A(n6132), .B(n6133), .Z(n6137) );
  XNOR U6830 ( .A(n6136), .B(n6137), .Z(n6138) );
  NANDN U6831 ( .A(n6111), .B(n6110), .Z(n6115) );
  NAND U6832 ( .A(n6113), .B(n6112), .Z(n6114) );
  NAND U6833 ( .A(n6115), .B(n6114), .Z(n6139) );
  XOR U6834 ( .A(n6138), .B(n6139), .Z(n6123) );
  NAND U6835 ( .A(n6116), .B(sreg[1219]), .Z(n6120) );
  OR U6836 ( .A(n6118), .B(n6117), .Z(n6119) );
  AND U6837 ( .A(n6120), .B(n6119), .Z(n6122) );
  XNOR U6838 ( .A(n6122), .B(sreg[1220]), .Z(n6121) );
  XNOR U6839 ( .A(n6123), .B(n6121), .Z(c[1220]) );
  AND U6840 ( .A(b[2]), .B(a[199]), .Z(n6151) );
  AND U6841 ( .A(a[200]), .B(b[1]), .Z(n6149) );
  AND U6842 ( .A(a[198]), .B(b[3]), .Z(n6148) );
  XOR U6843 ( .A(n6149), .B(n6148), .Z(n6150) );
  XOR U6844 ( .A(n6151), .B(n6150), .Z(n6154) );
  NAND U6845 ( .A(b[0]), .B(a[201]), .Z(n6155) );
  XOR U6846 ( .A(n6154), .B(n6155), .Z(n6157) );
  OR U6847 ( .A(n6125), .B(n6124), .Z(n6129) );
  NANDN U6848 ( .A(n6127), .B(n6126), .Z(n6128) );
  NAND U6849 ( .A(n6129), .B(n6128), .Z(n6156) );
  XNOR U6850 ( .A(n6157), .B(n6156), .Z(n6142) );
  NANDN U6851 ( .A(n6131), .B(n6130), .Z(n6135) );
  NAND U6852 ( .A(n6133), .B(n6132), .Z(n6134) );
  NAND U6853 ( .A(n6135), .B(n6134), .Z(n6143) );
  XNOR U6854 ( .A(n6142), .B(n6143), .Z(n6144) );
  NANDN U6855 ( .A(n6137), .B(n6136), .Z(n6141) );
  NANDN U6856 ( .A(n6139), .B(n6138), .Z(n6140) );
  NAND U6857 ( .A(n6141), .B(n6140), .Z(n6145) );
  XNOR U6858 ( .A(n6144), .B(n6145), .Z(n6160) );
  XOR U6859 ( .A(sreg[1221]), .B(n6160), .Z(n6162) );
  XNOR U6860 ( .A(n6161), .B(n6162), .Z(c[1221]) );
  NANDN U6861 ( .A(n6143), .B(n6142), .Z(n6147) );
  NANDN U6862 ( .A(n6145), .B(n6144), .Z(n6146) );
  NAND U6863 ( .A(n6147), .B(n6146), .Z(n6183) );
  AND U6864 ( .A(b[2]), .B(a[200]), .Z(n6177) );
  AND U6865 ( .A(a[201]), .B(b[1]), .Z(n6175) );
  AND U6866 ( .A(a[199]), .B(b[3]), .Z(n6174) );
  XOR U6867 ( .A(n6175), .B(n6174), .Z(n6176) );
  XOR U6868 ( .A(n6177), .B(n6176), .Z(n6168) );
  NAND U6869 ( .A(b[0]), .B(a[202]), .Z(n6169) );
  XOR U6870 ( .A(n6168), .B(n6169), .Z(n6171) );
  OR U6871 ( .A(n6149), .B(n6148), .Z(n6153) );
  NANDN U6872 ( .A(n6151), .B(n6150), .Z(n6152) );
  NAND U6873 ( .A(n6153), .B(n6152), .Z(n6170) );
  XNOR U6874 ( .A(n6171), .B(n6170), .Z(n6180) );
  NANDN U6875 ( .A(n6155), .B(n6154), .Z(n6159) );
  OR U6876 ( .A(n6157), .B(n6156), .Z(n6158) );
  NAND U6877 ( .A(n6159), .B(n6158), .Z(n6181) );
  XNOR U6878 ( .A(n6180), .B(n6181), .Z(n6182) );
  XOR U6879 ( .A(n6183), .B(n6182), .Z(n6167) );
  NANDN U6880 ( .A(n6160), .B(sreg[1221]), .Z(n6164) );
  NANDN U6881 ( .A(n6162), .B(n6161), .Z(n6163) );
  NAND U6882 ( .A(n6164), .B(n6163), .Z(n6166) );
  XNOR U6883 ( .A(sreg[1222]), .B(n6166), .Z(n6165) );
  XOR U6884 ( .A(n6167), .B(n6165), .Z(c[1222]) );
  NANDN U6885 ( .A(n6169), .B(n6168), .Z(n6173) );
  OR U6886 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U6887 ( .A(n6173), .B(n6172), .Z(n6198) );
  AND U6888 ( .A(b[2]), .B(a[201]), .Z(n6189) );
  AND U6889 ( .A(a[202]), .B(b[1]), .Z(n6187) );
  AND U6890 ( .A(a[200]), .B(b[3]), .Z(n6186) );
  XOR U6891 ( .A(n6187), .B(n6186), .Z(n6188) );
  XOR U6892 ( .A(n6189), .B(n6188), .Z(n6192) );
  NAND U6893 ( .A(b[0]), .B(a[203]), .Z(n6193) );
  XNOR U6894 ( .A(n6192), .B(n6193), .Z(n6194) );
  OR U6895 ( .A(n6175), .B(n6174), .Z(n6179) );
  NANDN U6896 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U6897 ( .A(n6179), .B(n6178), .Z(n6195) );
  XNOR U6898 ( .A(n6194), .B(n6195), .Z(n6199) );
  XNOR U6899 ( .A(n6198), .B(n6199), .Z(n6200) );
  NANDN U6900 ( .A(n6181), .B(n6180), .Z(n6185) );
  NAND U6901 ( .A(n6183), .B(n6182), .Z(n6184) );
  AND U6902 ( .A(n6185), .B(n6184), .Z(n6201) );
  XOR U6903 ( .A(n6200), .B(n6201), .Z(n6204) );
  XNOR U6904 ( .A(sreg[1223]), .B(n6204), .Z(n6205) );
  XOR U6905 ( .A(n6206), .B(n6205), .Z(c[1223]) );
  AND U6906 ( .A(b[2]), .B(a[202]), .Z(n6219) );
  AND U6907 ( .A(a[203]), .B(b[1]), .Z(n6217) );
  AND U6908 ( .A(a[201]), .B(b[3]), .Z(n6216) );
  XOR U6909 ( .A(n6217), .B(n6216), .Z(n6218) );
  XOR U6910 ( .A(n6219), .B(n6218), .Z(n6222) );
  NAND U6911 ( .A(b[0]), .B(a[204]), .Z(n6223) );
  XOR U6912 ( .A(n6222), .B(n6223), .Z(n6225) );
  OR U6913 ( .A(n6187), .B(n6186), .Z(n6191) );
  NANDN U6914 ( .A(n6189), .B(n6188), .Z(n6190) );
  NAND U6915 ( .A(n6191), .B(n6190), .Z(n6224) );
  XNOR U6916 ( .A(n6225), .B(n6224), .Z(n6210) );
  NANDN U6917 ( .A(n6193), .B(n6192), .Z(n6197) );
  NAND U6918 ( .A(n6195), .B(n6194), .Z(n6196) );
  NAND U6919 ( .A(n6197), .B(n6196), .Z(n6211) );
  XNOR U6920 ( .A(n6210), .B(n6211), .Z(n6212) );
  NANDN U6921 ( .A(n6199), .B(n6198), .Z(n6203) );
  NAND U6922 ( .A(n6201), .B(n6200), .Z(n6202) );
  AND U6923 ( .A(n6203), .B(n6202), .Z(n6213) );
  XNOR U6924 ( .A(n6212), .B(n6213), .Z(n6229) );
  NAND U6925 ( .A(sreg[1223]), .B(n6204), .Z(n6208) );
  OR U6926 ( .A(n6206), .B(n6205), .Z(n6207) );
  AND U6927 ( .A(n6208), .B(n6207), .Z(n6228) );
  XNOR U6928 ( .A(n6228), .B(sreg[1224]), .Z(n6209) );
  XOR U6929 ( .A(n6229), .B(n6209), .Z(c[1224]) );
  NANDN U6930 ( .A(n6211), .B(n6210), .Z(n6215) );
  NAND U6931 ( .A(n6213), .B(n6212), .Z(n6214) );
  NAND U6932 ( .A(n6215), .B(n6214), .Z(n6248) );
  AND U6933 ( .A(b[2]), .B(a[203]), .Z(n6242) );
  AND U6934 ( .A(a[204]), .B(b[1]), .Z(n6240) );
  AND U6935 ( .A(a[202]), .B(b[3]), .Z(n6239) );
  XOR U6936 ( .A(n6240), .B(n6239), .Z(n6241) );
  XOR U6937 ( .A(n6242), .B(n6241), .Z(n6233) );
  NAND U6938 ( .A(b[0]), .B(a[205]), .Z(n6234) );
  XOR U6939 ( .A(n6233), .B(n6234), .Z(n6236) );
  OR U6940 ( .A(n6217), .B(n6216), .Z(n6221) );
  NANDN U6941 ( .A(n6219), .B(n6218), .Z(n6220) );
  NAND U6942 ( .A(n6221), .B(n6220), .Z(n6235) );
  XNOR U6943 ( .A(n6236), .B(n6235), .Z(n6245) );
  NANDN U6944 ( .A(n6223), .B(n6222), .Z(n6227) );
  OR U6945 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U6946 ( .A(n6227), .B(n6226), .Z(n6246) );
  XNOR U6947 ( .A(n6245), .B(n6246), .Z(n6247) );
  XOR U6948 ( .A(n6248), .B(n6247), .Z(n6232) );
  XOR U6949 ( .A(sreg[1225]), .B(n6231), .Z(n6230) );
  XOR U6950 ( .A(n6232), .B(n6230), .Z(c[1225]) );
  NANDN U6951 ( .A(n6234), .B(n6233), .Z(n6238) );
  OR U6952 ( .A(n6236), .B(n6235), .Z(n6237) );
  NAND U6953 ( .A(n6238), .B(n6237), .Z(n6268) );
  AND U6954 ( .A(b[2]), .B(a[204]), .Z(n6259) );
  AND U6955 ( .A(a[205]), .B(b[1]), .Z(n6257) );
  AND U6956 ( .A(a[203]), .B(b[3]), .Z(n6256) );
  XOR U6957 ( .A(n6257), .B(n6256), .Z(n6258) );
  XOR U6958 ( .A(n6259), .B(n6258), .Z(n6262) );
  NAND U6959 ( .A(b[0]), .B(a[206]), .Z(n6263) );
  XNOR U6960 ( .A(n6262), .B(n6263), .Z(n6264) );
  OR U6961 ( .A(n6240), .B(n6239), .Z(n6244) );
  NANDN U6962 ( .A(n6242), .B(n6241), .Z(n6243) );
  AND U6963 ( .A(n6244), .B(n6243), .Z(n6265) );
  XNOR U6964 ( .A(n6264), .B(n6265), .Z(n6269) );
  XNOR U6965 ( .A(n6268), .B(n6269), .Z(n6270) );
  NANDN U6966 ( .A(n6246), .B(n6245), .Z(n6250) );
  NAND U6967 ( .A(n6248), .B(n6247), .Z(n6249) );
  AND U6968 ( .A(n6250), .B(n6249), .Z(n6271) );
  XOR U6969 ( .A(n6270), .B(n6271), .Z(n6251) );
  XNOR U6970 ( .A(sreg[1226]), .B(n6251), .Z(n6252) );
  XOR U6971 ( .A(n6253), .B(n6252), .Z(c[1226]) );
  NAND U6972 ( .A(sreg[1226]), .B(n6251), .Z(n6255) );
  OR U6973 ( .A(n6253), .B(n6252), .Z(n6254) );
  AND U6974 ( .A(n6255), .B(n6254), .Z(n6295) );
  IV U6975 ( .A(sreg[1227]), .Z(n6293) );
  AND U6976 ( .A(b[2]), .B(a[205]), .Z(n6284) );
  AND U6977 ( .A(a[206]), .B(b[1]), .Z(n6282) );
  AND U6978 ( .A(a[204]), .B(b[3]), .Z(n6281) );
  XOR U6979 ( .A(n6282), .B(n6281), .Z(n6283) );
  XOR U6980 ( .A(n6284), .B(n6283), .Z(n6287) );
  NAND U6981 ( .A(b[0]), .B(a[207]), .Z(n6288) );
  XOR U6982 ( .A(n6287), .B(n6288), .Z(n6290) );
  OR U6983 ( .A(n6257), .B(n6256), .Z(n6261) );
  NANDN U6984 ( .A(n6259), .B(n6258), .Z(n6260) );
  NAND U6985 ( .A(n6261), .B(n6260), .Z(n6289) );
  XNOR U6986 ( .A(n6290), .B(n6289), .Z(n6275) );
  NANDN U6987 ( .A(n6263), .B(n6262), .Z(n6267) );
  NAND U6988 ( .A(n6265), .B(n6264), .Z(n6266) );
  NAND U6989 ( .A(n6267), .B(n6266), .Z(n6276) );
  XNOR U6990 ( .A(n6275), .B(n6276), .Z(n6277) );
  NANDN U6991 ( .A(n6269), .B(n6268), .Z(n6273) );
  NAND U6992 ( .A(n6271), .B(n6270), .Z(n6272) );
  NAND U6993 ( .A(n6273), .B(n6272), .Z(n6278) );
  XOR U6994 ( .A(n6277), .B(n6278), .Z(n6294) );
  XOR U6995 ( .A(n6293), .B(n6294), .Z(n6274) );
  XOR U6996 ( .A(n6295), .B(n6274), .Z(c[1227]) );
  NANDN U6997 ( .A(n6276), .B(n6275), .Z(n6280) );
  NANDN U6998 ( .A(n6278), .B(n6277), .Z(n6279) );
  NAND U6999 ( .A(n6280), .B(n6279), .Z(n6305) );
  AND U7000 ( .A(b[2]), .B(a[206]), .Z(n6311) );
  AND U7001 ( .A(a[207]), .B(b[1]), .Z(n6309) );
  AND U7002 ( .A(a[205]), .B(b[3]), .Z(n6308) );
  XOR U7003 ( .A(n6309), .B(n6308), .Z(n6310) );
  XOR U7004 ( .A(n6311), .B(n6310), .Z(n6314) );
  NAND U7005 ( .A(b[0]), .B(a[208]), .Z(n6315) );
  XOR U7006 ( .A(n6314), .B(n6315), .Z(n6317) );
  OR U7007 ( .A(n6282), .B(n6281), .Z(n6286) );
  NANDN U7008 ( .A(n6284), .B(n6283), .Z(n6285) );
  NAND U7009 ( .A(n6286), .B(n6285), .Z(n6316) );
  XNOR U7010 ( .A(n6317), .B(n6316), .Z(n6302) );
  NANDN U7011 ( .A(n6288), .B(n6287), .Z(n6292) );
  OR U7012 ( .A(n6290), .B(n6289), .Z(n6291) );
  NAND U7013 ( .A(n6292), .B(n6291), .Z(n6303) );
  XNOR U7014 ( .A(n6302), .B(n6303), .Z(n6304) );
  XOR U7015 ( .A(n6305), .B(n6304), .Z(n6301) );
  NANDN U7016 ( .A(n6294), .B(n6293), .Z(n6298) );
  AND U7017 ( .A(n6294), .B(sreg[1227]), .Z(n6296) );
  NANDN U7018 ( .A(n6296), .B(n6295), .Z(n6297) );
  AND U7019 ( .A(n6298), .B(n6297), .Z(n6300) );
  XNOR U7020 ( .A(sreg[1228]), .B(n6300), .Z(n6299) );
  XOR U7021 ( .A(n6301), .B(n6299), .Z(c[1228]) );
  NANDN U7022 ( .A(n6303), .B(n6302), .Z(n6307) );
  NAND U7023 ( .A(n6305), .B(n6304), .Z(n6306) );
  NAND U7024 ( .A(n6307), .B(n6306), .Z(n6323) );
  AND U7025 ( .A(b[2]), .B(a[207]), .Z(n6329) );
  AND U7026 ( .A(a[208]), .B(b[1]), .Z(n6327) );
  AND U7027 ( .A(a[206]), .B(b[3]), .Z(n6326) );
  XOR U7028 ( .A(n6327), .B(n6326), .Z(n6328) );
  XOR U7029 ( .A(n6329), .B(n6328), .Z(n6332) );
  NAND U7030 ( .A(b[0]), .B(a[209]), .Z(n6333) );
  XOR U7031 ( .A(n6332), .B(n6333), .Z(n6335) );
  OR U7032 ( .A(n6309), .B(n6308), .Z(n6313) );
  NANDN U7033 ( .A(n6311), .B(n6310), .Z(n6312) );
  NAND U7034 ( .A(n6313), .B(n6312), .Z(n6334) );
  XNOR U7035 ( .A(n6335), .B(n6334), .Z(n6320) );
  NANDN U7036 ( .A(n6315), .B(n6314), .Z(n6319) );
  OR U7037 ( .A(n6317), .B(n6316), .Z(n6318) );
  NAND U7038 ( .A(n6319), .B(n6318), .Z(n6321) );
  XNOR U7039 ( .A(n6320), .B(n6321), .Z(n6322) );
  XNOR U7040 ( .A(n6323), .B(n6322), .Z(n6338) );
  XNOR U7041 ( .A(n6338), .B(sreg[1229]), .Z(n6339) );
  XOR U7042 ( .A(n6340), .B(n6339), .Z(c[1229]) );
  NANDN U7043 ( .A(n6321), .B(n6320), .Z(n6325) );
  NAND U7044 ( .A(n6323), .B(n6322), .Z(n6324) );
  NAND U7045 ( .A(n6325), .B(n6324), .Z(n6349) );
  AND U7046 ( .A(b[2]), .B(a[208]), .Z(n6355) );
  AND U7047 ( .A(a[209]), .B(b[1]), .Z(n6353) );
  AND U7048 ( .A(a[207]), .B(b[3]), .Z(n6352) );
  XOR U7049 ( .A(n6353), .B(n6352), .Z(n6354) );
  XOR U7050 ( .A(n6355), .B(n6354), .Z(n6358) );
  NAND U7051 ( .A(b[0]), .B(a[210]), .Z(n6359) );
  XOR U7052 ( .A(n6358), .B(n6359), .Z(n6361) );
  OR U7053 ( .A(n6327), .B(n6326), .Z(n6331) );
  NANDN U7054 ( .A(n6329), .B(n6328), .Z(n6330) );
  NAND U7055 ( .A(n6331), .B(n6330), .Z(n6360) );
  XNOR U7056 ( .A(n6361), .B(n6360), .Z(n6346) );
  NANDN U7057 ( .A(n6333), .B(n6332), .Z(n6337) );
  OR U7058 ( .A(n6335), .B(n6334), .Z(n6336) );
  NAND U7059 ( .A(n6337), .B(n6336), .Z(n6347) );
  XNOR U7060 ( .A(n6346), .B(n6347), .Z(n6348) );
  XOR U7061 ( .A(n6349), .B(n6348), .Z(n6345) );
  NAND U7062 ( .A(n6338), .B(sreg[1229]), .Z(n6342) );
  OR U7063 ( .A(n6340), .B(n6339), .Z(n6341) );
  NAND U7064 ( .A(n6342), .B(n6341), .Z(n6344) );
  XNOR U7065 ( .A(sreg[1230]), .B(n6344), .Z(n6343) );
  XOR U7066 ( .A(n6345), .B(n6343), .Z(c[1230]) );
  NANDN U7067 ( .A(n6347), .B(n6346), .Z(n6351) );
  NAND U7068 ( .A(n6349), .B(n6348), .Z(n6350) );
  NAND U7069 ( .A(n6351), .B(n6350), .Z(n6367) );
  AND U7070 ( .A(b[2]), .B(a[209]), .Z(n6373) );
  AND U7071 ( .A(a[210]), .B(b[1]), .Z(n6371) );
  AND U7072 ( .A(a[208]), .B(b[3]), .Z(n6370) );
  XOR U7073 ( .A(n6371), .B(n6370), .Z(n6372) );
  XOR U7074 ( .A(n6373), .B(n6372), .Z(n6376) );
  NAND U7075 ( .A(b[0]), .B(a[211]), .Z(n6377) );
  XOR U7076 ( .A(n6376), .B(n6377), .Z(n6379) );
  OR U7077 ( .A(n6353), .B(n6352), .Z(n6357) );
  NANDN U7078 ( .A(n6355), .B(n6354), .Z(n6356) );
  NAND U7079 ( .A(n6357), .B(n6356), .Z(n6378) );
  XNOR U7080 ( .A(n6379), .B(n6378), .Z(n6364) );
  NANDN U7081 ( .A(n6359), .B(n6358), .Z(n6363) );
  OR U7082 ( .A(n6361), .B(n6360), .Z(n6362) );
  NAND U7083 ( .A(n6363), .B(n6362), .Z(n6365) );
  XNOR U7084 ( .A(n6364), .B(n6365), .Z(n6366) );
  XNOR U7085 ( .A(n6367), .B(n6366), .Z(n6382) );
  XNOR U7086 ( .A(n6382), .B(sreg[1231]), .Z(n6383) );
  XOR U7087 ( .A(n6384), .B(n6383), .Z(c[1231]) );
  NANDN U7088 ( .A(n6365), .B(n6364), .Z(n6369) );
  NAND U7089 ( .A(n6367), .B(n6366), .Z(n6368) );
  NAND U7090 ( .A(n6369), .B(n6368), .Z(n6395) );
  AND U7091 ( .A(b[2]), .B(a[210]), .Z(n6401) );
  AND U7092 ( .A(a[211]), .B(b[1]), .Z(n6399) );
  AND U7093 ( .A(a[209]), .B(b[3]), .Z(n6398) );
  XOR U7094 ( .A(n6399), .B(n6398), .Z(n6400) );
  XOR U7095 ( .A(n6401), .B(n6400), .Z(n6404) );
  NAND U7096 ( .A(b[0]), .B(a[212]), .Z(n6405) );
  XOR U7097 ( .A(n6404), .B(n6405), .Z(n6407) );
  OR U7098 ( .A(n6371), .B(n6370), .Z(n6375) );
  NANDN U7099 ( .A(n6373), .B(n6372), .Z(n6374) );
  NAND U7100 ( .A(n6375), .B(n6374), .Z(n6406) );
  XNOR U7101 ( .A(n6407), .B(n6406), .Z(n6392) );
  NANDN U7102 ( .A(n6377), .B(n6376), .Z(n6381) );
  OR U7103 ( .A(n6379), .B(n6378), .Z(n6380) );
  NAND U7104 ( .A(n6381), .B(n6380), .Z(n6393) );
  XNOR U7105 ( .A(n6392), .B(n6393), .Z(n6394) );
  XNOR U7106 ( .A(n6395), .B(n6394), .Z(n6387) );
  XOR U7107 ( .A(sreg[1232]), .B(n6387), .Z(n6388) );
  NAND U7108 ( .A(n6382), .B(sreg[1231]), .Z(n6386) );
  OR U7109 ( .A(n6384), .B(n6383), .Z(n6385) );
  NAND U7110 ( .A(n6386), .B(n6385), .Z(n6389) );
  XOR U7111 ( .A(n6388), .B(n6389), .Z(c[1232]) );
  OR U7112 ( .A(n6387), .B(sreg[1232]), .Z(n6391) );
  NANDN U7113 ( .A(n6389), .B(n6388), .Z(n6390) );
  AND U7114 ( .A(n6391), .B(n6390), .Z(n6429) );
  NANDN U7115 ( .A(n6393), .B(n6392), .Z(n6397) );
  NAND U7116 ( .A(n6395), .B(n6394), .Z(n6396) );
  NAND U7117 ( .A(n6397), .B(n6396), .Z(n6414) );
  AND U7118 ( .A(b[2]), .B(a[211]), .Z(n6420) );
  AND U7119 ( .A(a[212]), .B(b[1]), .Z(n6418) );
  AND U7120 ( .A(a[210]), .B(b[3]), .Z(n6417) );
  XOR U7121 ( .A(n6418), .B(n6417), .Z(n6419) );
  XOR U7122 ( .A(n6420), .B(n6419), .Z(n6423) );
  NAND U7123 ( .A(b[0]), .B(a[213]), .Z(n6424) );
  XOR U7124 ( .A(n6423), .B(n6424), .Z(n6426) );
  OR U7125 ( .A(n6399), .B(n6398), .Z(n6403) );
  NANDN U7126 ( .A(n6401), .B(n6400), .Z(n6402) );
  NAND U7127 ( .A(n6403), .B(n6402), .Z(n6425) );
  XNOR U7128 ( .A(n6426), .B(n6425), .Z(n6411) );
  NANDN U7129 ( .A(n6405), .B(n6404), .Z(n6409) );
  OR U7130 ( .A(n6407), .B(n6406), .Z(n6408) );
  NAND U7131 ( .A(n6409), .B(n6408), .Z(n6412) );
  XNOR U7132 ( .A(n6411), .B(n6412), .Z(n6413) );
  XNOR U7133 ( .A(n6414), .B(n6413), .Z(n6430) );
  XOR U7134 ( .A(sreg[1233]), .B(n6430), .Z(n6410) );
  XOR U7135 ( .A(n6429), .B(n6410), .Z(c[1233]) );
  NANDN U7136 ( .A(n6412), .B(n6411), .Z(n6416) );
  NAND U7137 ( .A(n6414), .B(n6413), .Z(n6415) );
  NAND U7138 ( .A(n6416), .B(n6415), .Z(n6437) );
  AND U7139 ( .A(b[2]), .B(a[212]), .Z(n6443) );
  AND U7140 ( .A(a[213]), .B(b[1]), .Z(n6441) );
  AND U7141 ( .A(a[211]), .B(b[3]), .Z(n6440) );
  XOR U7142 ( .A(n6441), .B(n6440), .Z(n6442) );
  XOR U7143 ( .A(n6443), .B(n6442), .Z(n6446) );
  NAND U7144 ( .A(b[0]), .B(a[214]), .Z(n6447) );
  XOR U7145 ( .A(n6446), .B(n6447), .Z(n6449) );
  OR U7146 ( .A(n6418), .B(n6417), .Z(n6422) );
  NANDN U7147 ( .A(n6420), .B(n6419), .Z(n6421) );
  NAND U7148 ( .A(n6422), .B(n6421), .Z(n6448) );
  XNOR U7149 ( .A(n6449), .B(n6448), .Z(n6434) );
  NANDN U7150 ( .A(n6424), .B(n6423), .Z(n6428) );
  OR U7151 ( .A(n6426), .B(n6425), .Z(n6427) );
  NAND U7152 ( .A(n6428), .B(n6427), .Z(n6435) );
  XNOR U7153 ( .A(n6434), .B(n6435), .Z(n6436) );
  XOR U7154 ( .A(n6437), .B(n6436), .Z(n6433) );
  XOR U7155 ( .A(sreg[1234]), .B(n6432), .Z(n6431) );
  XOR U7156 ( .A(n6433), .B(n6431), .Z(c[1234]) );
  NANDN U7157 ( .A(n6435), .B(n6434), .Z(n6439) );
  NAND U7158 ( .A(n6437), .B(n6436), .Z(n6438) );
  NAND U7159 ( .A(n6439), .B(n6438), .Z(n6455) );
  AND U7160 ( .A(b[2]), .B(a[213]), .Z(n6461) );
  AND U7161 ( .A(a[214]), .B(b[1]), .Z(n6459) );
  AND U7162 ( .A(a[212]), .B(b[3]), .Z(n6458) );
  XOR U7163 ( .A(n6459), .B(n6458), .Z(n6460) );
  XOR U7164 ( .A(n6461), .B(n6460), .Z(n6464) );
  NAND U7165 ( .A(b[0]), .B(a[215]), .Z(n6465) );
  XOR U7166 ( .A(n6464), .B(n6465), .Z(n6467) );
  OR U7167 ( .A(n6441), .B(n6440), .Z(n6445) );
  NANDN U7168 ( .A(n6443), .B(n6442), .Z(n6444) );
  NAND U7169 ( .A(n6445), .B(n6444), .Z(n6466) );
  XNOR U7170 ( .A(n6467), .B(n6466), .Z(n6452) );
  NANDN U7171 ( .A(n6447), .B(n6446), .Z(n6451) );
  OR U7172 ( .A(n6449), .B(n6448), .Z(n6450) );
  NAND U7173 ( .A(n6451), .B(n6450), .Z(n6453) );
  XNOR U7174 ( .A(n6452), .B(n6453), .Z(n6454) );
  XNOR U7175 ( .A(n6455), .B(n6454), .Z(n6470) );
  XNOR U7176 ( .A(n6470), .B(sreg[1235]), .Z(n6471) );
  XOR U7177 ( .A(n6472), .B(n6471), .Z(c[1235]) );
  NANDN U7178 ( .A(n6453), .B(n6452), .Z(n6457) );
  NAND U7179 ( .A(n6455), .B(n6454), .Z(n6456) );
  NAND U7180 ( .A(n6457), .B(n6456), .Z(n6478) );
  AND U7181 ( .A(b[2]), .B(a[214]), .Z(n6484) );
  AND U7182 ( .A(a[215]), .B(b[1]), .Z(n6482) );
  AND U7183 ( .A(a[213]), .B(b[3]), .Z(n6481) );
  XOR U7184 ( .A(n6482), .B(n6481), .Z(n6483) );
  XOR U7185 ( .A(n6484), .B(n6483), .Z(n6487) );
  NAND U7186 ( .A(b[0]), .B(a[216]), .Z(n6488) );
  XOR U7187 ( .A(n6487), .B(n6488), .Z(n6490) );
  OR U7188 ( .A(n6459), .B(n6458), .Z(n6463) );
  NANDN U7189 ( .A(n6461), .B(n6460), .Z(n6462) );
  NAND U7190 ( .A(n6463), .B(n6462), .Z(n6489) );
  XNOR U7191 ( .A(n6490), .B(n6489), .Z(n6475) );
  NANDN U7192 ( .A(n6465), .B(n6464), .Z(n6469) );
  OR U7193 ( .A(n6467), .B(n6466), .Z(n6468) );
  NAND U7194 ( .A(n6469), .B(n6468), .Z(n6476) );
  XNOR U7195 ( .A(n6475), .B(n6476), .Z(n6477) );
  XNOR U7196 ( .A(n6478), .B(n6477), .Z(n6493) );
  XNOR U7197 ( .A(n6493), .B(sreg[1236]), .Z(n6495) );
  NAND U7198 ( .A(n6470), .B(sreg[1235]), .Z(n6474) );
  OR U7199 ( .A(n6472), .B(n6471), .Z(n6473) );
  AND U7200 ( .A(n6474), .B(n6473), .Z(n6494) );
  XOR U7201 ( .A(n6495), .B(n6494), .Z(c[1236]) );
  NANDN U7202 ( .A(n6476), .B(n6475), .Z(n6480) );
  NAND U7203 ( .A(n6478), .B(n6477), .Z(n6479) );
  NAND U7204 ( .A(n6480), .B(n6479), .Z(n6504) );
  AND U7205 ( .A(b[2]), .B(a[215]), .Z(n6510) );
  AND U7206 ( .A(a[216]), .B(b[1]), .Z(n6508) );
  AND U7207 ( .A(a[214]), .B(b[3]), .Z(n6507) );
  XOR U7208 ( .A(n6508), .B(n6507), .Z(n6509) );
  XOR U7209 ( .A(n6510), .B(n6509), .Z(n6513) );
  NAND U7210 ( .A(b[0]), .B(a[217]), .Z(n6514) );
  XOR U7211 ( .A(n6513), .B(n6514), .Z(n6516) );
  OR U7212 ( .A(n6482), .B(n6481), .Z(n6486) );
  NANDN U7213 ( .A(n6484), .B(n6483), .Z(n6485) );
  NAND U7214 ( .A(n6486), .B(n6485), .Z(n6515) );
  XNOR U7215 ( .A(n6516), .B(n6515), .Z(n6501) );
  NANDN U7216 ( .A(n6488), .B(n6487), .Z(n6492) );
  OR U7217 ( .A(n6490), .B(n6489), .Z(n6491) );
  NAND U7218 ( .A(n6492), .B(n6491), .Z(n6502) );
  XNOR U7219 ( .A(n6501), .B(n6502), .Z(n6503) );
  XNOR U7220 ( .A(n6504), .B(n6503), .Z(n6500) );
  NAND U7221 ( .A(n6493), .B(sreg[1236]), .Z(n6497) );
  OR U7222 ( .A(n6495), .B(n6494), .Z(n6496) );
  AND U7223 ( .A(n6497), .B(n6496), .Z(n6499) );
  XNOR U7224 ( .A(n6499), .B(sreg[1237]), .Z(n6498) );
  XOR U7225 ( .A(n6500), .B(n6498), .Z(c[1237]) );
  NANDN U7226 ( .A(n6502), .B(n6501), .Z(n6506) );
  NAND U7227 ( .A(n6504), .B(n6503), .Z(n6505) );
  NAND U7228 ( .A(n6506), .B(n6505), .Z(n6522) );
  AND U7229 ( .A(b[2]), .B(a[216]), .Z(n6528) );
  AND U7230 ( .A(a[217]), .B(b[1]), .Z(n6526) );
  AND U7231 ( .A(a[215]), .B(b[3]), .Z(n6525) );
  XOR U7232 ( .A(n6526), .B(n6525), .Z(n6527) );
  XOR U7233 ( .A(n6528), .B(n6527), .Z(n6531) );
  NAND U7234 ( .A(b[0]), .B(a[218]), .Z(n6532) );
  XOR U7235 ( .A(n6531), .B(n6532), .Z(n6534) );
  OR U7236 ( .A(n6508), .B(n6507), .Z(n6512) );
  NANDN U7237 ( .A(n6510), .B(n6509), .Z(n6511) );
  NAND U7238 ( .A(n6512), .B(n6511), .Z(n6533) );
  XNOR U7239 ( .A(n6534), .B(n6533), .Z(n6519) );
  NANDN U7240 ( .A(n6514), .B(n6513), .Z(n6518) );
  OR U7241 ( .A(n6516), .B(n6515), .Z(n6517) );
  NAND U7242 ( .A(n6518), .B(n6517), .Z(n6520) );
  XNOR U7243 ( .A(n6519), .B(n6520), .Z(n6521) );
  XNOR U7244 ( .A(n6522), .B(n6521), .Z(n6537) );
  XNOR U7245 ( .A(n6537), .B(sreg[1238]), .Z(n6539) );
  XNOR U7246 ( .A(n6538), .B(n6539), .Z(c[1238]) );
  NANDN U7247 ( .A(n6520), .B(n6519), .Z(n6524) );
  NAND U7248 ( .A(n6522), .B(n6521), .Z(n6523) );
  NAND U7249 ( .A(n6524), .B(n6523), .Z(n6545) );
  AND U7250 ( .A(b[2]), .B(a[217]), .Z(n6557) );
  AND U7251 ( .A(a[218]), .B(b[1]), .Z(n6555) );
  AND U7252 ( .A(a[216]), .B(b[3]), .Z(n6554) );
  XOR U7253 ( .A(n6555), .B(n6554), .Z(n6556) );
  XOR U7254 ( .A(n6557), .B(n6556), .Z(n6548) );
  NAND U7255 ( .A(b[0]), .B(a[219]), .Z(n6549) );
  XOR U7256 ( .A(n6548), .B(n6549), .Z(n6551) );
  OR U7257 ( .A(n6526), .B(n6525), .Z(n6530) );
  NANDN U7258 ( .A(n6528), .B(n6527), .Z(n6529) );
  NAND U7259 ( .A(n6530), .B(n6529), .Z(n6550) );
  XNOR U7260 ( .A(n6551), .B(n6550), .Z(n6542) );
  NANDN U7261 ( .A(n6532), .B(n6531), .Z(n6536) );
  OR U7262 ( .A(n6534), .B(n6533), .Z(n6535) );
  NAND U7263 ( .A(n6536), .B(n6535), .Z(n6543) );
  XNOR U7264 ( .A(n6542), .B(n6543), .Z(n6544) );
  XNOR U7265 ( .A(n6545), .B(n6544), .Z(n6561) );
  XOR U7266 ( .A(sreg[1239]), .B(n6561), .Z(n6562) );
  NAND U7267 ( .A(n6537), .B(sreg[1238]), .Z(n6541) );
  NANDN U7268 ( .A(n6539), .B(n6538), .Z(n6540) );
  NAND U7269 ( .A(n6541), .B(n6540), .Z(n6563) );
  XOR U7270 ( .A(n6562), .B(n6563), .Z(c[1239]) );
  NANDN U7271 ( .A(n6543), .B(n6542), .Z(n6547) );
  NAND U7272 ( .A(n6545), .B(n6544), .Z(n6546) );
  NAND U7273 ( .A(n6547), .B(n6546), .Z(n6573) );
  NANDN U7274 ( .A(n6549), .B(n6548), .Z(n6553) );
  OR U7275 ( .A(n6551), .B(n6550), .Z(n6552) );
  AND U7276 ( .A(n6553), .B(n6552), .Z(n6572) );
  AND U7277 ( .A(b[2]), .B(a[218]), .Z(n6577) );
  AND U7278 ( .A(a[219]), .B(b[1]), .Z(n6575) );
  AND U7279 ( .A(a[217]), .B(b[3]), .Z(n6574) );
  XOR U7280 ( .A(n6575), .B(n6574), .Z(n6576) );
  XOR U7281 ( .A(n6577), .B(n6576), .Z(n6580) );
  NAND U7282 ( .A(b[0]), .B(a[220]), .Z(n6581) );
  XOR U7283 ( .A(n6580), .B(n6581), .Z(n6583) );
  OR U7284 ( .A(n6555), .B(n6554), .Z(n6559) );
  NANDN U7285 ( .A(n6557), .B(n6556), .Z(n6558) );
  NAND U7286 ( .A(n6559), .B(n6558), .Z(n6582) );
  XOR U7287 ( .A(n6583), .B(n6582), .Z(n6571) );
  XNOR U7288 ( .A(n6572), .B(n6571), .Z(n6560) );
  XNOR U7289 ( .A(n6573), .B(n6560), .Z(n6566) );
  XOR U7290 ( .A(sreg[1240]), .B(n6566), .Z(n6567) );
  OR U7291 ( .A(n6561), .B(sreg[1239]), .Z(n6565) );
  NANDN U7292 ( .A(n6563), .B(n6562), .Z(n6564) );
  AND U7293 ( .A(n6565), .B(n6564), .Z(n6568) );
  XOR U7294 ( .A(n6567), .B(n6568), .Z(c[1240]) );
  OR U7295 ( .A(n6566), .B(sreg[1240]), .Z(n6570) );
  NANDN U7296 ( .A(n6568), .B(n6567), .Z(n6569) );
  AND U7297 ( .A(n6570), .B(n6569), .Z(n6587) );
  AND U7298 ( .A(b[2]), .B(a[219]), .Z(n6598) );
  AND U7299 ( .A(a[220]), .B(b[1]), .Z(n6596) );
  AND U7300 ( .A(a[218]), .B(b[3]), .Z(n6595) );
  XOR U7301 ( .A(n6596), .B(n6595), .Z(n6597) );
  XOR U7302 ( .A(n6598), .B(n6597), .Z(n6601) );
  NAND U7303 ( .A(b[0]), .B(a[221]), .Z(n6602) );
  XOR U7304 ( .A(n6601), .B(n6602), .Z(n6604) );
  OR U7305 ( .A(n6575), .B(n6574), .Z(n6579) );
  NANDN U7306 ( .A(n6577), .B(n6576), .Z(n6578) );
  NAND U7307 ( .A(n6579), .B(n6578), .Z(n6603) );
  XNOR U7308 ( .A(n6604), .B(n6603), .Z(n6589) );
  NANDN U7309 ( .A(n6581), .B(n6580), .Z(n6585) );
  OR U7310 ( .A(n6583), .B(n6582), .Z(n6584) );
  NAND U7311 ( .A(n6585), .B(n6584), .Z(n6590) );
  XNOR U7312 ( .A(n6589), .B(n6590), .Z(n6591) );
  XNOR U7313 ( .A(n6592), .B(n6591), .Z(n6588) );
  XNOR U7314 ( .A(sreg[1241]), .B(n6588), .Z(n6586) );
  XOR U7315 ( .A(n6587), .B(n6586), .Z(c[1241]) );
  NANDN U7316 ( .A(n6590), .B(n6589), .Z(n6594) );
  NANDN U7317 ( .A(n6592), .B(n6591), .Z(n6593) );
  NAND U7318 ( .A(n6594), .B(n6593), .Z(n6610) );
  AND U7319 ( .A(b[2]), .B(a[220]), .Z(n6616) );
  AND U7320 ( .A(a[221]), .B(b[1]), .Z(n6614) );
  AND U7321 ( .A(a[219]), .B(b[3]), .Z(n6613) );
  XOR U7322 ( .A(n6614), .B(n6613), .Z(n6615) );
  XOR U7323 ( .A(n6616), .B(n6615), .Z(n6619) );
  NAND U7324 ( .A(b[0]), .B(a[222]), .Z(n6620) );
  XOR U7325 ( .A(n6619), .B(n6620), .Z(n6622) );
  OR U7326 ( .A(n6596), .B(n6595), .Z(n6600) );
  NANDN U7327 ( .A(n6598), .B(n6597), .Z(n6599) );
  NAND U7328 ( .A(n6600), .B(n6599), .Z(n6621) );
  XNOR U7329 ( .A(n6622), .B(n6621), .Z(n6607) );
  NANDN U7330 ( .A(n6602), .B(n6601), .Z(n6606) );
  OR U7331 ( .A(n6604), .B(n6603), .Z(n6605) );
  NAND U7332 ( .A(n6606), .B(n6605), .Z(n6608) );
  XNOR U7333 ( .A(n6607), .B(n6608), .Z(n6609) );
  XNOR U7334 ( .A(n6610), .B(n6609), .Z(n6626) );
  XOR U7335 ( .A(sreg[1242]), .B(n6626), .Z(n6627) );
  XOR U7336 ( .A(n6628), .B(n6627), .Z(c[1242]) );
  NANDN U7337 ( .A(n6608), .B(n6607), .Z(n6612) );
  NAND U7338 ( .A(n6610), .B(n6609), .Z(n6611) );
  NAND U7339 ( .A(n6612), .B(n6611), .Z(n6636) );
  AND U7340 ( .A(b[2]), .B(a[221]), .Z(n6640) );
  AND U7341 ( .A(a[222]), .B(b[1]), .Z(n6638) );
  AND U7342 ( .A(a[220]), .B(b[3]), .Z(n6637) );
  XOR U7343 ( .A(n6638), .B(n6637), .Z(n6639) );
  XOR U7344 ( .A(n6640), .B(n6639), .Z(n6643) );
  NAND U7345 ( .A(b[0]), .B(a[223]), .Z(n6644) );
  XOR U7346 ( .A(n6643), .B(n6644), .Z(n6645) );
  OR U7347 ( .A(n6614), .B(n6613), .Z(n6618) );
  NANDN U7348 ( .A(n6616), .B(n6615), .Z(n6617) );
  AND U7349 ( .A(n6618), .B(n6617), .Z(n6646) );
  XOR U7350 ( .A(n6645), .B(n6646), .Z(n6634) );
  NANDN U7351 ( .A(n6620), .B(n6619), .Z(n6624) );
  OR U7352 ( .A(n6622), .B(n6621), .Z(n6623) );
  AND U7353 ( .A(n6624), .B(n6623), .Z(n6635) );
  XOR U7354 ( .A(n6634), .B(n6635), .Z(n6625) );
  XOR U7355 ( .A(n6636), .B(n6625), .Z(n6633) );
  OR U7356 ( .A(n6626), .B(sreg[1242]), .Z(n6630) );
  NANDN U7357 ( .A(n6628), .B(n6627), .Z(n6629) );
  AND U7358 ( .A(n6630), .B(n6629), .Z(n6632) );
  XOR U7359 ( .A(sreg[1243]), .B(n6632), .Z(n6631) );
  XNOR U7360 ( .A(n6633), .B(n6631), .Z(c[1243]) );
  AND U7361 ( .A(b[2]), .B(a[222]), .Z(n6656) );
  AND U7362 ( .A(a[223]), .B(b[1]), .Z(n6654) );
  AND U7363 ( .A(a[221]), .B(b[3]), .Z(n6653) );
  XOR U7364 ( .A(n6654), .B(n6653), .Z(n6655) );
  XOR U7365 ( .A(n6656), .B(n6655), .Z(n6659) );
  NAND U7366 ( .A(b[0]), .B(a[224]), .Z(n6660) );
  XOR U7367 ( .A(n6659), .B(n6660), .Z(n6662) );
  OR U7368 ( .A(n6638), .B(n6637), .Z(n6642) );
  NANDN U7369 ( .A(n6640), .B(n6639), .Z(n6641) );
  NAND U7370 ( .A(n6642), .B(n6641), .Z(n6661) );
  XNOR U7371 ( .A(n6662), .B(n6661), .Z(n6647) );
  XNOR U7372 ( .A(n6647), .B(n6648), .Z(n6650) );
  XOR U7373 ( .A(n6649), .B(n6650), .Z(n6665) );
  XOR U7374 ( .A(n6665), .B(sreg[1244]), .Z(n6667) );
  XNOR U7375 ( .A(n6666), .B(n6667), .Z(c[1244]) );
  NANDN U7376 ( .A(n6648), .B(n6647), .Z(n6652) );
  NAND U7377 ( .A(n6650), .B(n6649), .Z(n6651) );
  NAND U7378 ( .A(n6652), .B(n6651), .Z(n6676) );
  AND U7379 ( .A(b[2]), .B(a[223]), .Z(n6682) );
  AND U7380 ( .A(a[224]), .B(b[1]), .Z(n6680) );
  AND U7381 ( .A(a[222]), .B(b[3]), .Z(n6679) );
  XOR U7382 ( .A(n6680), .B(n6679), .Z(n6681) );
  XOR U7383 ( .A(n6682), .B(n6681), .Z(n6685) );
  NAND U7384 ( .A(b[0]), .B(a[225]), .Z(n6686) );
  XOR U7385 ( .A(n6685), .B(n6686), .Z(n6688) );
  OR U7386 ( .A(n6654), .B(n6653), .Z(n6658) );
  NANDN U7387 ( .A(n6656), .B(n6655), .Z(n6657) );
  NAND U7388 ( .A(n6658), .B(n6657), .Z(n6687) );
  XNOR U7389 ( .A(n6688), .B(n6687), .Z(n6673) );
  NANDN U7390 ( .A(n6660), .B(n6659), .Z(n6664) );
  OR U7391 ( .A(n6662), .B(n6661), .Z(n6663) );
  NAND U7392 ( .A(n6664), .B(n6663), .Z(n6674) );
  XNOR U7393 ( .A(n6673), .B(n6674), .Z(n6675) );
  XOR U7394 ( .A(n6676), .B(n6675), .Z(n6672) );
  NANDN U7395 ( .A(n6665), .B(sreg[1244]), .Z(n6669) );
  NANDN U7396 ( .A(n6667), .B(n6666), .Z(n6668) );
  NAND U7397 ( .A(n6669), .B(n6668), .Z(n6671) );
  XNOR U7398 ( .A(sreg[1245]), .B(n6671), .Z(n6670) );
  XOR U7399 ( .A(n6672), .B(n6670), .Z(c[1245]) );
  NANDN U7400 ( .A(n6674), .B(n6673), .Z(n6678) );
  NAND U7401 ( .A(n6676), .B(n6675), .Z(n6677) );
  NAND U7402 ( .A(n6678), .B(n6677), .Z(n6694) );
  AND U7403 ( .A(b[2]), .B(a[224]), .Z(n6700) );
  AND U7404 ( .A(a[225]), .B(b[1]), .Z(n6698) );
  AND U7405 ( .A(a[223]), .B(b[3]), .Z(n6697) );
  XOR U7406 ( .A(n6698), .B(n6697), .Z(n6699) );
  XOR U7407 ( .A(n6700), .B(n6699), .Z(n6703) );
  NAND U7408 ( .A(b[0]), .B(a[226]), .Z(n6704) );
  XOR U7409 ( .A(n6703), .B(n6704), .Z(n6706) );
  OR U7410 ( .A(n6680), .B(n6679), .Z(n6684) );
  NANDN U7411 ( .A(n6682), .B(n6681), .Z(n6683) );
  NAND U7412 ( .A(n6684), .B(n6683), .Z(n6705) );
  XNOR U7413 ( .A(n6706), .B(n6705), .Z(n6691) );
  NANDN U7414 ( .A(n6686), .B(n6685), .Z(n6690) );
  OR U7415 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U7416 ( .A(n6690), .B(n6689), .Z(n6692) );
  XNOR U7417 ( .A(n6691), .B(n6692), .Z(n6693) );
  XNOR U7418 ( .A(n6694), .B(n6693), .Z(n6709) );
  XOR U7419 ( .A(sreg[1246]), .B(n6709), .Z(n6711) );
  XNOR U7420 ( .A(n6710), .B(n6711), .Z(c[1246]) );
  NANDN U7421 ( .A(n6692), .B(n6691), .Z(n6696) );
  NAND U7422 ( .A(n6694), .B(n6693), .Z(n6695) );
  NAND U7423 ( .A(n6696), .B(n6695), .Z(n6718) );
  AND U7424 ( .A(b[2]), .B(a[225]), .Z(n6724) );
  AND U7425 ( .A(a[226]), .B(b[1]), .Z(n6722) );
  AND U7426 ( .A(a[224]), .B(b[3]), .Z(n6721) );
  XOR U7427 ( .A(n6722), .B(n6721), .Z(n6723) );
  XOR U7428 ( .A(n6724), .B(n6723), .Z(n6727) );
  NAND U7429 ( .A(b[0]), .B(a[227]), .Z(n6728) );
  XOR U7430 ( .A(n6727), .B(n6728), .Z(n6730) );
  OR U7431 ( .A(n6698), .B(n6697), .Z(n6702) );
  NANDN U7432 ( .A(n6700), .B(n6699), .Z(n6701) );
  NAND U7433 ( .A(n6702), .B(n6701), .Z(n6729) );
  XNOR U7434 ( .A(n6730), .B(n6729), .Z(n6715) );
  NANDN U7435 ( .A(n6704), .B(n6703), .Z(n6708) );
  OR U7436 ( .A(n6706), .B(n6705), .Z(n6707) );
  NAND U7437 ( .A(n6708), .B(n6707), .Z(n6716) );
  XNOR U7438 ( .A(n6715), .B(n6716), .Z(n6717) );
  XOR U7439 ( .A(n6718), .B(n6717), .Z(n6734) );
  OR U7440 ( .A(n6709), .B(sreg[1246]), .Z(n6713) );
  NAND U7441 ( .A(n6711), .B(n6710), .Z(n6712) );
  AND U7442 ( .A(n6713), .B(n6712), .Z(n6733) );
  XNOR U7443 ( .A(sreg[1247]), .B(n6733), .Z(n6714) );
  XOR U7444 ( .A(n6734), .B(n6714), .Z(c[1247]) );
  NANDN U7445 ( .A(n6716), .B(n6715), .Z(n6720) );
  NAND U7446 ( .A(n6718), .B(n6717), .Z(n6719) );
  NAND U7447 ( .A(n6720), .B(n6719), .Z(n6739) );
  AND U7448 ( .A(b[2]), .B(a[226]), .Z(n6745) );
  AND U7449 ( .A(a[227]), .B(b[1]), .Z(n6743) );
  AND U7450 ( .A(a[225]), .B(b[3]), .Z(n6742) );
  XOR U7451 ( .A(n6743), .B(n6742), .Z(n6744) );
  XOR U7452 ( .A(n6745), .B(n6744), .Z(n6748) );
  NAND U7453 ( .A(b[0]), .B(a[228]), .Z(n6749) );
  XOR U7454 ( .A(n6748), .B(n6749), .Z(n6751) );
  OR U7455 ( .A(n6722), .B(n6721), .Z(n6726) );
  NANDN U7456 ( .A(n6724), .B(n6723), .Z(n6725) );
  NAND U7457 ( .A(n6726), .B(n6725), .Z(n6750) );
  XNOR U7458 ( .A(n6751), .B(n6750), .Z(n6736) );
  NANDN U7459 ( .A(n6728), .B(n6727), .Z(n6732) );
  OR U7460 ( .A(n6730), .B(n6729), .Z(n6731) );
  NAND U7461 ( .A(n6732), .B(n6731), .Z(n6737) );
  XNOR U7462 ( .A(n6736), .B(n6737), .Z(n6738) );
  XOR U7463 ( .A(n6739), .B(n6738), .Z(n6755) );
  XNOR U7464 ( .A(sreg[1248]), .B(n6754), .Z(n6735) );
  XOR U7465 ( .A(n6755), .B(n6735), .Z(c[1248]) );
  NANDN U7466 ( .A(n6737), .B(n6736), .Z(n6741) );
  NAND U7467 ( .A(n6739), .B(n6738), .Z(n6740) );
  NAND U7468 ( .A(n6741), .B(n6740), .Z(n6760) );
  AND U7469 ( .A(b[2]), .B(a[227]), .Z(n6766) );
  AND U7470 ( .A(a[228]), .B(b[1]), .Z(n6764) );
  AND U7471 ( .A(a[226]), .B(b[3]), .Z(n6763) );
  XOR U7472 ( .A(n6764), .B(n6763), .Z(n6765) );
  XOR U7473 ( .A(n6766), .B(n6765), .Z(n6769) );
  NAND U7474 ( .A(b[0]), .B(a[229]), .Z(n6770) );
  XOR U7475 ( .A(n6769), .B(n6770), .Z(n6772) );
  OR U7476 ( .A(n6743), .B(n6742), .Z(n6747) );
  NANDN U7477 ( .A(n6745), .B(n6744), .Z(n6746) );
  NAND U7478 ( .A(n6747), .B(n6746), .Z(n6771) );
  XNOR U7479 ( .A(n6772), .B(n6771), .Z(n6757) );
  NANDN U7480 ( .A(n6749), .B(n6748), .Z(n6753) );
  OR U7481 ( .A(n6751), .B(n6750), .Z(n6752) );
  NAND U7482 ( .A(n6753), .B(n6752), .Z(n6758) );
  XNOR U7483 ( .A(n6757), .B(n6758), .Z(n6759) );
  XNOR U7484 ( .A(n6760), .B(n6759), .Z(n6776) );
  XOR U7485 ( .A(n6775), .B(sreg[1249]), .Z(n6756) );
  XOR U7486 ( .A(n6776), .B(n6756), .Z(c[1249]) );
  NANDN U7487 ( .A(n6758), .B(n6757), .Z(n6762) );
  NAND U7488 ( .A(n6760), .B(n6759), .Z(n6761) );
  NAND U7489 ( .A(n6762), .B(n6761), .Z(n6783) );
  AND U7490 ( .A(b[2]), .B(a[228]), .Z(n6789) );
  AND U7491 ( .A(a[229]), .B(b[1]), .Z(n6787) );
  AND U7492 ( .A(a[227]), .B(b[3]), .Z(n6786) );
  XOR U7493 ( .A(n6787), .B(n6786), .Z(n6788) );
  XOR U7494 ( .A(n6789), .B(n6788), .Z(n6792) );
  NAND U7495 ( .A(b[0]), .B(a[230]), .Z(n6793) );
  XOR U7496 ( .A(n6792), .B(n6793), .Z(n6795) );
  OR U7497 ( .A(n6764), .B(n6763), .Z(n6768) );
  NANDN U7498 ( .A(n6766), .B(n6765), .Z(n6767) );
  NAND U7499 ( .A(n6768), .B(n6767), .Z(n6794) );
  XNOR U7500 ( .A(n6795), .B(n6794), .Z(n6780) );
  NANDN U7501 ( .A(n6770), .B(n6769), .Z(n6774) );
  OR U7502 ( .A(n6772), .B(n6771), .Z(n6773) );
  NAND U7503 ( .A(n6774), .B(n6773), .Z(n6781) );
  XNOR U7504 ( .A(n6780), .B(n6781), .Z(n6782) );
  XOR U7505 ( .A(n6783), .B(n6782), .Z(n6779) );
  XOR U7506 ( .A(sreg[1250]), .B(n6778), .Z(n6777) );
  XOR U7507 ( .A(n6779), .B(n6777), .Z(c[1250]) );
  NANDN U7508 ( .A(n6781), .B(n6780), .Z(n6785) );
  NAND U7509 ( .A(n6783), .B(n6782), .Z(n6784) );
  NAND U7510 ( .A(n6785), .B(n6784), .Z(n6801) );
  AND U7511 ( .A(b[2]), .B(a[229]), .Z(n6807) );
  AND U7512 ( .A(a[230]), .B(b[1]), .Z(n6805) );
  AND U7513 ( .A(a[228]), .B(b[3]), .Z(n6804) );
  XOR U7514 ( .A(n6805), .B(n6804), .Z(n6806) );
  XOR U7515 ( .A(n6807), .B(n6806), .Z(n6810) );
  NAND U7516 ( .A(b[0]), .B(a[231]), .Z(n6811) );
  XOR U7517 ( .A(n6810), .B(n6811), .Z(n6813) );
  OR U7518 ( .A(n6787), .B(n6786), .Z(n6791) );
  NANDN U7519 ( .A(n6789), .B(n6788), .Z(n6790) );
  NAND U7520 ( .A(n6791), .B(n6790), .Z(n6812) );
  XNOR U7521 ( .A(n6813), .B(n6812), .Z(n6798) );
  NANDN U7522 ( .A(n6793), .B(n6792), .Z(n6797) );
  OR U7523 ( .A(n6795), .B(n6794), .Z(n6796) );
  NAND U7524 ( .A(n6797), .B(n6796), .Z(n6799) );
  XNOR U7525 ( .A(n6798), .B(n6799), .Z(n6800) );
  XNOR U7526 ( .A(n6801), .B(n6800), .Z(n6816) );
  XNOR U7527 ( .A(n6816), .B(sreg[1251]), .Z(n6817) );
  XOR U7528 ( .A(n6818), .B(n6817), .Z(c[1251]) );
  NANDN U7529 ( .A(n6799), .B(n6798), .Z(n6803) );
  NAND U7530 ( .A(n6801), .B(n6800), .Z(n6802) );
  NAND U7531 ( .A(n6803), .B(n6802), .Z(n6827) );
  AND U7532 ( .A(b[2]), .B(a[230]), .Z(n6833) );
  AND U7533 ( .A(a[231]), .B(b[1]), .Z(n6831) );
  AND U7534 ( .A(a[229]), .B(b[3]), .Z(n6830) );
  XOR U7535 ( .A(n6831), .B(n6830), .Z(n6832) );
  XOR U7536 ( .A(n6833), .B(n6832), .Z(n6836) );
  NAND U7537 ( .A(b[0]), .B(a[232]), .Z(n6837) );
  XOR U7538 ( .A(n6836), .B(n6837), .Z(n6839) );
  OR U7539 ( .A(n6805), .B(n6804), .Z(n6809) );
  NANDN U7540 ( .A(n6807), .B(n6806), .Z(n6808) );
  NAND U7541 ( .A(n6809), .B(n6808), .Z(n6838) );
  XNOR U7542 ( .A(n6839), .B(n6838), .Z(n6824) );
  NANDN U7543 ( .A(n6811), .B(n6810), .Z(n6815) );
  OR U7544 ( .A(n6813), .B(n6812), .Z(n6814) );
  NAND U7545 ( .A(n6815), .B(n6814), .Z(n6825) );
  XNOR U7546 ( .A(n6824), .B(n6825), .Z(n6826) );
  XOR U7547 ( .A(n6827), .B(n6826), .Z(n6823) );
  NAND U7548 ( .A(n6816), .B(sreg[1251]), .Z(n6820) );
  OR U7549 ( .A(n6818), .B(n6817), .Z(n6819) );
  NAND U7550 ( .A(n6820), .B(n6819), .Z(n6822) );
  XNOR U7551 ( .A(sreg[1252]), .B(n6822), .Z(n6821) );
  XOR U7552 ( .A(n6823), .B(n6821), .Z(c[1252]) );
  NANDN U7553 ( .A(n6825), .B(n6824), .Z(n6829) );
  NAND U7554 ( .A(n6827), .B(n6826), .Z(n6828) );
  NAND U7555 ( .A(n6829), .B(n6828), .Z(n6845) );
  AND U7556 ( .A(b[2]), .B(a[231]), .Z(n6851) );
  AND U7557 ( .A(a[232]), .B(b[1]), .Z(n6849) );
  AND U7558 ( .A(a[230]), .B(b[3]), .Z(n6848) );
  XOR U7559 ( .A(n6849), .B(n6848), .Z(n6850) );
  XOR U7560 ( .A(n6851), .B(n6850), .Z(n6854) );
  NAND U7561 ( .A(b[0]), .B(a[233]), .Z(n6855) );
  XOR U7562 ( .A(n6854), .B(n6855), .Z(n6857) );
  OR U7563 ( .A(n6831), .B(n6830), .Z(n6835) );
  NANDN U7564 ( .A(n6833), .B(n6832), .Z(n6834) );
  NAND U7565 ( .A(n6835), .B(n6834), .Z(n6856) );
  XNOR U7566 ( .A(n6857), .B(n6856), .Z(n6842) );
  NANDN U7567 ( .A(n6837), .B(n6836), .Z(n6841) );
  OR U7568 ( .A(n6839), .B(n6838), .Z(n6840) );
  NAND U7569 ( .A(n6841), .B(n6840), .Z(n6843) );
  XNOR U7570 ( .A(n6842), .B(n6843), .Z(n6844) );
  XNOR U7571 ( .A(n6845), .B(n6844), .Z(n6860) );
  XNOR U7572 ( .A(n6860), .B(sreg[1253]), .Z(n6861) );
  XOR U7573 ( .A(n6862), .B(n6861), .Z(c[1253]) );
  NANDN U7574 ( .A(n6843), .B(n6842), .Z(n6847) );
  NAND U7575 ( .A(n6845), .B(n6844), .Z(n6846) );
  NAND U7576 ( .A(n6847), .B(n6846), .Z(n6868) );
  AND U7577 ( .A(b[2]), .B(a[232]), .Z(n6874) );
  AND U7578 ( .A(a[233]), .B(b[1]), .Z(n6872) );
  AND U7579 ( .A(a[231]), .B(b[3]), .Z(n6871) );
  XOR U7580 ( .A(n6872), .B(n6871), .Z(n6873) );
  XOR U7581 ( .A(n6874), .B(n6873), .Z(n6877) );
  NAND U7582 ( .A(b[0]), .B(a[234]), .Z(n6878) );
  XOR U7583 ( .A(n6877), .B(n6878), .Z(n6880) );
  OR U7584 ( .A(n6849), .B(n6848), .Z(n6853) );
  NANDN U7585 ( .A(n6851), .B(n6850), .Z(n6852) );
  NAND U7586 ( .A(n6853), .B(n6852), .Z(n6879) );
  XNOR U7587 ( .A(n6880), .B(n6879), .Z(n6865) );
  NANDN U7588 ( .A(n6855), .B(n6854), .Z(n6859) );
  OR U7589 ( .A(n6857), .B(n6856), .Z(n6858) );
  NAND U7590 ( .A(n6859), .B(n6858), .Z(n6866) );
  XNOR U7591 ( .A(n6865), .B(n6866), .Z(n6867) );
  XNOR U7592 ( .A(n6868), .B(n6867), .Z(n6883) );
  XOR U7593 ( .A(sreg[1254]), .B(n6883), .Z(n6884) );
  NAND U7594 ( .A(n6860), .B(sreg[1253]), .Z(n6864) );
  OR U7595 ( .A(n6862), .B(n6861), .Z(n6863) );
  NAND U7596 ( .A(n6864), .B(n6863), .Z(n6885) );
  XOR U7597 ( .A(n6884), .B(n6885), .Z(c[1254]) );
  NANDN U7598 ( .A(n6866), .B(n6865), .Z(n6870) );
  NAND U7599 ( .A(n6868), .B(n6867), .Z(n6869) );
  NAND U7600 ( .A(n6870), .B(n6869), .Z(n6891) );
  AND U7601 ( .A(b[2]), .B(a[233]), .Z(n6897) );
  AND U7602 ( .A(a[234]), .B(b[1]), .Z(n6895) );
  AND U7603 ( .A(a[232]), .B(b[3]), .Z(n6894) );
  XOR U7604 ( .A(n6895), .B(n6894), .Z(n6896) );
  XOR U7605 ( .A(n6897), .B(n6896), .Z(n6900) );
  NAND U7606 ( .A(b[0]), .B(a[235]), .Z(n6901) );
  XOR U7607 ( .A(n6900), .B(n6901), .Z(n6903) );
  OR U7608 ( .A(n6872), .B(n6871), .Z(n6876) );
  NANDN U7609 ( .A(n6874), .B(n6873), .Z(n6875) );
  NAND U7610 ( .A(n6876), .B(n6875), .Z(n6902) );
  XNOR U7611 ( .A(n6903), .B(n6902), .Z(n6888) );
  NANDN U7612 ( .A(n6878), .B(n6877), .Z(n6882) );
  OR U7613 ( .A(n6880), .B(n6879), .Z(n6881) );
  NAND U7614 ( .A(n6882), .B(n6881), .Z(n6889) );
  XNOR U7615 ( .A(n6888), .B(n6889), .Z(n6890) );
  XNOR U7616 ( .A(n6891), .B(n6890), .Z(n6906) );
  XNOR U7617 ( .A(n6906), .B(sreg[1255]), .Z(n6908) );
  OR U7618 ( .A(n6883), .B(sreg[1254]), .Z(n6887) );
  NANDN U7619 ( .A(n6885), .B(n6884), .Z(n6886) );
  NAND U7620 ( .A(n6887), .B(n6886), .Z(n6907) );
  XOR U7621 ( .A(n6908), .B(n6907), .Z(c[1255]) );
  NANDN U7622 ( .A(n6889), .B(n6888), .Z(n6893) );
  NAND U7623 ( .A(n6891), .B(n6890), .Z(n6892) );
  NAND U7624 ( .A(n6893), .B(n6892), .Z(n6914) );
  AND U7625 ( .A(b[2]), .B(a[234]), .Z(n6920) );
  AND U7626 ( .A(a[235]), .B(b[1]), .Z(n6918) );
  AND U7627 ( .A(a[233]), .B(b[3]), .Z(n6917) );
  XOR U7628 ( .A(n6918), .B(n6917), .Z(n6919) );
  XOR U7629 ( .A(n6920), .B(n6919), .Z(n6923) );
  NAND U7630 ( .A(b[0]), .B(a[236]), .Z(n6924) );
  XOR U7631 ( .A(n6923), .B(n6924), .Z(n6926) );
  OR U7632 ( .A(n6895), .B(n6894), .Z(n6899) );
  NANDN U7633 ( .A(n6897), .B(n6896), .Z(n6898) );
  NAND U7634 ( .A(n6899), .B(n6898), .Z(n6925) );
  XNOR U7635 ( .A(n6926), .B(n6925), .Z(n6911) );
  NANDN U7636 ( .A(n6901), .B(n6900), .Z(n6905) );
  OR U7637 ( .A(n6903), .B(n6902), .Z(n6904) );
  NAND U7638 ( .A(n6905), .B(n6904), .Z(n6912) );
  XNOR U7639 ( .A(n6911), .B(n6912), .Z(n6913) );
  XNOR U7640 ( .A(n6914), .B(n6913), .Z(n6929) );
  XNOR U7641 ( .A(n6929), .B(sreg[1256]), .Z(n6931) );
  NAND U7642 ( .A(n6906), .B(sreg[1255]), .Z(n6910) );
  OR U7643 ( .A(n6908), .B(n6907), .Z(n6909) );
  AND U7644 ( .A(n6910), .B(n6909), .Z(n6930) );
  XOR U7645 ( .A(n6931), .B(n6930), .Z(c[1256]) );
  NANDN U7646 ( .A(n6912), .B(n6911), .Z(n6916) );
  NAND U7647 ( .A(n6914), .B(n6913), .Z(n6915) );
  NAND U7648 ( .A(n6916), .B(n6915), .Z(n6942) );
  AND U7649 ( .A(b[2]), .B(a[235]), .Z(n6948) );
  AND U7650 ( .A(a[236]), .B(b[1]), .Z(n6946) );
  AND U7651 ( .A(a[234]), .B(b[3]), .Z(n6945) );
  XOR U7652 ( .A(n6946), .B(n6945), .Z(n6947) );
  XOR U7653 ( .A(n6948), .B(n6947), .Z(n6951) );
  NAND U7654 ( .A(b[0]), .B(a[237]), .Z(n6952) );
  XOR U7655 ( .A(n6951), .B(n6952), .Z(n6954) );
  OR U7656 ( .A(n6918), .B(n6917), .Z(n6922) );
  NANDN U7657 ( .A(n6920), .B(n6919), .Z(n6921) );
  NAND U7658 ( .A(n6922), .B(n6921), .Z(n6953) );
  XNOR U7659 ( .A(n6954), .B(n6953), .Z(n6939) );
  NANDN U7660 ( .A(n6924), .B(n6923), .Z(n6928) );
  OR U7661 ( .A(n6926), .B(n6925), .Z(n6927) );
  NAND U7662 ( .A(n6928), .B(n6927), .Z(n6940) );
  XNOR U7663 ( .A(n6939), .B(n6940), .Z(n6941) );
  XNOR U7664 ( .A(n6942), .B(n6941), .Z(n6934) );
  XOR U7665 ( .A(sreg[1257]), .B(n6934), .Z(n6935) );
  NAND U7666 ( .A(n6929), .B(sreg[1256]), .Z(n6933) );
  OR U7667 ( .A(n6931), .B(n6930), .Z(n6932) );
  NAND U7668 ( .A(n6933), .B(n6932), .Z(n6936) );
  XOR U7669 ( .A(n6935), .B(n6936), .Z(c[1257]) );
  OR U7670 ( .A(n6934), .B(sreg[1257]), .Z(n6938) );
  NANDN U7671 ( .A(n6936), .B(n6935), .Z(n6937) );
  AND U7672 ( .A(n6938), .B(n6937), .Z(n6976) );
  NANDN U7673 ( .A(n6940), .B(n6939), .Z(n6944) );
  NAND U7674 ( .A(n6942), .B(n6941), .Z(n6943) );
  NAND U7675 ( .A(n6944), .B(n6943), .Z(n6961) );
  AND U7676 ( .A(b[2]), .B(a[236]), .Z(n6967) );
  AND U7677 ( .A(a[237]), .B(b[1]), .Z(n6965) );
  AND U7678 ( .A(a[235]), .B(b[3]), .Z(n6964) );
  XOR U7679 ( .A(n6965), .B(n6964), .Z(n6966) );
  XOR U7680 ( .A(n6967), .B(n6966), .Z(n6970) );
  NAND U7681 ( .A(b[0]), .B(a[238]), .Z(n6971) );
  XOR U7682 ( .A(n6970), .B(n6971), .Z(n6973) );
  OR U7683 ( .A(n6946), .B(n6945), .Z(n6950) );
  NANDN U7684 ( .A(n6948), .B(n6947), .Z(n6949) );
  NAND U7685 ( .A(n6950), .B(n6949), .Z(n6972) );
  XNOR U7686 ( .A(n6973), .B(n6972), .Z(n6958) );
  NANDN U7687 ( .A(n6952), .B(n6951), .Z(n6956) );
  OR U7688 ( .A(n6954), .B(n6953), .Z(n6955) );
  NAND U7689 ( .A(n6956), .B(n6955), .Z(n6959) );
  XNOR U7690 ( .A(n6958), .B(n6959), .Z(n6960) );
  XNOR U7691 ( .A(n6961), .B(n6960), .Z(n6977) );
  XOR U7692 ( .A(sreg[1258]), .B(n6977), .Z(n6957) );
  XOR U7693 ( .A(n6976), .B(n6957), .Z(c[1258]) );
  NANDN U7694 ( .A(n6959), .B(n6958), .Z(n6963) );
  NAND U7695 ( .A(n6961), .B(n6960), .Z(n6962) );
  NAND U7696 ( .A(n6963), .B(n6962), .Z(n6984) );
  AND U7697 ( .A(b[2]), .B(a[237]), .Z(n6990) );
  AND U7698 ( .A(a[238]), .B(b[1]), .Z(n6988) );
  AND U7699 ( .A(a[236]), .B(b[3]), .Z(n6987) );
  XOR U7700 ( .A(n6988), .B(n6987), .Z(n6989) );
  XOR U7701 ( .A(n6990), .B(n6989), .Z(n6993) );
  NAND U7702 ( .A(b[0]), .B(a[239]), .Z(n6994) );
  XOR U7703 ( .A(n6993), .B(n6994), .Z(n6996) );
  OR U7704 ( .A(n6965), .B(n6964), .Z(n6969) );
  NANDN U7705 ( .A(n6967), .B(n6966), .Z(n6968) );
  NAND U7706 ( .A(n6969), .B(n6968), .Z(n6995) );
  XNOR U7707 ( .A(n6996), .B(n6995), .Z(n6981) );
  NANDN U7708 ( .A(n6971), .B(n6970), .Z(n6975) );
  OR U7709 ( .A(n6973), .B(n6972), .Z(n6974) );
  NAND U7710 ( .A(n6975), .B(n6974), .Z(n6982) );
  XNOR U7711 ( .A(n6981), .B(n6982), .Z(n6983) );
  XNOR U7712 ( .A(n6984), .B(n6983), .Z(n6980) );
  XOR U7713 ( .A(n6979), .B(sreg[1259]), .Z(n6978) );
  XOR U7714 ( .A(n6980), .B(n6978), .Z(c[1259]) );
  NANDN U7715 ( .A(n6982), .B(n6981), .Z(n6986) );
  NAND U7716 ( .A(n6984), .B(n6983), .Z(n6985) );
  NAND U7717 ( .A(n6986), .B(n6985), .Z(n7002) );
  AND U7718 ( .A(b[2]), .B(a[238]), .Z(n7014) );
  AND U7719 ( .A(a[239]), .B(b[1]), .Z(n7012) );
  AND U7720 ( .A(a[237]), .B(b[3]), .Z(n7011) );
  XOR U7721 ( .A(n7012), .B(n7011), .Z(n7013) );
  XOR U7722 ( .A(n7014), .B(n7013), .Z(n7005) );
  NAND U7723 ( .A(b[0]), .B(a[240]), .Z(n7006) );
  XOR U7724 ( .A(n7005), .B(n7006), .Z(n7008) );
  OR U7725 ( .A(n6988), .B(n6987), .Z(n6992) );
  NANDN U7726 ( .A(n6990), .B(n6989), .Z(n6991) );
  NAND U7727 ( .A(n6992), .B(n6991), .Z(n7007) );
  XNOR U7728 ( .A(n7008), .B(n7007), .Z(n6999) );
  NANDN U7729 ( .A(n6994), .B(n6993), .Z(n6998) );
  OR U7730 ( .A(n6996), .B(n6995), .Z(n6997) );
  NAND U7731 ( .A(n6998), .B(n6997), .Z(n7000) );
  XNOR U7732 ( .A(n6999), .B(n7000), .Z(n7001) );
  XNOR U7733 ( .A(n7002), .B(n7001), .Z(n7018) );
  XNOR U7734 ( .A(n7018), .B(sreg[1260]), .Z(n7020) );
  XNOR U7735 ( .A(n7019), .B(n7020), .Z(c[1260]) );
  NANDN U7736 ( .A(n7000), .B(n6999), .Z(n7004) );
  NAND U7737 ( .A(n7002), .B(n7001), .Z(n7003) );
  NAND U7738 ( .A(n7004), .B(n7003), .Z(n7025) );
  NANDN U7739 ( .A(n7006), .B(n7005), .Z(n7010) );
  OR U7740 ( .A(n7008), .B(n7007), .Z(n7009) );
  AND U7741 ( .A(n7010), .B(n7009), .Z(n7024) );
  AND U7742 ( .A(b[2]), .B(a[239]), .Z(n7029) );
  AND U7743 ( .A(a[240]), .B(b[1]), .Z(n7027) );
  AND U7744 ( .A(a[238]), .B(b[3]), .Z(n7026) );
  XOR U7745 ( .A(n7027), .B(n7026), .Z(n7028) );
  XOR U7746 ( .A(n7029), .B(n7028), .Z(n7032) );
  NAND U7747 ( .A(b[0]), .B(a[241]), .Z(n7033) );
  XOR U7748 ( .A(n7032), .B(n7033), .Z(n7035) );
  OR U7749 ( .A(n7012), .B(n7011), .Z(n7016) );
  NANDN U7750 ( .A(n7014), .B(n7013), .Z(n7015) );
  NAND U7751 ( .A(n7016), .B(n7015), .Z(n7034) );
  XOR U7752 ( .A(n7035), .B(n7034), .Z(n7023) );
  XNOR U7753 ( .A(n7024), .B(n7023), .Z(n7017) );
  XNOR U7754 ( .A(n7025), .B(n7017), .Z(n7038) );
  XOR U7755 ( .A(sreg[1261]), .B(n7038), .Z(n7039) );
  NAND U7756 ( .A(n7018), .B(sreg[1260]), .Z(n7022) );
  NANDN U7757 ( .A(n7020), .B(n7019), .Z(n7021) );
  NAND U7758 ( .A(n7022), .B(n7021), .Z(n7040) );
  XOR U7759 ( .A(n7039), .B(n7040), .Z(c[1261]) );
  AND U7760 ( .A(b[2]), .B(a[240]), .Z(n7055) );
  AND U7761 ( .A(a[241]), .B(b[1]), .Z(n7053) );
  AND U7762 ( .A(a[239]), .B(b[3]), .Z(n7052) );
  XOR U7763 ( .A(n7053), .B(n7052), .Z(n7054) );
  XOR U7764 ( .A(n7055), .B(n7054), .Z(n7058) );
  NAND U7765 ( .A(b[0]), .B(a[242]), .Z(n7059) );
  XOR U7766 ( .A(n7058), .B(n7059), .Z(n7061) );
  OR U7767 ( .A(n7027), .B(n7026), .Z(n7031) );
  NANDN U7768 ( .A(n7029), .B(n7028), .Z(n7030) );
  NAND U7769 ( .A(n7031), .B(n7030), .Z(n7060) );
  XNOR U7770 ( .A(n7061), .B(n7060), .Z(n7046) );
  NANDN U7771 ( .A(n7033), .B(n7032), .Z(n7037) );
  OR U7772 ( .A(n7035), .B(n7034), .Z(n7036) );
  NAND U7773 ( .A(n7037), .B(n7036), .Z(n7047) );
  XNOR U7774 ( .A(n7046), .B(n7047), .Z(n7048) );
  XOR U7775 ( .A(n7049), .B(n7048), .Z(n7045) );
  OR U7776 ( .A(n7038), .B(sreg[1261]), .Z(n7042) );
  NANDN U7777 ( .A(n7040), .B(n7039), .Z(n7041) );
  AND U7778 ( .A(n7042), .B(n7041), .Z(n7044) );
  XNOR U7779 ( .A(sreg[1262]), .B(n7044), .Z(n7043) );
  XNOR U7780 ( .A(n7045), .B(n7043), .Z(c[1262]) );
  NANDN U7781 ( .A(n7047), .B(n7046), .Z(n7051) );
  NANDN U7782 ( .A(n7049), .B(n7048), .Z(n7050) );
  NAND U7783 ( .A(n7051), .B(n7050), .Z(n7072) );
  AND U7784 ( .A(b[2]), .B(a[241]), .Z(n7078) );
  AND U7785 ( .A(a[242]), .B(b[1]), .Z(n7076) );
  AND U7786 ( .A(a[240]), .B(b[3]), .Z(n7075) );
  XOR U7787 ( .A(n7076), .B(n7075), .Z(n7077) );
  XOR U7788 ( .A(n7078), .B(n7077), .Z(n7081) );
  NAND U7789 ( .A(b[0]), .B(a[243]), .Z(n7082) );
  XOR U7790 ( .A(n7081), .B(n7082), .Z(n7084) );
  OR U7791 ( .A(n7053), .B(n7052), .Z(n7057) );
  NANDN U7792 ( .A(n7055), .B(n7054), .Z(n7056) );
  NAND U7793 ( .A(n7057), .B(n7056), .Z(n7083) );
  XNOR U7794 ( .A(n7084), .B(n7083), .Z(n7069) );
  NANDN U7795 ( .A(n7059), .B(n7058), .Z(n7063) );
  OR U7796 ( .A(n7061), .B(n7060), .Z(n7062) );
  NAND U7797 ( .A(n7063), .B(n7062), .Z(n7070) );
  XNOR U7798 ( .A(n7069), .B(n7070), .Z(n7071) );
  XNOR U7799 ( .A(n7072), .B(n7071), .Z(n7064) );
  XNOR U7800 ( .A(n7064), .B(sreg[1263]), .Z(n7065) );
  XOR U7801 ( .A(n7066), .B(n7065), .Z(c[1263]) );
  NAND U7802 ( .A(n7064), .B(sreg[1263]), .Z(n7068) );
  OR U7803 ( .A(n7066), .B(n7065), .Z(n7067) );
  NAND U7804 ( .A(n7068), .B(n7067), .Z(n7102) );
  NANDN U7805 ( .A(n7070), .B(n7069), .Z(n7074) );
  NAND U7806 ( .A(n7072), .B(n7071), .Z(n7073) );
  AND U7807 ( .A(n7074), .B(n7073), .Z(n7091) );
  AND U7808 ( .A(b[2]), .B(a[242]), .Z(n7099) );
  AND U7809 ( .A(a[243]), .B(b[1]), .Z(n7097) );
  AND U7810 ( .A(a[241]), .B(b[3]), .Z(n7096) );
  XOR U7811 ( .A(n7097), .B(n7096), .Z(n7098) );
  XOR U7812 ( .A(n7099), .B(n7098), .Z(n7092) );
  NAND U7813 ( .A(b[0]), .B(a[244]), .Z(n7093) );
  XOR U7814 ( .A(n7092), .B(n7093), .Z(n7094) );
  OR U7815 ( .A(n7076), .B(n7075), .Z(n7080) );
  NANDN U7816 ( .A(n7078), .B(n7077), .Z(n7079) );
  AND U7817 ( .A(n7080), .B(n7079), .Z(n7095) );
  XOR U7818 ( .A(n7094), .B(n7095), .Z(n7089) );
  NANDN U7819 ( .A(n7082), .B(n7081), .Z(n7086) );
  OR U7820 ( .A(n7084), .B(n7083), .Z(n7085) );
  AND U7821 ( .A(n7086), .B(n7085), .Z(n7090) );
  XOR U7822 ( .A(n7089), .B(n7090), .Z(n7087) );
  XNOR U7823 ( .A(n7091), .B(n7087), .Z(n7103) );
  XOR U7824 ( .A(sreg[1264]), .B(n7103), .Z(n7088) );
  XNOR U7825 ( .A(n7102), .B(n7088), .Z(c[1264]) );
  AND U7826 ( .A(b[2]), .B(a[243]), .Z(n7108) );
  AND U7827 ( .A(a[244]), .B(b[1]), .Z(n7106) );
  AND U7828 ( .A(a[242]), .B(b[3]), .Z(n7105) );
  XOR U7829 ( .A(n7106), .B(n7105), .Z(n7107) );
  XOR U7830 ( .A(n7108), .B(n7107), .Z(n7111) );
  NAND U7831 ( .A(b[0]), .B(a[245]), .Z(n7112) );
  XNOR U7832 ( .A(n7111), .B(n7112), .Z(n7113) );
  OR U7833 ( .A(n7097), .B(n7096), .Z(n7101) );
  NANDN U7834 ( .A(n7099), .B(n7098), .Z(n7100) );
  AND U7835 ( .A(n7101), .B(n7100), .Z(n7114) );
  XNOR U7836 ( .A(n7113), .B(n7114), .Z(n7118) );
  XNOR U7837 ( .A(n7117), .B(n7118), .Z(n7119) );
  XNOR U7838 ( .A(n7120), .B(n7119), .Z(n7123) );
  XNOR U7839 ( .A(sreg[1265]), .B(n7124), .Z(n7104) );
  XOR U7840 ( .A(n7123), .B(n7104), .Z(c[1265]) );
  AND U7841 ( .A(b[2]), .B(a[244]), .Z(n7135) );
  AND U7842 ( .A(a[245]), .B(b[1]), .Z(n7133) );
  AND U7843 ( .A(a[243]), .B(b[3]), .Z(n7132) );
  XOR U7844 ( .A(n7133), .B(n7132), .Z(n7134) );
  XOR U7845 ( .A(n7135), .B(n7134), .Z(n7138) );
  NAND U7846 ( .A(b[0]), .B(a[246]), .Z(n7139) );
  XOR U7847 ( .A(n7138), .B(n7139), .Z(n7141) );
  OR U7848 ( .A(n7106), .B(n7105), .Z(n7110) );
  NANDN U7849 ( .A(n7108), .B(n7107), .Z(n7109) );
  NAND U7850 ( .A(n7110), .B(n7109), .Z(n7140) );
  XNOR U7851 ( .A(n7141), .B(n7140), .Z(n7126) );
  NANDN U7852 ( .A(n7112), .B(n7111), .Z(n7116) );
  NAND U7853 ( .A(n7114), .B(n7113), .Z(n7115) );
  NAND U7854 ( .A(n7116), .B(n7115), .Z(n7127) );
  XNOR U7855 ( .A(n7126), .B(n7127), .Z(n7128) );
  NANDN U7856 ( .A(n7118), .B(n7117), .Z(n7122) );
  NANDN U7857 ( .A(n7120), .B(n7119), .Z(n7121) );
  NAND U7858 ( .A(n7122), .B(n7121), .Z(n7129) );
  XOR U7859 ( .A(n7128), .B(n7129), .Z(n7145) );
  XOR U7860 ( .A(sreg[1266]), .B(n7144), .Z(n7125) );
  XNOR U7861 ( .A(n7145), .B(n7125), .Z(c[1266]) );
  NANDN U7862 ( .A(n7127), .B(n7126), .Z(n7131) );
  NANDN U7863 ( .A(n7129), .B(n7128), .Z(n7130) );
  NAND U7864 ( .A(n7131), .B(n7130), .Z(n7162) );
  AND U7865 ( .A(b[2]), .B(a[245]), .Z(n7156) );
  AND U7866 ( .A(a[246]), .B(b[1]), .Z(n7154) );
  AND U7867 ( .A(a[244]), .B(b[3]), .Z(n7153) );
  XOR U7868 ( .A(n7154), .B(n7153), .Z(n7155) );
  XOR U7869 ( .A(n7156), .B(n7155), .Z(n7147) );
  NAND U7870 ( .A(b[0]), .B(a[247]), .Z(n7148) );
  XOR U7871 ( .A(n7147), .B(n7148), .Z(n7150) );
  OR U7872 ( .A(n7133), .B(n7132), .Z(n7137) );
  NANDN U7873 ( .A(n7135), .B(n7134), .Z(n7136) );
  NAND U7874 ( .A(n7137), .B(n7136), .Z(n7149) );
  XNOR U7875 ( .A(n7150), .B(n7149), .Z(n7159) );
  NANDN U7876 ( .A(n7139), .B(n7138), .Z(n7143) );
  OR U7877 ( .A(n7141), .B(n7140), .Z(n7142) );
  NAND U7878 ( .A(n7143), .B(n7142), .Z(n7160) );
  XNOR U7879 ( .A(n7159), .B(n7160), .Z(n7161) );
  XOR U7880 ( .A(n7162), .B(n7161), .Z(n7166) );
  XNOR U7881 ( .A(sreg[1267]), .B(n7165), .Z(n7146) );
  XOR U7882 ( .A(n7166), .B(n7146), .Z(c[1267]) );
  NANDN U7883 ( .A(n7148), .B(n7147), .Z(n7152) );
  OR U7884 ( .A(n7150), .B(n7149), .Z(n7151) );
  NAND U7885 ( .A(n7152), .B(n7151), .Z(n7180) );
  AND U7886 ( .A(b[2]), .B(a[246]), .Z(n7171) );
  AND U7887 ( .A(a[247]), .B(b[1]), .Z(n7169) );
  AND U7888 ( .A(a[245]), .B(b[3]), .Z(n7168) );
  XOR U7889 ( .A(n7169), .B(n7168), .Z(n7170) );
  XOR U7890 ( .A(n7171), .B(n7170), .Z(n7174) );
  NAND U7891 ( .A(b[0]), .B(a[248]), .Z(n7175) );
  XNOR U7892 ( .A(n7174), .B(n7175), .Z(n7176) );
  OR U7893 ( .A(n7154), .B(n7153), .Z(n7158) );
  NANDN U7894 ( .A(n7156), .B(n7155), .Z(n7157) );
  AND U7895 ( .A(n7158), .B(n7157), .Z(n7177) );
  XNOR U7896 ( .A(n7176), .B(n7177), .Z(n7181) );
  XNOR U7897 ( .A(n7180), .B(n7181), .Z(n7182) );
  NANDN U7898 ( .A(n7160), .B(n7159), .Z(n7164) );
  NAND U7899 ( .A(n7162), .B(n7161), .Z(n7163) );
  AND U7900 ( .A(n7164), .B(n7163), .Z(n7183) );
  XNOR U7901 ( .A(n7182), .B(n7183), .Z(n7187) );
  XNOR U7902 ( .A(sreg[1268]), .B(n7186), .Z(n7167) );
  XOR U7903 ( .A(n7187), .B(n7167), .Z(c[1268]) );
  AND U7904 ( .A(b[2]), .B(a[247]), .Z(n7200) );
  AND U7905 ( .A(a[248]), .B(b[1]), .Z(n7198) );
  AND U7906 ( .A(a[246]), .B(b[3]), .Z(n7197) );
  XOR U7907 ( .A(n7198), .B(n7197), .Z(n7199) );
  XOR U7908 ( .A(n7200), .B(n7199), .Z(n7203) );
  NAND U7909 ( .A(b[0]), .B(a[249]), .Z(n7204) );
  XOR U7910 ( .A(n7203), .B(n7204), .Z(n7206) );
  OR U7911 ( .A(n7169), .B(n7168), .Z(n7173) );
  NANDN U7912 ( .A(n7171), .B(n7170), .Z(n7172) );
  NAND U7913 ( .A(n7173), .B(n7172), .Z(n7205) );
  XNOR U7914 ( .A(n7206), .B(n7205), .Z(n7191) );
  NANDN U7915 ( .A(n7175), .B(n7174), .Z(n7179) );
  NAND U7916 ( .A(n7177), .B(n7176), .Z(n7178) );
  NAND U7917 ( .A(n7179), .B(n7178), .Z(n7192) );
  XNOR U7918 ( .A(n7191), .B(n7192), .Z(n7193) );
  NANDN U7919 ( .A(n7181), .B(n7180), .Z(n7185) );
  NAND U7920 ( .A(n7183), .B(n7182), .Z(n7184) );
  AND U7921 ( .A(n7185), .B(n7184), .Z(n7194) );
  XNOR U7922 ( .A(n7193), .B(n7194), .Z(n7190) );
  XOR U7923 ( .A(n7189), .B(sreg[1269]), .Z(n7188) );
  XOR U7924 ( .A(n7190), .B(n7188), .Z(c[1269]) );
  NANDN U7925 ( .A(n7192), .B(n7191), .Z(n7196) );
  NAND U7926 ( .A(n7194), .B(n7193), .Z(n7195) );
  NAND U7927 ( .A(n7196), .B(n7195), .Z(n7212) );
  AND U7928 ( .A(b[2]), .B(a[248]), .Z(n7218) );
  AND U7929 ( .A(a[249]), .B(b[1]), .Z(n7216) );
  AND U7930 ( .A(a[247]), .B(b[3]), .Z(n7215) );
  XOR U7931 ( .A(n7216), .B(n7215), .Z(n7217) );
  XOR U7932 ( .A(n7218), .B(n7217), .Z(n7221) );
  NAND U7933 ( .A(b[0]), .B(a[250]), .Z(n7222) );
  XOR U7934 ( .A(n7221), .B(n7222), .Z(n7224) );
  OR U7935 ( .A(n7198), .B(n7197), .Z(n7202) );
  NANDN U7936 ( .A(n7200), .B(n7199), .Z(n7201) );
  NAND U7937 ( .A(n7202), .B(n7201), .Z(n7223) );
  XNOR U7938 ( .A(n7224), .B(n7223), .Z(n7209) );
  NANDN U7939 ( .A(n7204), .B(n7203), .Z(n7208) );
  OR U7940 ( .A(n7206), .B(n7205), .Z(n7207) );
  NAND U7941 ( .A(n7208), .B(n7207), .Z(n7210) );
  XNOR U7942 ( .A(n7209), .B(n7210), .Z(n7211) );
  XNOR U7943 ( .A(n7212), .B(n7211), .Z(n7227) );
  XNOR U7944 ( .A(n7227), .B(sreg[1270]), .Z(n7229) );
  XNOR U7945 ( .A(n7228), .B(n7229), .Z(c[1270]) );
  NANDN U7946 ( .A(n7210), .B(n7209), .Z(n7214) );
  NAND U7947 ( .A(n7212), .B(n7211), .Z(n7213) );
  NAND U7948 ( .A(n7214), .B(n7213), .Z(n7238) );
  AND U7949 ( .A(b[2]), .B(a[249]), .Z(n7244) );
  AND U7950 ( .A(a[250]), .B(b[1]), .Z(n7242) );
  AND U7951 ( .A(a[248]), .B(b[3]), .Z(n7241) );
  XOR U7952 ( .A(n7242), .B(n7241), .Z(n7243) );
  XOR U7953 ( .A(n7244), .B(n7243), .Z(n7247) );
  NAND U7954 ( .A(b[0]), .B(a[251]), .Z(n7248) );
  XOR U7955 ( .A(n7247), .B(n7248), .Z(n7250) );
  OR U7956 ( .A(n7216), .B(n7215), .Z(n7220) );
  NANDN U7957 ( .A(n7218), .B(n7217), .Z(n7219) );
  NAND U7958 ( .A(n7220), .B(n7219), .Z(n7249) );
  XNOR U7959 ( .A(n7250), .B(n7249), .Z(n7235) );
  NANDN U7960 ( .A(n7222), .B(n7221), .Z(n7226) );
  OR U7961 ( .A(n7224), .B(n7223), .Z(n7225) );
  NAND U7962 ( .A(n7226), .B(n7225), .Z(n7236) );
  XNOR U7963 ( .A(n7235), .B(n7236), .Z(n7237) );
  XNOR U7964 ( .A(n7238), .B(n7237), .Z(n7234) );
  NAND U7965 ( .A(n7227), .B(sreg[1270]), .Z(n7231) );
  NANDN U7966 ( .A(n7229), .B(n7228), .Z(n7230) );
  AND U7967 ( .A(n7231), .B(n7230), .Z(n7233) );
  XNOR U7968 ( .A(n7233), .B(sreg[1271]), .Z(n7232) );
  XOR U7969 ( .A(n7234), .B(n7232), .Z(c[1271]) );
  NANDN U7970 ( .A(n7236), .B(n7235), .Z(n7240) );
  NAND U7971 ( .A(n7238), .B(n7237), .Z(n7239) );
  NAND U7972 ( .A(n7240), .B(n7239), .Z(n7256) );
  AND U7973 ( .A(b[2]), .B(a[250]), .Z(n7262) );
  AND U7974 ( .A(a[251]), .B(b[1]), .Z(n7260) );
  AND U7975 ( .A(a[249]), .B(b[3]), .Z(n7259) );
  XOR U7976 ( .A(n7260), .B(n7259), .Z(n7261) );
  XOR U7977 ( .A(n7262), .B(n7261), .Z(n7265) );
  NAND U7978 ( .A(b[0]), .B(a[252]), .Z(n7266) );
  XOR U7979 ( .A(n7265), .B(n7266), .Z(n7268) );
  OR U7980 ( .A(n7242), .B(n7241), .Z(n7246) );
  NANDN U7981 ( .A(n7244), .B(n7243), .Z(n7245) );
  NAND U7982 ( .A(n7246), .B(n7245), .Z(n7267) );
  XNOR U7983 ( .A(n7268), .B(n7267), .Z(n7253) );
  NANDN U7984 ( .A(n7248), .B(n7247), .Z(n7252) );
  OR U7985 ( .A(n7250), .B(n7249), .Z(n7251) );
  NAND U7986 ( .A(n7252), .B(n7251), .Z(n7254) );
  XNOR U7987 ( .A(n7253), .B(n7254), .Z(n7255) );
  XNOR U7988 ( .A(n7256), .B(n7255), .Z(n7271) );
  XNOR U7989 ( .A(n7271), .B(sreg[1272]), .Z(n7273) );
  XNOR U7990 ( .A(n7272), .B(n7273), .Z(c[1272]) );
  NANDN U7991 ( .A(n7254), .B(n7253), .Z(n7258) );
  NAND U7992 ( .A(n7256), .B(n7255), .Z(n7257) );
  NAND U7993 ( .A(n7258), .B(n7257), .Z(n7282) );
  AND U7994 ( .A(b[2]), .B(a[251]), .Z(n7288) );
  AND U7995 ( .A(a[252]), .B(b[1]), .Z(n7286) );
  AND U7996 ( .A(a[250]), .B(b[3]), .Z(n7285) );
  XOR U7997 ( .A(n7286), .B(n7285), .Z(n7287) );
  XOR U7998 ( .A(n7288), .B(n7287), .Z(n7291) );
  NAND U7999 ( .A(b[0]), .B(a[253]), .Z(n7292) );
  XOR U8000 ( .A(n7291), .B(n7292), .Z(n7294) );
  OR U8001 ( .A(n7260), .B(n7259), .Z(n7264) );
  NANDN U8002 ( .A(n7262), .B(n7261), .Z(n7263) );
  NAND U8003 ( .A(n7264), .B(n7263), .Z(n7293) );
  XNOR U8004 ( .A(n7294), .B(n7293), .Z(n7279) );
  NANDN U8005 ( .A(n7266), .B(n7265), .Z(n7270) );
  OR U8006 ( .A(n7268), .B(n7267), .Z(n7269) );
  NAND U8007 ( .A(n7270), .B(n7269), .Z(n7280) );
  XNOR U8008 ( .A(n7279), .B(n7280), .Z(n7281) );
  XOR U8009 ( .A(n7282), .B(n7281), .Z(n7278) );
  NAND U8010 ( .A(n7271), .B(sreg[1272]), .Z(n7275) );
  NANDN U8011 ( .A(n7273), .B(n7272), .Z(n7274) );
  NAND U8012 ( .A(n7275), .B(n7274), .Z(n7277) );
  XNOR U8013 ( .A(sreg[1273]), .B(n7277), .Z(n7276) );
  XOR U8014 ( .A(n7278), .B(n7276), .Z(c[1273]) );
  NANDN U8015 ( .A(n7280), .B(n7279), .Z(n7284) );
  NAND U8016 ( .A(n7282), .B(n7281), .Z(n7283) );
  NAND U8017 ( .A(n7284), .B(n7283), .Z(n7300) );
  AND U8018 ( .A(b[2]), .B(a[252]), .Z(n7306) );
  AND U8019 ( .A(a[253]), .B(b[1]), .Z(n7304) );
  AND U8020 ( .A(a[251]), .B(b[3]), .Z(n7303) );
  XOR U8021 ( .A(n7304), .B(n7303), .Z(n7305) );
  XOR U8022 ( .A(n7306), .B(n7305), .Z(n7309) );
  NAND U8023 ( .A(b[0]), .B(a[254]), .Z(n7310) );
  XOR U8024 ( .A(n7309), .B(n7310), .Z(n7312) );
  OR U8025 ( .A(n7286), .B(n7285), .Z(n7290) );
  NANDN U8026 ( .A(n7288), .B(n7287), .Z(n7289) );
  NAND U8027 ( .A(n7290), .B(n7289), .Z(n7311) );
  XNOR U8028 ( .A(n7312), .B(n7311), .Z(n7297) );
  NANDN U8029 ( .A(n7292), .B(n7291), .Z(n7296) );
  OR U8030 ( .A(n7294), .B(n7293), .Z(n7295) );
  NAND U8031 ( .A(n7296), .B(n7295), .Z(n7298) );
  XNOR U8032 ( .A(n7297), .B(n7298), .Z(n7299) );
  XNOR U8033 ( .A(n7300), .B(n7299), .Z(n7315) );
  XNOR U8034 ( .A(n7315), .B(sreg[1274]), .Z(n7316) );
  XOR U8035 ( .A(n7317), .B(n7316), .Z(c[1274]) );
  NANDN U8036 ( .A(n7298), .B(n7297), .Z(n7302) );
  NAND U8037 ( .A(n7300), .B(n7299), .Z(n7301) );
  NAND U8038 ( .A(n7302), .B(n7301), .Z(n7328) );
  AND U8039 ( .A(b[2]), .B(a[253]), .Z(n7334) );
  AND U8040 ( .A(a[254]), .B(b[1]), .Z(n7332) );
  AND U8041 ( .A(a[252]), .B(b[3]), .Z(n7331) );
  XOR U8042 ( .A(n7332), .B(n7331), .Z(n7333) );
  XOR U8043 ( .A(n7334), .B(n7333), .Z(n7337) );
  NAND U8044 ( .A(b[0]), .B(a[255]), .Z(n7338) );
  XOR U8045 ( .A(n7337), .B(n7338), .Z(n7340) );
  OR U8046 ( .A(n7304), .B(n7303), .Z(n7308) );
  NANDN U8047 ( .A(n7306), .B(n7305), .Z(n7307) );
  NAND U8048 ( .A(n7308), .B(n7307), .Z(n7339) );
  XNOR U8049 ( .A(n7340), .B(n7339), .Z(n7325) );
  NANDN U8050 ( .A(n7310), .B(n7309), .Z(n7314) );
  OR U8051 ( .A(n7312), .B(n7311), .Z(n7313) );
  NAND U8052 ( .A(n7314), .B(n7313), .Z(n7326) );
  XNOR U8053 ( .A(n7325), .B(n7326), .Z(n7327) );
  XNOR U8054 ( .A(n7328), .B(n7327), .Z(n7320) );
  XOR U8055 ( .A(sreg[1275]), .B(n7320), .Z(n7321) );
  NAND U8056 ( .A(n7315), .B(sreg[1274]), .Z(n7319) );
  OR U8057 ( .A(n7317), .B(n7316), .Z(n7318) );
  NAND U8058 ( .A(n7319), .B(n7318), .Z(n7322) );
  XOR U8059 ( .A(n7321), .B(n7322), .Z(c[1275]) );
  OR U8060 ( .A(n7320), .B(sreg[1275]), .Z(n7324) );
  NANDN U8061 ( .A(n7322), .B(n7321), .Z(n7323) );
  NAND U8062 ( .A(n7324), .B(n7323), .Z(n7363) );
  NANDN U8063 ( .A(n7326), .B(n7325), .Z(n7330) );
  NAND U8064 ( .A(n7328), .B(n7327), .Z(n7329) );
  NAND U8065 ( .A(n7330), .B(n7329), .Z(n7346) );
  AND U8066 ( .A(b[2]), .B(a[254]), .Z(n7352) );
  AND U8067 ( .A(a[255]), .B(b[1]), .Z(n7350) );
  AND U8068 ( .A(a[253]), .B(b[3]), .Z(n7349) );
  XOR U8069 ( .A(n7350), .B(n7349), .Z(n7351) );
  XOR U8070 ( .A(n7352), .B(n7351), .Z(n7355) );
  NAND U8071 ( .A(b[0]), .B(a[256]), .Z(n7356) );
  XOR U8072 ( .A(n7355), .B(n7356), .Z(n7358) );
  OR U8073 ( .A(n7332), .B(n7331), .Z(n7336) );
  NANDN U8074 ( .A(n7334), .B(n7333), .Z(n7335) );
  NAND U8075 ( .A(n7336), .B(n7335), .Z(n7357) );
  XNOR U8076 ( .A(n7358), .B(n7357), .Z(n7343) );
  NANDN U8077 ( .A(n7338), .B(n7337), .Z(n7342) );
  OR U8078 ( .A(n7340), .B(n7339), .Z(n7341) );
  NAND U8079 ( .A(n7342), .B(n7341), .Z(n7344) );
  XNOR U8080 ( .A(n7343), .B(n7344), .Z(n7345) );
  XNOR U8081 ( .A(n7346), .B(n7345), .Z(n7361) );
  XNOR U8082 ( .A(n7361), .B(sreg[1276]), .Z(n7362) );
  XOR U8083 ( .A(n7363), .B(n7362), .Z(c[1276]) );
  NANDN U8084 ( .A(n7344), .B(n7343), .Z(n7348) );
  NAND U8085 ( .A(n7346), .B(n7345), .Z(n7347) );
  NAND U8086 ( .A(n7348), .B(n7347), .Z(n7369) );
  AND U8087 ( .A(b[2]), .B(a[255]), .Z(n7375) );
  AND U8088 ( .A(a[256]), .B(b[1]), .Z(n7373) );
  AND U8089 ( .A(a[254]), .B(b[3]), .Z(n7372) );
  XOR U8090 ( .A(n7373), .B(n7372), .Z(n7374) );
  XOR U8091 ( .A(n7375), .B(n7374), .Z(n7378) );
  NAND U8092 ( .A(b[0]), .B(a[257]), .Z(n7379) );
  XOR U8093 ( .A(n7378), .B(n7379), .Z(n7381) );
  OR U8094 ( .A(n7350), .B(n7349), .Z(n7354) );
  NANDN U8095 ( .A(n7352), .B(n7351), .Z(n7353) );
  NAND U8096 ( .A(n7354), .B(n7353), .Z(n7380) );
  XNOR U8097 ( .A(n7381), .B(n7380), .Z(n7366) );
  NANDN U8098 ( .A(n7356), .B(n7355), .Z(n7360) );
  OR U8099 ( .A(n7358), .B(n7357), .Z(n7359) );
  NAND U8100 ( .A(n7360), .B(n7359), .Z(n7367) );
  XNOR U8101 ( .A(n7366), .B(n7367), .Z(n7368) );
  XNOR U8102 ( .A(n7369), .B(n7368), .Z(n7384) );
  XNOR U8103 ( .A(n7384), .B(sreg[1277]), .Z(n7386) );
  NAND U8104 ( .A(n7361), .B(sreg[1276]), .Z(n7365) );
  OR U8105 ( .A(n7363), .B(n7362), .Z(n7364) );
  AND U8106 ( .A(n7365), .B(n7364), .Z(n7385) );
  XOR U8107 ( .A(n7386), .B(n7385), .Z(c[1277]) );
  NANDN U8108 ( .A(n7367), .B(n7366), .Z(n7371) );
  NAND U8109 ( .A(n7369), .B(n7368), .Z(n7370) );
  NAND U8110 ( .A(n7371), .B(n7370), .Z(n7393) );
  AND U8111 ( .A(b[2]), .B(a[256]), .Z(n7399) );
  AND U8112 ( .A(a[257]), .B(b[1]), .Z(n7397) );
  AND U8113 ( .A(a[255]), .B(b[3]), .Z(n7396) );
  XOR U8114 ( .A(n7397), .B(n7396), .Z(n7398) );
  XOR U8115 ( .A(n7399), .B(n7398), .Z(n7402) );
  NAND U8116 ( .A(b[0]), .B(a[258]), .Z(n7403) );
  XOR U8117 ( .A(n7402), .B(n7403), .Z(n7405) );
  OR U8118 ( .A(n7373), .B(n7372), .Z(n7377) );
  NANDN U8119 ( .A(n7375), .B(n7374), .Z(n7376) );
  NAND U8120 ( .A(n7377), .B(n7376), .Z(n7404) );
  XNOR U8121 ( .A(n7405), .B(n7404), .Z(n7390) );
  NANDN U8122 ( .A(n7379), .B(n7378), .Z(n7383) );
  OR U8123 ( .A(n7381), .B(n7380), .Z(n7382) );
  NAND U8124 ( .A(n7383), .B(n7382), .Z(n7391) );
  XNOR U8125 ( .A(n7390), .B(n7391), .Z(n7392) );
  XNOR U8126 ( .A(n7393), .B(n7392), .Z(n7409) );
  NAND U8127 ( .A(n7384), .B(sreg[1277]), .Z(n7388) );
  OR U8128 ( .A(n7386), .B(n7385), .Z(n7387) );
  AND U8129 ( .A(n7388), .B(n7387), .Z(n7408) );
  XNOR U8130 ( .A(n7408), .B(sreg[1278]), .Z(n7389) );
  XOR U8131 ( .A(n7409), .B(n7389), .Z(c[1278]) );
  NANDN U8132 ( .A(n7391), .B(n7390), .Z(n7395) );
  NAND U8133 ( .A(n7393), .B(n7392), .Z(n7394) );
  NAND U8134 ( .A(n7395), .B(n7394), .Z(n7416) );
  AND U8135 ( .A(b[2]), .B(a[257]), .Z(n7422) );
  AND U8136 ( .A(a[258]), .B(b[1]), .Z(n7420) );
  AND U8137 ( .A(a[256]), .B(b[3]), .Z(n7419) );
  XOR U8138 ( .A(n7420), .B(n7419), .Z(n7421) );
  XOR U8139 ( .A(n7422), .B(n7421), .Z(n7425) );
  NAND U8140 ( .A(b[0]), .B(a[259]), .Z(n7426) );
  XOR U8141 ( .A(n7425), .B(n7426), .Z(n7428) );
  OR U8142 ( .A(n7397), .B(n7396), .Z(n7401) );
  NANDN U8143 ( .A(n7399), .B(n7398), .Z(n7400) );
  NAND U8144 ( .A(n7401), .B(n7400), .Z(n7427) );
  XNOR U8145 ( .A(n7428), .B(n7427), .Z(n7413) );
  NANDN U8146 ( .A(n7403), .B(n7402), .Z(n7407) );
  OR U8147 ( .A(n7405), .B(n7404), .Z(n7406) );
  NAND U8148 ( .A(n7407), .B(n7406), .Z(n7414) );
  XNOR U8149 ( .A(n7413), .B(n7414), .Z(n7415) );
  XNOR U8150 ( .A(n7416), .B(n7415), .Z(n7412) );
  XOR U8151 ( .A(n7411), .B(sreg[1279]), .Z(n7410) );
  XOR U8152 ( .A(n7412), .B(n7410), .Z(c[1279]) );
  NANDN U8153 ( .A(n7414), .B(n7413), .Z(n7418) );
  NAND U8154 ( .A(n7416), .B(n7415), .Z(n7417) );
  NAND U8155 ( .A(n7418), .B(n7417), .Z(n7434) );
  AND U8156 ( .A(b[2]), .B(a[258]), .Z(n7440) );
  AND U8157 ( .A(a[259]), .B(b[1]), .Z(n7438) );
  AND U8158 ( .A(a[257]), .B(b[3]), .Z(n7437) );
  XOR U8159 ( .A(n7438), .B(n7437), .Z(n7439) );
  XOR U8160 ( .A(n7440), .B(n7439), .Z(n7443) );
  NAND U8161 ( .A(b[0]), .B(a[260]), .Z(n7444) );
  XOR U8162 ( .A(n7443), .B(n7444), .Z(n7446) );
  OR U8163 ( .A(n7420), .B(n7419), .Z(n7424) );
  NANDN U8164 ( .A(n7422), .B(n7421), .Z(n7423) );
  NAND U8165 ( .A(n7424), .B(n7423), .Z(n7445) );
  XNOR U8166 ( .A(n7446), .B(n7445), .Z(n7431) );
  NANDN U8167 ( .A(n7426), .B(n7425), .Z(n7430) );
  OR U8168 ( .A(n7428), .B(n7427), .Z(n7429) );
  NAND U8169 ( .A(n7430), .B(n7429), .Z(n7432) );
  XNOR U8170 ( .A(n7431), .B(n7432), .Z(n7433) );
  XNOR U8171 ( .A(n7434), .B(n7433), .Z(n7449) );
  XOR U8172 ( .A(sreg[1280]), .B(n7449), .Z(n7450) );
  XOR U8173 ( .A(n7451), .B(n7450), .Z(c[1280]) );
  NANDN U8174 ( .A(n7432), .B(n7431), .Z(n7436) );
  NAND U8175 ( .A(n7434), .B(n7433), .Z(n7435) );
  NAND U8176 ( .A(n7436), .B(n7435), .Z(n7458) );
  AND U8177 ( .A(b[2]), .B(a[259]), .Z(n7464) );
  AND U8178 ( .A(a[260]), .B(b[1]), .Z(n7462) );
  AND U8179 ( .A(a[258]), .B(b[3]), .Z(n7461) );
  XOR U8180 ( .A(n7462), .B(n7461), .Z(n7463) );
  XOR U8181 ( .A(n7464), .B(n7463), .Z(n7467) );
  NAND U8182 ( .A(b[0]), .B(a[261]), .Z(n7468) );
  XOR U8183 ( .A(n7467), .B(n7468), .Z(n7470) );
  OR U8184 ( .A(n7438), .B(n7437), .Z(n7442) );
  NANDN U8185 ( .A(n7440), .B(n7439), .Z(n7441) );
  NAND U8186 ( .A(n7442), .B(n7441), .Z(n7469) );
  XNOR U8187 ( .A(n7470), .B(n7469), .Z(n7455) );
  NANDN U8188 ( .A(n7444), .B(n7443), .Z(n7448) );
  OR U8189 ( .A(n7446), .B(n7445), .Z(n7447) );
  NAND U8190 ( .A(n7448), .B(n7447), .Z(n7456) );
  XNOR U8191 ( .A(n7455), .B(n7456), .Z(n7457) );
  XOR U8192 ( .A(n7458), .B(n7457), .Z(n7474) );
  OR U8193 ( .A(n7449), .B(sreg[1280]), .Z(n7453) );
  NANDN U8194 ( .A(n7451), .B(n7450), .Z(n7452) );
  AND U8195 ( .A(n7453), .B(n7452), .Z(n7473) );
  XNOR U8196 ( .A(sreg[1281]), .B(n7473), .Z(n7454) );
  XOR U8197 ( .A(n7474), .B(n7454), .Z(c[1281]) );
  NANDN U8198 ( .A(n7456), .B(n7455), .Z(n7460) );
  NAND U8199 ( .A(n7458), .B(n7457), .Z(n7459) );
  NAND U8200 ( .A(n7460), .B(n7459), .Z(n7479) );
  AND U8201 ( .A(b[2]), .B(a[260]), .Z(n7485) );
  AND U8202 ( .A(a[261]), .B(b[1]), .Z(n7483) );
  AND U8203 ( .A(a[259]), .B(b[3]), .Z(n7482) );
  XOR U8204 ( .A(n7483), .B(n7482), .Z(n7484) );
  XOR U8205 ( .A(n7485), .B(n7484), .Z(n7488) );
  NAND U8206 ( .A(b[0]), .B(a[262]), .Z(n7489) );
  XOR U8207 ( .A(n7488), .B(n7489), .Z(n7491) );
  OR U8208 ( .A(n7462), .B(n7461), .Z(n7466) );
  NANDN U8209 ( .A(n7464), .B(n7463), .Z(n7465) );
  NAND U8210 ( .A(n7466), .B(n7465), .Z(n7490) );
  XNOR U8211 ( .A(n7491), .B(n7490), .Z(n7476) );
  NANDN U8212 ( .A(n7468), .B(n7467), .Z(n7472) );
  OR U8213 ( .A(n7470), .B(n7469), .Z(n7471) );
  NAND U8214 ( .A(n7472), .B(n7471), .Z(n7477) );
  XNOR U8215 ( .A(n7476), .B(n7477), .Z(n7478) );
  XOR U8216 ( .A(n7479), .B(n7478), .Z(n7495) );
  XNOR U8217 ( .A(sreg[1282]), .B(n7494), .Z(n7475) );
  XOR U8218 ( .A(n7495), .B(n7475), .Z(c[1282]) );
  NANDN U8219 ( .A(n7477), .B(n7476), .Z(n7481) );
  NAND U8220 ( .A(n7479), .B(n7478), .Z(n7480) );
  NAND U8221 ( .A(n7481), .B(n7480), .Z(n7500) );
  AND U8222 ( .A(b[2]), .B(a[261]), .Z(n7506) );
  AND U8223 ( .A(a[262]), .B(b[1]), .Z(n7504) );
  AND U8224 ( .A(a[260]), .B(b[3]), .Z(n7503) );
  XOR U8225 ( .A(n7504), .B(n7503), .Z(n7505) );
  XOR U8226 ( .A(n7506), .B(n7505), .Z(n7509) );
  NAND U8227 ( .A(b[0]), .B(a[263]), .Z(n7510) );
  XOR U8228 ( .A(n7509), .B(n7510), .Z(n7512) );
  OR U8229 ( .A(n7483), .B(n7482), .Z(n7487) );
  NANDN U8230 ( .A(n7485), .B(n7484), .Z(n7486) );
  NAND U8231 ( .A(n7487), .B(n7486), .Z(n7511) );
  XNOR U8232 ( .A(n7512), .B(n7511), .Z(n7497) );
  NANDN U8233 ( .A(n7489), .B(n7488), .Z(n7493) );
  OR U8234 ( .A(n7491), .B(n7490), .Z(n7492) );
  NAND U8235 ( .A(n7493), .B(n7492), .Z(n7498) );
  XNOR U8236 ( .A(n7497), .B(n7498), .Z(n7499) );
  XOR U8237 ( .A(n7500), .B(n7499), .Z(n7516) );
  XNOR U8238 ( .A(sreg[1283]), .B(n7515), .Z(n7496) );
  XOR U8239 ( .A(n7516), .B(n7496), .Z(c[1283]) );
  NANDN U8240 ( .A(n7498), .B(n7497), .Z(n7502) );
  NAND U8241 ( .A(n7500), .B(n7499), .Z(n7501) );
  NAND U8242 ( .A(n7502), .B(n7501), .Z(n7521) );
  AND U8243 ( .A(b[2]), .B(a[262]), .Z(n7527) );
  AND U8244 ( .A(a[263]), .B(b[1]), .Z(n7525) );
  AND U8245 ( .A(a[261]), .B(b[3]), .Z(n7524) );
  XOR U8246 ( .A(n7525), .B(n7524), .Z(n7526) );
  XOR U8247 ( .A(n7527), .B(n7526), .Z(n7530) );
  NAND U8248 ( .A(b[0]), .B(a[264]), .Z(n7531) );
  XOR U8249 ( .A(n7530), .B(n7531), .Z(n7533) );
  OR U8250 ( .A(n7504), .B(n7503), .Z(n7508) );
  NANDN U8251 ( .A(n7506), .B(n7505), .Z(n7507) );
  NAND U8252 ( .A(n7508), .B(n7507), .Z(n7532) );
  XNOR U8253 ( .A(n7533), .B(n7532), .Z(n7518) );
  NANDN U8254 ( .A(n7510), .B(n7509), .Z(n7514) );
  OR U8255 ( .A(n7512), .B(n7511), .Z(n7513) );
  NAND U8256 ( .A(n7514), .B(n7513), .Z(n7519) );
  XNOR U8257 ( .A(n7518), .B(n7519), .Z(n7520) );
  XOR U8258 ( .A(n7521), .B(n7520), .Z(n7537) );
  XNOR U8259 ( .A(sreg[1284]), .B(n7536), .Z(n7517) );
  XOR U8260 ( .A(n7537), .B(n7517), .Z(c[1284]) );
  NANDN U8261 ( .A(n7519), .B(n7518), .Z(n7523) );
  NAND U8262 ( .A(n7521), .B(n7520), .Z(n7522) );
  NAND U8263 ( .A(n7523), .B(n7522), .Z(n7544) );
  AND U8264 ( .A(b[2]), .B(a[263]), .Z(n7550) );
  AND U8265 ( .A(a[264]), .B(b[1]), .Z(n7548) );
  AND U8266 ( .A(a[262]), .B(b[3]), .Z(n7547) );
  XOR U8267 ( .A(n7548), .B(n7547), .Z(n7549) );
  XOR U8268 ( .A(n7550), .B(n7549), .Z(n7553) );
  NAND U8269 ( .A(b[0]), .B(a[265]), .Z(n7554) );
  XOR U8270 ( .A(n7553), .B(n7554), .Z(n7556) );
  OR U8271 ( .A(n7525), .B(n7524), .Z(n7529) );
  NANDN U8272 ( .A(n7527), .B(n7526), .Z(n7528) );
  NAND U8273 ( .A(n7529), .B(n7528), .Z(n7555) );
  XNOR U8274 ( .A(n7556), .B(n7555), .Z(n7541) );
  NANDN U8275 ( .A(n7531), .B(n7530), .Z(n7535) );
  OR U8276 ( .A(n7533), .B(n7532), .Z(n7534) );
  NAND U8277 ( .A(n7535), .B(n7534), .Z(n7542) );
  XNOR U8278 ( .A(n7541), .B(n7542), .Z(n7543) );
  XNOR U8279 ( .A(n7544), .B(n7543), .Z(n7540) );
  XOR U8280 ( .A(n7539), .B(sreg[1285]), .Z(n7538) );
  XOR U8281 ( .A(n7540), .B(n7538), .Z(c[1285]) );
  NANDN U8282 ( .A(n7542), .B(n7541), .Z(n7546) );
  NAND U8283 ( .A(n7544), .B(n7543), .Z(n7545) );
  NAND U8284 ( .A(n7546), .B(n7545), .Z(n7562) );
  AND U8285 ( .A(b[2]), .B(a[264]), .Z(n7568) );
  AND U8286 ( .A(a[265]), .B(b[1]), .Z(n7566) );
  AND U8287 ( .A(a[263]), .B(b[3]), .Z(n7565) );
  XOR U8288 ( .A(n7566), .B(n7565), .Z(n7567) );
  XOR U8289 ( .A(n7568), .B(n7567), .Z(n7571) );
  NAND U8290 ( .A(b[0]), .B(a[266]), .Z(n7572) );
  XOR U8291 ( .A(n7571), .B(n7572), .Z(n7574) );
  OR U8292 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U8293 ( .A(n7550), .B(n7549), .Z(n7551) );
  NAND U8294 ( .A(n7552), .B(n7551), .Z(n7573) );
  XNOR U8295 ( .A(n7574), .B(n7573), .Z(n7559) );
  NANDN U8296 ( .A(n7554), .B(n7553), .Z(n7558) );
  OR U8297 ( .A(n7556), .B(n7555), .Z(n7557) );
  NAND U8298 ( .A(n7558), .B(n7557), .Z(n7560) );
  XNOR U8299 ( .A(n7559), .B(n7560), .Z(n7561) );
  XNOR U8300 ( .A(n7562), .B(n7561), .Z(n7577) );
  XNOR U8301 ( .A(n7577), .B(sreg[1286]), .Z(n7579) );
  XNOR U8302 ( .A(n7578), .B(n7579), .Z(c[1286]) );
  NANDN U8303 ( .A(n7560), .B(n7559), .Z(n7564) );
  NAND U8304 ( .A(n7562), .B(n7561), .Z(n7563) );
  NAND U8305 ( .A(n7564), .B(n7563), .Z(n7586) );
  AND U8306 ( .A(b[2]), .B(a[265]), .Z(n7592) );
  AND U8307 ( .A(a[266]), .B(b[1]), .Z(n7590) );
  AND U8308 ( .A(a[264]), .B(b[3]), .Z(n7589) );
  XOR U8309 ( .A(n7590), .B(n7589), .Z(n7591) );
  XOR U8310 ( .A(n7592), .B(n7591), .Z(n7595) );
  NAND U8311 ( .A(b[0]), .B(a[267]), .Z(n7596) );
  XOR U8312 ( .A(n7595), .B(n7596), .Z(n7598) );
  OR U8313 ( .A(n7566), .B(n7565), .Z(n7570) );
  NANDN U8314 ( .A(n7568), .B(n7567), .Z(n7569) );
  NAND U8315 ( .A(n7570), .B(n7569), .Z(n7597) );
  XNOR U8316 ( .A(n7598), .B(n7597), .Z(n7583) );
  NANDN U8317 ( .A(n7572), .B(n7571), .Z(n7576) );
  OR U8318 ( .A(n7574), .B(n7573), .Z(n7575) );
  NAND U8319 ( .A(n7576), .B(n7575), .Z(n7584) );
  XNOR U8320 ( .A(n7583), .B(n7584), .Z(n7585) );
  XNOR U8321 ( .A(n7586), .B(n7585), .Z(n7602) );
  NAND U8322 ( .A(n7577), .B(sreg[1286]), .Z(n7581) );
  NANDN U8323 ( .A(n7579), .B(n7578), .Z(n7580) );
  AND U8324 ( .A(n7581), .B(n7580), .Z(n7601) );
  XNOR U8325 ( .A(n7601), .B(sreg[1287]), .Z(n7582) );
  XOR U8326 ( .A(n7602), .B(n7582), .Z(c[1287]) );
  NANDN U8327 ( .A(n7584), .B(n7583), .Z(n7588) );
  NAND U8328 ( .A(n7586), .B(n7585), .Z(n7587) );
  NAND U8329 ( .A(n7588), .B(n7587), .Z(n7609) );
  AND U8330 ( .A(b[2]), .B(a[266]), .Z(n7615) );
  AND U8331 ( .A(a[267]), .B(b[1]), .Z(n7613) );
  AND U8332 ( .A(a[265]), .B(b[3]), .Z(n7612) );
  XOR U8333 ( .A(n7613), .B(n7612), .Z(n7614) );
  XOR U8334 ( .A(n7615), .B(n7614), .Z(n7618) );
  NAND U8335 ( .A(b[0]), .B(a[268]), .Z(n7619) );
  XOR U8336 ( .A(n7618), .B(n7619), .Z(n7621) );
  OR U8337 ( .A(n7590), .B(n7589), .Z(n7594) );
  NANDN U8338 ( .A(n7592), .B(n7591), .Z(n7593) );
  NAND U8339 ( .A(n7594), .B(n7593), .Z(n7620) );
  XNOR U8340 ( .A(n7621), .B(n7620), .Z(n7606) );
  NANDN U8341 ( .A(n7596), .B(n7595), .Z(n7600) );
  OR U8342 ( .A(n7598), .B(n7597), .Z(n7599) );
  NAND U8343 ( .A(n7600), .B(n7599), .Z(n7607) );
  XNOR U8344 ( .A(n7606), .B(n7607), .Z(n7608) );
  XOR U8345 ( .A(n7609), .B(n7608), .Z(n7605) );
  XOR U8346 ( .A(sreg[1288]), .B(n7604), .Z(n7603) );
  XOR U8347 ( .A(n7605), .B(n7603), .Z(c[1288]) );
  NANDN U8348 ( .A(n7607), .B(n7606), .Z(n7611) );
  NAND U8349 ( .A(n7609), .B(n7608), .Z(n7610) );
  NAND U8350 ( .A(n7611), .B(n7610), .Z(n7627) );
  AND U8351 ( .A(b[2]), .B(a[267]), .Z(n7633) );
  AND U8352 ( .A(a[268]), .B(b[1]), .Z(n7631) );
  AND U8353 ( .A(a[266]), .B(b[3]), .Z(n7630) );
  XOR U8354 ( .A(n7631), .B(n7630), .Z(n7632) );
  XOR U8355 ( .A(n7633), .B(n7632), .Z(n7636) );
  NAND U8356 ( .A(b[0]), .B(a[269]), .Z(n7637) );
  XOR U8357 ( .A(n7636), .B(n7637), .Z(n7639) );
  OR U8358 ( .A(n7613), .B(n7612), .Z(n7617) );
  NANDN U8359 ( .A(n7615), .B(n7614), .Z(n7616) );
  NAND U8360 ( .A(n7617), .B(n7616), .Z(n7638) );
  XNOR U8361 ( .A(n7639), .B(n7638), .Z(n7624) );
  NANDN U8362 ( .A(n7619), .B(n7618), .Z(n7623) );
  OR U8363 ( .A(n7621), .B(n7620), .Z(n7622) );
  NAND U8364 ( .A(n7623), .B(n7622), .Z(n7625) );
  XNOR U8365 ( .A(n7624), .B(n7625), .Z(n7626) );
  XNOR U8366 ( .A(n7627), .B(n7626), .Z(n7642) );
  XNOR U8367 ( .A(n7642), .B(sreg[1289]), .Z(n7643) );
  XOR U8368 ( .A(n7644), .B(n7643), .Z(c[1289]) );
  NANDN U8369 ( .A(n7625), .B(n7624), .Z(n7629) );
  NAND U8370 ( .A(n7627), .B(n7626), .Z(n7628) );
  NAND U8371 ( .A(n7629), .B(n7628), .Z(n7651) );
  AND U8372 ( .A(b[2]), .B(a[268]), .Z(n7657) );
  AND U8373 ( .A(a[269]), .B(b[1]), .Z(n7655) );
  AND U8374 ( .A(a[267]), .B(b[3]), .Z(n7654) );
  XOR U8375 ( .A(n7655), .B(n7654), .Z(n7656) );
  XOR U8376 ( .A(n7657), .B(n7656), .Z(n7660) );
  NAND U8377 ( .A(b[0]), .B(a[270]), .Z(n7661) );
  XOR U8378 ( .A(n7660), .B(n7661), .Z(n7663) );
  OR U8379 ( .A(n7631), .B(n7630), .Z(n7635) );
  NANDN U8380 ( .A(n7633), .B(n7632), .Z(n7634) );
  NAND U8381 ( .A(n7635), .B(n7634), .Z(n7662) );
  XNOR U8382 ( .A(n7663), .B(n7662), .Z(n7648) );
  NANDN U8383 ( .A(n7637), .B(n7636), .Z(n7641) );
  OR U8384 ( .A(n7639), .B(n7638), .Z(n7640) );
  NAND U8385 ( .A(n7641), .B(n7640), .Z(n7649) );
  XNOR U8386 ( .A(n7648), .B(n7649), .Z(n7650) );
  XNOR U8387 ( .A(n7651), .B(n7650), .Z(n7667) );
  NAND U8388 ( .A(n7642), .B(sreg[1289]), .Z(n7646) );
  OR U8389 ( .A(n7644), .B(n7643), .Z(n7645) );
  AND U8390 ( .A(n7646), .B(n7645), .Z(n7666) );
  XNOR U8391 ( .A(n7666), .B(sreg[1290]), .Z(n7647) );
  XOR U8392 ( .A(n7667), .B(n7647), .Z(c[1290]) );
  NANDN U8393 ( .A(n7649), .B(n7648), .Z(n7653) );
  NAND U8394 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U8395 ( .A(n7653), .B(n7652), .Z(n7672) );
  AND U8396 ( .A(b[2]), .B(a[269]), .Z(n7678) );
  AND U8397 ( .A(a[270]), .B(b[1]), .Z(n7676) );
  AND U8398 ( .A(a[268]), .B(b[3]), .Z(n7675) );
  XOR U8399 ( .A(n7676), .B(n7675), .Z(n7677) );
  XOR U8400 ( .A(n7678), .B(n7677), .Z(n7681) );
  NAND U8401 ( .A(b[0]), .B(a[271]), .Z(n7682) );
  XOR U8402 ( .A(n7681), .B(n7682), .Z(n7684) );
  OR U8403 ( .A(n7655), .B(n7654), .Z(n7659) );
  NANDN U8404 ( .A(n7657), .B(n7656), .Z(n7658) );
  NAND U8405 ( .A(n7659), .B(n7658), .Z(n7683) );
  XNOR U8406 ( .A(n7684), .B(n7683), .Z(n7669) );
  NANDN U8407 ( .A(n7661), .B(n7660), .Z(n7665) );
  OR U8408 ( .A(n7663), .B(n7662), .Z(n7664) );
  NAND U8409 ( .A(n7665), .B(n7664), .Z(n7670) );
  XNOR U8410 ( .A(n7669), .B(n7670), .Z(n7671) );
  XOR U8411 ( .A(n7672), .B(n7671), .Z(n7688) );
  XOR U8412 ( .A(sreg[1291]), .B(n7687), .Z(n7668) );
  XOR U8413 ( .A(n7688), .B(n7668), .Z(c[1291]) );
  NANDN U8414 ( .A(n7670), .B(n7669), .Z(n7674) );
  NAND U8415 ( .A(n7672), .B(n7671), .Z(n7673) );
  NAND U8416 ( .A(n7674), .B(n7673), .Z(n7695) );
  AND U8417 ( .A(b[2]), .B(a[270]), .Z(n7707) );
  AND U8418 ( .A(a[271]), .B(b[1]), .Z(n7705) );
  AND U8419 ( .A(a[269]), .B(b[3]), .Z(n7704) );
  XOR U8420 ( .A(n7705), .B(n7704), .Z(n7706) );
  XOR U8421 ( .A(n7707), .B(n7706), .Z(n7698) );
  NAND U8422 ( .A(b[0]), .B(a[272]), .Z(n7699) );
  XOR U8423 ( .A(n7698), .B(n7699), .Z(n7701) );
  OR U8424 ( .A(n7676), .B(n7675), .Z(n7680) );
  NANDN U8425 ( .A(n7678), .B(n7677), .Z(n7679) );
  NAND U8426 ( .A(n7680), .B(n7679), .Z(n7700) );
  XNOR U8427 ( .A(n7701), .B(n7700), .Z(n7692) );
  NANDN U8428 ( .A(n7682), .B(n7681), .Z(n7686) );
  OR U8429 ( .A(n7684), .B(n7683), .Z(n7685) );
  NAND U8430 ( .A(n7686), .B(n7685), .Z(n7693) );
  XNOR U8431 ( .A(n7692), .B(n7693), .Z(n7694) );
  XOR U8432 ( .A(n7695), .B(n7694), .Z(n7691) );
  XNOR U8433 ( .A(sreg[1292]), .B(n7690), .Z(n7689) );
  XOR U8434 ( .A(n7691), .B(n7689), .Z(c[1292]) );
  IV U8435 ( .A(sreg[1293]), .Z(n7712) );
  NANDN U8436 ( .A(n7693), .B(n7692), .Z(n7697) );
  NAND U8437 ( .A(n7695), .B(n7694), .Z(n7696) );
  AND U8438 ( .A(n7697), .B(n7696), .Z(n7720) );
  NANDN U8439 ( .A(n7699), .B(n7698), .Z(n7703) );
  OR U8440 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U8441 ( .A(n7703), .B(n7702), .Z(n7719) );
  AND U8442 ( .A(b[2]), .B(a[271]), .Z(n7724) );
  AND U8443 ( .A(a[272]), .B(b[1]), .Z(n7722) );
  AND U8444 ( .A(a[270]), .B(b[3]), .Z(n7721) );
  XOR U8445 ( .A(n7722), .B(n7721), .Z(n7723) );
  XOR U8446 ( .A(n7724), .B(n7723), .Z(n7727) );
  NAND U8447 ( .A(b[0]), .B(a[273]), .Z(n7728) );
  XOR U8448 ( .A(n7727), .B(n7728), .Z(n7730) );
  OR U8449 ( .A(n7705), .B(n7704), .Z(n7709) );
  NANDN U8450 ( .A(n7707), .B(n7706), .Z(n7708) );
  NAND U8451 ( .A(n7709), .B(n7708), .Z(n7729) );
  XOR U8452 ( .A(n7730), .B(n7729), .Z(n7718) );
  XNOR U8453 ( .A(n7719), .B(n7718), .Z(n7710) );
  XOR U8454 ( .A(n7720), .B(n7710), .Z(n7713) );
  XOR U8455 ( .A(n7712), .B(n7713), .Z(n7711) );
  XOR U8456 ( .A(n7714), .B(n7711), .Z(c[1293]) );
  NANDN U8457 ( .A(n7713), .B(n7712), .Z(n7717) );
  AND U8458 ( .A(n7713), .B(sreg[1293]), .Z(n7715) );
  NANDN U8459 ( .A(n7715), .B(n7714), .Z(n7716) );
  NAND U8460 ( .A(n7717), .B(n7716), .Z(n7753) );
  AND U8461 ( .A(b[2]), .B(a[272]), .Z(n7742) );
  AND U8462 ( .A(a[273]), .B(b[1]), .Z(n7740) );
  AND U8463 ( .A(a[271]), .B(b[3]), .Z(n7739) );
  XOR U8464 ( .A(n7740), .B(n7739), .Z(n7741) );
  XOR U8465 ( .A(n7742), .B(n7741), .Z(n7745) );
  NAND U8466 ( .A(b[0]), .B(a[274]), .Z(n7746) );
  XOR U8467 ( .A(n7745), .B(n7746), .Z(n7748) );
  OR U8468 ( .A(n7722), .B(n7721), .Z(n7726) );
  NANDN U8469 ( .A(n7724), .B(n7723), .Z(n7725) );
  NAND U8470 ( .A(n7726), .B(n7725), .Z(n7747) );
  XNOR U8471 ( .A(n7748), .B(n7747), .Z(n7733) );
  NANDN U8472 ( .A(n7728), .B(n7727), .Z(n7732) );
  OR U8473 ( .A(n7730), .B(n7729), .Z(n7731) );
  NAND U8474 ( .A(n7732), .B(n7731), .Z(n7734) );
  XNOR U8475 ( .A(n7733), .B(n7734), .Z(n7735) );
  XOR U8476 ( .A(n7736), .B(n7735), .Z(n7751) );
  XNOR U8477 ( .A(n7751), .B(sreg[1294]), .Z(n7752) );
  XOR U8478 ( .A(n7753), .B(n7752), .Z(c[1294]) );
  NANDN U8479 ( .A(n7734), .B(n7733), .Z(n7738) );
  NANDN U8480 ( .A(n7736), .B(n7735), .Z(n7737) );
  NAND U8481 ( .A(n7738), .B(n7737), .Z(n7762) );
  AND U8482 ( .A(b[2]), .B(a[273]), .Z(n7768) );
  AND U8483 ( .A(a[274]), .B(b[1]), .Z(n7766) );
  AND U8484 ( .A(a[272]), .B(b[3]), .Z(n7765) );
  XOR U8485 ( .A(n7766), .B(n7765), .Z(n7767) );
  XOR U8486 ( .A(n7768), .B(n7767), .Z(n7771) );
  NAND U8487 ( .A(b[0]), .B(a[275]), .Z(n7772) );
  XOR U8488 ( .A(n7771), .B(n7772), .Z(n7774) );
  OR U8489 ( .A(n7740), .B(n7739), .Z(n7744) );
  NANDN U8490 ( .A(n7742), .B(n7741), .Z(n7743) );
  NAND U8491 ( .A(n7744), .B(n7743), .Z(n7773) );
  XNOR U8492 ( .A(n7774), .B(n7773), .Z(n7759) );
  NANDN U8493 ( .A(n7746), .B(n7745), .Z(n7750) );
  OR U8494 ( .A(n7748), .B(n7747), .Z(n7749) );
  NAND U8495 ( .A(n7750), .B(n7749), .Z(n7760) );
  XNOR U8496 ( .A(n7759), .B(n7760), .Z(n7761) );
  XNOR U8497 ( .A(n7762), .B(n7761), .Z(n7758) );
  NAND U8498 ( .A(n7751), .B(sreg[1294]), .Z(n7755) );
  OR U8499 ( .A(n7753), .B(n7752), .Z(n7754) );
  AND U8500 ( .A(n7755), .B(n7754), .Z(n7757) );
  XNOR U8501 ( .A(n7757), .B(sreg[1295]), .Z(n7756) );
  XOR U8502 ( .A(n7758), .B(n7756), .Z(c[1295]) );
  NANDN U8503 ( .A(n7760), .B(n7759), .Z(n7764) );
  NAND U8504 ( .A(n7762), .B(n7761), .Z(n7763) );
  AND U8505 ( .A(n7764), .B(n7763), .Z(n7780) );
  AND U8506 ( .A(b[2]), .B(a[274]), .Z(n7784) );
  AND U8507 ( .A(a[275]), .B(b[1]), .Z(n7782) );
  AND U8508 ( .A(a[273]), .B(b[3]), .Z(n7781) );
  XOR U8509 ( .A(n7782), .B(n7781), .Z(n7783) );
  XOR U8510 ( .A(n7784), .B(n7783), .Z(n7787) );
  NAND U8511 ( .A(b[0]), .B(a[276]), .Z(n7788) );
  XOR U8512 ( .A(n7787), .B(n7788), .Z(n7789) );
  OR U8513 ( .A(n7766), .B(n7765), .Z(n7770) );
  NANDN U8514 ( .A(n7768), .B(n7767), .Z(n7769) );
  AND U8515 ( .A(n7770), .B(n7769), .Z(n7790) );
  XOR U8516 ( .A(n7789), .B(n7790), .Z(n7778) );
  NANDN U8517 ( .A(n7772), .B(n7771), .Z(n7776) );
  OR U8518 ( .A(n7774), .B(n7773), .Z(n7775) );
  AND U8519 ( .A(n7776), .B(n7775), .Z(n7779) );
  XOR U8520 ( .A(n7778), .B(n7779), .Z(n7777) );
  XOR U8521 ( .A(n7780), .B(n7777), .Z(n7791) );
  XNOR U8522 ( .A(sreg[1296]), .B(n7791), .Z(n7793) );
  XNOR U8523 ( .A(n7792), .B(n7793), .Z(c[1296]) );
  AND U8524 ( .A(b[2]), .B(a[275]), .Z(n7806) );
  AND U8525 ( .A(a[276]), .B(b[1]), .Z(n7804) );
  AND U8526 ( .A(a[274]), .B(b[3]), .Z(n7803) );
  XOR U8527 ( .A(n7804), .B(n7803), .Z(n7805) );
  XOR U8528 ( .A(n7806), .B(n7805), .Z(n7809) );
  NAND U8529 ( .A(b[0]), .B(a[277]), .Z(n7810) );
  XOR U8530 ( .A(n7809), .B(n7810), .Z(n7812) );
  OR U8531 ( .A(n7782), .B(n7781), .Z(n7786) );
  NANDN U8532 ( .A(n7784), .B(n7783), .Z(n7785) );
  NAND U8533 ( .A(n7786), .B(n7785), .Z(n7811) );
  XNOR U8534 ( .A(n7812), .B(n7811), .Z(n7797) );
  XNOR U8535 ( .A(n7797), .B(n7798), .Z(n7800) );
  XOR U8536 ( .A(n7799), .B(n7800), .Z(n7816) );
  NAND U8537 ( .A(sreg[1296]), .B(n7791), .Z(n7795) );
  NANDN U8538 ( .A(n7793), .B(n7792), .Z(n7794) );
  NAND U8539 ( .A(n7795), .B(n7794), .Z(n7815) );
  XNOR U8540 ( .A(sreg[1297]), .B(n7815), .Z(n7796) );
  XOR U8541 ( .A(n7816), .B(n7796), .Z(c[1297]) );
  NANDN U8542 ( .A(n7798), .B(n7797), .Z(n7802) );
  NAND U8543 ( .A(n7800), .B(n7799), .Z(n7801) );
  NAND U8544 ( .A(n7802), .B(n7801), .Z(n7835) );
  AND U8545 ( .A(b[2]), .B(a[276]), .Z(n7829) );
  AND U8546 ( .A(a[277]), .B(b[1]), .Z(n7827) );
  AND U8547 ( .A(a[275]), .B(b[3]), .Z(n7826) );
  XOR U8548 ( .A(n7827), .B(n7826), .Z(n7828) );
  XOR U8549 ( .A(n7829), .B(n7828), .Z(n7820) );
  NAND U8550 ( .A(b[0]), .B(a[278]), .Z(n7821) );
  XOR U8551 ( .A(n7820), .B(n7821), .Z(n7823) );
  OR U8552 ( .A(n7804), .B(n7803), .Z(n7808) );
  NANDN U8553 ( .A(n7806), .B(n7805), .Z(n7807) );
  NAND U8554 ( .A(n7808), .B(n7807), .Z(n7822) );
  XNOR U8555 ( .A(n7823), .B(n7822), .Z(n7832) );
  NANDN U8556 ( .A(n7810), .B(n7809), .Z(n7814) );
  OR U8557 ( .A(n7812), .B(n7811), .Z(n7813) );
  NAND U8558 ( .A(n7814), .B(n7813), .Z(n7833) );
  XNOR U8559 ( .A(n7832), .B(n7833), .Z(n7834) );
  XNOR U8560 ( .A(n7835), .B(n7834), .Z(n7819) );
  XOR U8561 ( .A(n7818), .B(sreg[1298]), .Z(n7817) );
  XOR U8562 ( .A(n7819), .B(n7817), .Z(c[1298]) );
  NANDN U8563 ( .A(n7821), .B(n7820), .Z(n7825) );
  OR U8564 ( .A(n7823), .B(n7822), .Z(n7824) );
  NAND U8565 ( .A(n7825), .B(n7824), .Z(n7850) );
  AND U8566 ( .A(b[2]), .B(a[277]), .Z(n7841) );
  AND U8567 ( .A(a[278]), .B(b[1]), .Z(n7839) );
  AND U8568 ( .A(a[276]), .B(b[3]), .Z(n7838) );
  XOR U8569 ( .A(n7839), .B(n7838), .Z(n7840) );
  XOR U8570 ( .A(n7841), .B(n7840), .Z(n7844) );
  NAND U8571 ( .A(b[0]), .B(a[279]), .Z(n7845) );
  XNOR U8572 ( .A(n7844), .B(n7845), .Z(n7846) );
  OR U8573 ( .A(n7827), .B(n7826), .Z(n7831) );
  NANDN U8574 ( .A(n7829), .B(n7828), .Z(n7830) );
  AND U8575 ( .A(n7831), .B(n7830), .Z(n7847) );
  XNOR U8576 ( .A(n7846), .B(n7847), .Z(n7851) );
  XNOR U8577 ( .A(n7850), .B(n7851), .Z(n7852) );
  NANDN U8578 ( .A(n7833), .B(n7832), .Z(n7837) );
  NAND U8579 ( .A(n7835), .B(n7834), .Z(n7836) );
  AND U8580 ( .A(n7837), .B(n7836), .Z(n7853) );
  XOR U8581 ( .A(n7852), .B(n7853), .Z(n7856) );
  XNOR U8582 ( .A(sreg[1299]), .B(n7856), .Z(n7858) );
  XNOR U8583 ( .A(n7857), .B(n7858), .Z(c[1299]) );
  AND U8584 ( .A(b[2]), .B(a[278]), .Z(n7873) );
  AND U8585 ( .A(a[279]), .B(b[1]), .Z(n7871) );
  AND U8586 ( .A(a[277]), .B(b[3]), .Z(n7870) );
  XOR U8587 ( .A(n7871), .B(n7870), .Z(n7872) );
  XOR U8588 ( .A(n7873), .B(n7872), .Z(n7876) );
  NAND U8589 ( .A(b[0]), .B(a[280]), .Z(n7877) );
  XOR U8590 ( .A(n7876), .B(n7877), .Z(n7879) );
  OR U8591 ( .A(n7839), .B(n7838), .Z(n7843) );
  NANDN U8592 ( .A(n7841), .B(n7840), .Z(n7842) );
  NAND U8593 ( .A(n7843), .B(n7842), .Z(n7878) );
  XNOR U8594 ( .A(n7879), .B(n7878), .Z(n7864) );
  NANDN U8595 ( .A(n7845), .B(n7844), .Z(n7849) );
  NAND U8596 ( .A(n7847), .B(n7846), .Z(n7848) );
  NAND U8597 ( .A(n7849), .B(n7848), .Z(n7865) );
  XNOR U8598 ( .A(n7864), .B(n7865), .Z(n7866) );
  NANDN U8599 ( .A(n7851), .B(n7850), .Z(n7855) );
  NAND U8600 ( .A(n7853), .B(n7852), .Z(n7854) );
  AND U8601 ( .A(n7855), .B(n7854), .Z(n7867) );
  XNOR U8602 ( .A(n7866), .B(n7867), .Z(n7863) );
  NAND U8603 ( .A(sreg[1299]), .B(n7856), .Z(n7860) );
  NANDN U8604 ( .A(n7858), .B(n7857), .Z(n7859) );
  AND U8605 ( .A(n7860), .B(n7859), .Z(n7862) );
  XNOR U8606 ( .A(n7862), .B(sreg[1300]), .Z(n7861) );
  XOR U8607 ( .A(n7863), .B(n7861), .Z(c[1300]) );
  NANDN U8608 ( .A(n7865), .B(n7864), .Z(n7869) );
  NAND U8609 ( .A(n7867), .B(n7866), .Z(n7868) );
  NAND U8610 ( .A(n7869), .B(n7868), .Z(n7885) );
  AND U8611 ( .A(b[2]), .B(a[279]), .Z(n7897) );
  AND U8612 ( .A(a[280]), .B(b[1]), .Z(n7895) );
  AND U8613 ( .A(a[278]), .B(b[3]), .Z(n7894) );
  XOR U8614 ( .A(n7895), .B(n7894), .Z(n7896) );
  XOR U8615 ( .A(n7897), .B(n7896), .Z(n7888) );
  NAND U8616 ( .A(b[0]), .B(a[281]), .Z(n7889) );
  XOR U8617 ( .A(n7888), .B(n7889), .Z(n7891) );
  OR U8618 ( .A(n7871), .B(n7870), .Z(n7875) );
  NANDN U8619 ( .A(n7873), .B(n7872), .Z(n7874) );
  NAND U8620 ( .A(n7875), .B(n7874), .Z(n7890) );
  XNOR U8621 ( .A(n7891), .B(n7890), .Z(n7882) );
  NANDN U8622 ( .A(n7877), .B(n7876), .Z(n7881) );
  OR U8623 ( .A(n7879), .B(n7878), .Z(n7880) );
  NAND U8624 ( .A(n7881), .B(n7880), .Z(n7883) );
  XNOR U8625 ( .A(n7882), .B(n7883), .Z(n7884) );
  XNOR U8626 ( .A(n7885), .B(n7884), .Z(n7900) );
  XNOR U8627 ( .A(n7900), .B(sreg[1301]), .Z(n7902) );
  XNOR U8628 ( .A(n7901), .B(n7902), .Z(c[1301]) );
  NANDN U8629 ( .A(n7883), .B(n7882), .Z(n7887) );
  NAND U8630 ( .A(n7885), .B(n7884), .Z(n7886) );
  NAND U8631 ( .A(n7887), .B(n7886), .Z(n7920) );
  NANDN U8632 ( .A(n7889), .B(n7888), .Z(n7893) );
  OR U8633 ( .A(n7891), .B(n7890), .Z(n7892) );
  NAND U8634 ( .A(n7893), .B(n7892), .Z(n7917) );
  AND U8635 ( .A(b[2]), .B(a[280]), .Z(n7908) );
  AND U8636 ( .A(a[281]), .B(b[1]), .Z(n7906) );
  AND U8637 ( .A(a[279]), .B(b[3]), .Z(n7905) );
  XOR U8638 ( .A(n7906), .B(n7905), .Z(n7907) );
  XOR U8639 ( .A(n7908), .B(n7907), .Z(n7911) );
  NAND U8640 ( .A(b[0]), .B(a[282]), .Z(n7912) );
  XNOR U8641 ( .A(n7911), .B(n7912), .Z(n7913) );
  OR U8642 ( .A(n7895), .B(n7894), .Z(n7899) );
  NANDN U8643 ( .A(n7897), .B(n7896), .Z(n7898) );
  AND U8644 ( .A(n7899), .B(n7898), .Z(n7914) );
  XNOR U8645 ( .A(n7913), .B(n7914), .Z(n7918) );
  XNOR U8646 ( .A(n7917), .B(n7918), .Z(n7919) );
  XNOR U8647 ( .A(n7920), .B(n7919), .Z(n7923) );
  XNOR U8648 ( .A(sreg[1302]), .B(n7923), .Z(n7925) );
  NAND U8649 ( .A(n7900), .B(sreg[1301]), .Z(n7904) );
  NANDN U8650 ( .A(n7902), .B(n7901), .Z(n7903) );
  AND U8651 ( .A(n7904), .B(n7903), .Z(n7924) );
  XOR U8652 ( .A(n7925), .B(n7924), .Z(c[1302]) );
  AND U8653 ( .A(b[2]), .B(a[281]), .Z(n7938) );
  AND U8654 ( .A(a[282]), .B(b[1]), .Z(n7936) );
  AND U8655 ( .A(a[280]), .B(b[3]), .Z(n7935) );
  XOR U8656 ( .A(n7936), .B(n7935), .Z(n7937) );
  XOR U8657 ( .A(n7938), .B(n7937), .Z(n7941) );
  NAND U8658 ( .A(b[0]), .B(a[283]), .Z(n7942) );
  XOR U8659 ( .A(n7941), .B(n7942), .Z(n7944) );
  OR U8660 ( .A(n7906), .B(n7905), .Z(n7910) );
  NANDN U8661 ( .A(n7908), .B(n7907), .Z(n7909) );
  NAND U8662 ( .A(n7910), .B(n7909), .Z(n7943) );
  XNOR U8663 ( .A(n7944), .B(n7943), .Z(n7929) );
  NANDN U8664 ( .A(n7912), .B(n7911), .Z(n7916) );
  NAND U8665 ( .A(n7914), .B(n7913), .Z(n7915) );
  NAND U8666 ( .A(n7916), .B(n7915), .Z(n7930) );
  XNOR U8667 ( .A(n7929), .B(n7930), .Z(n7931) );
  NANDN U8668 ( .A(n7918), .B(n7917), .Z(n7922) );
  NANDN U8669 ( .A(n7920), .B(n7919), .Z(n7921) );
  AND U8670 ( .A(n7922), .B(n7921), .Z(n7932) );
  XNOR U8671 ( .A(n7931), .B(n7932), .Z(n7948) );
  NAND U8672 ( .A(sreg[1302]), .B(n7923), .Z(n7927) );
  OR U8673 ( .A(n7925), .B(n7924), .Z(n7926) );
  AND U8674 ( .A(n7927), .B(n7926), .Z(n7947) );
  XNOR U8675 ( .A(n7947), .B(sreg[1303]), .Z(n7928) );
  XOR U8676 ( .A(n7948), .B(n7928), .Z(c[1303]) );
  NANDN U8677 ( .A(n7930), .B(n7929), .Z(n7934) );
  NAND U8678 ( .A(n7932), .B(n7931), .Z(n7933) );
  NAND U8679 ( .A(n7934), .B(n7933), .Z(n7953) );
  AND U8680 ( .A(b[2]), .B(a[282]), .Z(n7959) );
  AND U8681 ( .A(a[283]), .B(b[1]), .Z(n7957) );
  AND U8682 ( .A(a[281]), .B(b[3]), .Z(n7956) );
  XOR U8683 ( .A(n7957), .B(n7956), .Z(n7958) );
  XOR U8684 ( .A(n7959), .B(n7958), .Z(n7962) );
  NAND U8685 ( .A(b[0]), .B(a[284]), .Z(n7963) );
  XOR U8686 ( .A(n7962), .B(n7963), .Z(n7965) );
  OR U8687 ( .A(n7936), .B(n7935), .Z(n7940) );
  NANDN U8688 ( .A(n7938), .B(n7937), .Z(n7939) );
  NAND U8689 ( .A(n7940), .B(n7939), .Z(n7964) );
  XNOR U8690 ( .A(n7965), .B(n7964), .Z(n7950) );
  NANDN U8691 ( .A(n7942), .B(n7941), .Z(n7946) );
  OR U8692 ( .A(n7944), .B(n7943), .Z(n7945) );
  NAND U8693 ( .A(n7946), .B(n7945), .Z(n7951) );
  XNOR U8694 ( .A(n7950), .B(n7951), .Z(n7952) );
  XNOR U8695 ( .A(n7953), .B(n7952), .Z(n7969) );
  XOR U8696 ( .A(n7968), .B(sreg[1304]), .Z(n7949) );
  XOR U8697 ( .A(n7969), .B(n7949), .Z(c[1304]) );
  NANDN U8698 ( .A(n7951), .B(n7950), .Z(n7955) );
  NAND U8699 ( .A(n7953), .B(n7952), .Z(n7954) );
  NAND U8700 ( .A(n7955), .B(n7954), .Z(n7976) );
  AND U8701 ( .A(b[2]), .B(a[283]), .Z(n7982) );
  AND U8702 ( .A(a[284]), .B(b[1]), .Z(n7980) );
  AND U8703 ( .A(a[282]), .B(b[3]), .Z(n7979) );
  XOR U8704 ( .A(n7980), .B(n7979), .Z(n7981) );
  XOR U8705 ( .A(n7982), .B(n7981), .Z(n7985) );
  NAND U8706 ( .A(b[0]), .B(a[285]), .Z(n7986) );
  XOR U8707 ( .A(n7985), .B(n7986), .Z(n7988) );
  OR U8708 ( .A(n7957), .B(n7956), .Z(n7961) );
  NANDN U8709 ( .A(n7959), .B(n7958), .Z(n7960) );
  NAND U8710 ( .A(n7961), .B(n7960), .Z(n7987) );
  XNOR U8711 ( .A(n7988), .B(n7987), .Z(n7973) );
  NANDN U8712 ( .A(n7963), .B(n7962), .Z(n7967) );
  OR U8713 ( .A(n7965), .B(n7964), .Z(n7966) );
  NAND U8714 ( .A(n7967), .B(n7966), .Z(n7974) );
  XNOR U8715 ( .A(n7973), .B(n7974), .Z(n7975) );
  XNOR U8716 ( .A(n7976), .B(n7975), .Z(n7972) );
  XOR U8717 ( .A(n7971), .B(sreg[1305]), .Z(n7970) );
  XOR U8718 ( .A(n7972), .B(n7970), .Z(c[1305]) );
  NANDN U8719 ( .A(n7974), .B(n7973), .Z(n7978) );
  NAND U8720 ( .A(n7976), .B(n7975), .Z(n7977) );
  NAND U8721 ( .A(n7978), .B(n7977), .Z(n7994) );
  AND U8722 ( .A(b[2]), .B(a[284]), .Z(n8000) );
  AND U8723 ( .A(a[285]), .B(b[1]), .Z(n7998) );
  AND U8724 ( .A(a[283]), .B(b[3]), .Z(n7997) );
  XOR U8725 ( .A(n7998), .B(n7997), .Z(n7999) );
  XOR U8726 ( .A(n8000), .B(n7999), .Z(n8003) );
  NAND U8727 ( .A(b[0]), .B(a[286]), .Z(n8004) );
  XOR U8728 ( .A(n8003), .B(n8004), .Z(n8006) );
  OR U8729 ( .A(n7980), .B(n7979), .Z(n7984) );
  NANDN U8730 ( .A(n7982), .B(n7981), .Z(n7983) );
  NAND U8731 ( .A(n7984), .B(n7983), .Z(n8005) );
  XNOR U8732 ( .A(n8006), .B(n8005), .Z(n7991) );
  NANDN U8733 ( .A(n7986), .B(n7985), .Z(n7990) );
  OR U8734 ( .A(n7988), .B(n7987), .Z(n7989) );
  NAND U8735 ( .A(n7990), .B(n7989), .Z(n7992) );
  XNOR U8736 ( .A(n7991), .B(n7992), .Z(n7993) );
  XNOR U8737 ( .A(n7994), .B(n7993), .Z(n8009) );
  XNOR U8738 ( .A(n8009), .B(sreg[1306]), .Z(n8011) );
  XNOR U8739 ( .A(n8010), .B(n8011), .Z(c[1306]) );
  NANDN U8740 ( .A(n7992), .B(n7991), .Z(n7996) );
  NAND U8741 ( .A(n7994), .B(n7993), .Z(n7995) );
  NAND U8742 ( .A(n7996), .B(n7995), .Z(n8017) );
  AND U8743 ( .A(b[2]), .B(a[285]), .Z(n8023) );
  AND U8744 ( .A(a[286]), .B(b[1]), .Z(n8021) );
  AND U8745 ( .A(a[284]), .B(b[3]), .Z(n8020) );
  XOR U8746 ( .A(n8021), .B(n8020), .Z(n8022) );
  XOR U8747 ( .A(n8023), .B(n8022), .Z(n8026) );
  NAND U8748 ( .A(b[0]), .B(a[287]), .Z(n8027) );
  XOR U8749 ( .A(n8026), .B(n8027), .Z(n8029) );
  OR U8750 ( .A(n7998), .B(n7997), .Z(n8002) );
  NANDN U8751 ( .A(n8000), .B(n7999), .Z(n8001) );
  NAND U8752 ( .A(n8002), .B(n8001), .Z(n8028) );
  XNOR U8753 ( .A(n8029), .B(n8028), .Z(n8014) );
  NANDN U8754 ( .A(n8004), .B(n8003), .Z(n8008) );
  OR U8755 ( .A(n8006), .B(n8005), .Z(n8007) );
  NAND U8756 ( .A(n8008), .B(n8007), .Z(n8015) );
  XNOR U8757 ( .A(n8014), .B(n8015), .Z(n8016) );
  XNOR U8758 ( .A(n8017), .B(n8016), .Z(n8032) );
  XNOR U8759 ( .A(n8032), .B(sreg[1307]), .Z(n8034) );
  NAND U8760 ( .A(n8009), .B(sreg[1306]), .Z(n8013) );
  NANDN U8761 ( .A(n8011), .B(n8010), .Z(n8012) );
  AND U8762 ( .A(n8013), .B(n8012), .Z(n8033) );
  XOR U8763 ( .A(n8034), .B(n8033), .Z(c[1307]) );
  NANDN U8764 ( .A(n8015), .B(n8014), .Z(n8019) );
  NAND U8765 ( .A(n8017), .B(n8016), .Z(n8018) );
  NAND U8766 ( .A(n8019), .B(n8018), .Z(n8041) );
  AND U8767 ( .A(b[2]), .B(a[286]), .Z(n8053) );
  AND U8768 ( .A(a[287]), .B(b[1]), .Z(n8051) );
  AND U8769 ( .A(a[285]), .B(b[3]), .Z(n8050) );
  XOR U8770 ( .A(n8051), .B(n8050), .Z(n8052) );
  XOR U8771 ( .A(n8053), .B(n8052), .Z(n8044) );
  NAND U8772 ( .A(b[0]), .B(a[288]), .Z(n8045) );
  XOR U8773 ( .A(n8044), .B(n8045), .Z(n8047) );
  OR U8774 ( .A(n8021), .B(n8020), .Z(n8025) );
  NANDN U8775 ( .A(n8023), .B(n8022), .Z(n8024) );
  NAND U8776 ( .A(n8025), .B(n8024), .Z(n8046) );
  XNOR U8777 ( .A(n8047), .B(n8046), .Z(n8038) );
  NANDN U8778 ( .A(n8027), .B(n8026), .Z(n8031) );
  OR U8779 ( .A(n8029), .B(n8028), .Z(n8030) );
  NAND U8780 ( .A(n8031), .B(n8030), .Z(n8039) );
  XNOR U8781 ( .A(n8038), .B(n8039), .Z(n8040) );
  XOR U8782 ( .A(n8041), .B(n8040), .Z(n8058) );
  NAND U8783 ( .A(n8032), .B(sreg[1307]), .Z(n8036) );
  OR U8784 ( .A(n8034), .B(n8033), .Z(n8035) );
  NAND U8785 ( .A(n8036), .B(n8035), .Z(n8057) );
  XNOR U8786 ( .A(sreg[1308]), .B(n8057), .Z(n8037) );
  XOR U8787 ( .A(n8058), .B(n8037), .Z(c[1308]) );
  NANDN U8788 ( .A(n8039), .B(n8038), .Z(n8043) );
  NAND U8789 ( .A(n8041), .B(n8040), .Z(n8042) );
  NAND U8790 ( .A(n8043), .B(n8042), .Z(n8062) );
  NANDN U8791 ( .A(n8045), .B(n8044), .Z(n8049) );
  OR U8792 ( .A(n8047), .B(n8046), .Z(n8048) );
  AND U8793 ( .A(n8049), .B(n8048), .Z(n8061) );
  AND U8794 ( .A(b[2]), .B(a[287]), .Z(n8072) );
  AND U8795 ( .A(a[288]), .B(b[1]), .Z(n8070) );
  AND U8796 ( .A(a[286]), .B(b[3]), .Z(n8069) );
  XOR U8797 ( .A(n8070), .B(n8069), .Z(n8071) );
  XOR U8798 ( .A(n8072), .B(n8071), .Z(n8063) );
  NAND U8799 ( .A(b[0]), .B(a[289]), .Z(n8064) );
  XOR U8800 ( .A(n8063), .B(n8064), .Z(n8066) );
  OR U8801 ( .A(n8051), .B(n8050), .Z(n8055) );
  NANDN U8802 ( .A(n8053), .B(n8052), .Z(n8054) );
  NAND U8803 ( .A(n8055), .B(n8054), .Z(n8065) );
  XOR U8804 ( .A(n8066), .B(n8065), .Z(n8060) );
  XNOR U8805 ( .A(n8061), .B(n8060), .Z(n8056) );
  XNOR U8806 ( .A(n8062), .B(n8056), .Z(n8077) );
  XOR U8807 ( .A(n8076), .B(sreg[1309]), .Z(n8059) );
  XOR U8808 ( .A(n8077), .B(n8059), .Z(c[1309]) );
  NANDN U8809 ( .A(n8064), .B(n8063), .Z(n8068) );
  OR U8810 ( .A(n8066), .B(n8065), .Z(n8067) );
  AND U8811 ( .A(n8068), .B(n8067), .Z(n8082) );
  AND U8812 ( .A(b[2]), .B(a[288]), .Z(n8087) );
  AND U8813 ( .A(a[289]), .B(b[1]), .Z(n8085) );
  AND U8814 ( .A(a[287]), .B(b[3]), .Z(n8084) );
  XOR U8815 ( .A(n8085), .B(n8084), .Z(n8086) );
  XOR U8816 ( .A(n8087), .B(n8086), .Z(n8090) );
  NAND U8817 ( .A(b[0]), .B(a[290]), .Z(n8091) );
  XOR U8818 ( .A(n8090), .B(n8091), .Z(n8093) );
  OR U8819 ( .A(n8070), .B(n8069), .Z(n8074) );
  NANDN U8820 ( .A(n8072), .B(n8071), .Z(n8073) );
  NAND U8821 ( .A(n8074), .B(n8073), .Z(n8092) );
  XOR U8822 ( .A(n8093), .B(n8092), .Z(n8081) );
  XNOR U8823 ( .A(n8082), .B(n8081), .Z(n8075) );
  XOR U8824 ( .A(n8083), .B(n8075), .Z(n8080) );
  XOR U8825 ( .A(sreg[1310]), .B(n8079), .Z(n8078) );
  XNOR U8826 ( .A(n8080), .B(n8078), .Z(c[1310]) );
  AND U8827 ( .A(b[2]), .B(a[289]), .Z(n8110) );
  AND U8828 ( .A(a[290]), .B(b[1]), .Z(n8108) );
  AND U8829 ( .A(a[288]), .B(b[3]), .Z(n8107) );
  XOR U8830 ( .A(n8108), .B(n8107), .Z(n8109) );
  XOR U8831 ( .A(n8110), .B(n8109), .Z(n8113) );
  NAND U8832 ( .A(b[0]), .B(a[291]), .Z(n8114) );
  XOR U8833 ( .A(n8113), .B(n8114), .Z(n8116) );
  OR U8834 ( .A(n8085), .B(n8084), .Z(n8089) );
  NANDN U8835 ( .A(n8087), .B(n8086), .Z(n8088) );
  NAND U8836 ( .A(n8089), .B(n8088), .Z(n8115) );
  XNOR U8837 ( .A(n8116), .B(n8115), .Z(n8101) );
  NANDN U8838 ( .A(n8091), .B(n8090), .Z(n8095) );
  OR U8839 ( .A(n8093), .B(n8092), .Z(n8094) );
  NAND U8840 ( .A(n8095), .B(n8094), .Z(n8102) );
  XNOR U8841 ( .A(n8101), .B(n8102), .Z(n8103) );
  XOR U8842 ( .A(n8104), .B(n8103), .Z(n8096) );
  XNOR U8843 ( .A(n8096), .B(sreg[1311]), .Z(n8097) );
  XOR U8844 ( .A(n8098), .B(n8097), .Z(c[1311]) );
  NAND U8845 ( .A(n8096), .B(sreg[1311]), .Z(n8100) );
  OR U8846 ( .A(n8098), .B(n8097), .Z(n8099) );
  NAND U8847 ( .A(n8100), .B(n8099), .Z(n8121) );
  NANDN U8848 ( .A(n8102), .B(n8101), .Z(n8106) );
  NANDN U8849 ( .A(n8104), .B(n8103), .Z(n8105) );
  AND U8850 ( .A(n8106), .B(n8105), .Z(n8125) );
  AND U8851 ( .A(b[2]), .B(a[290]), .Z(n8133) );
  AND U8852 ( .A(a[291]), .B(b[1]), .Z(n8131) );
  AND U8853 ( .A(a[289]), .B(b[3]), .Z(n8130) );
  XOR U8854 ( .A(n8131), .B(n8130), .Z(n8132) );
  XOR U8855 ( .A(n8133), .B(n8132), .Z(n8126) );
  NAND U8856 ( .A(b[0]), .B(a[292]), .Z(n8127) );
  XOR U8857 ( .A(n8126), .B(n8127), .Z(n8128) );
  OR U8858 ( .A(n8108), .B(n8107), .Z(n8112) );
  NANDN U8859 ( .A(n8110), .B(n8109), .Z(n8111) );
  AND U8860 ( .A(n8112), .B(n8111), .Z(n8129) );
  XOR U8861 ( .A(n8128), .B(n8129), .Z(n8123) );
  NANDN U8862 ( .A(n8114), .B(n8113), .Z(n8118) );
  OR U8863 ( .A(n8116), .B(n8115), .Z(n8117) );
  AND U8864 ( .A(n8118), .B(n8117), .Z(n8124) );
  XOR U8865 ( .A(n8123), .B(n8124), .Z(n8119) );
  XNOR U8866 ( .A(n8125), .B(n8119), .Z(n8122) );
  XOR U8867 ( .A(sreg[1312]), .B(n8122), .Z(n8120) );
  XNOR U8868 ( .A(n8121), .B(n8120), .Z(c[1312]) );
  AND U8869 ( .A(b[2]), .B(a[291]), .Z(n8139) );
  AND U8870 ( .A(a[292]), .B(b[1]), .Z(n8137) );
  AND U8871 ( .A(a[290]), .B(b[3]), .Z(n8136) );
  XOR U8872 ( .A(n8137), .B(n8136), .Z(n8138) );
  XOR U8873 ( .A(n8139), .B(n8138), .Z(n8142) );
  NAND U8874 ( .A(b[0]), .B(a[293]), .Z(n8143) );
  XNOR U8875 ( .A(n8142), .B(n8143), .Z(n8144) );
  OR U8876 ( .A(n8131), .B(n8130), .Z(n8135) );
  NANDN U8877 ( .A(n8133), .B(n8132), .Z(n8134) );
  AND U8878 ( .A(n8135), .B(n8134), .Z(n8145) );
  XNOR U8879 ( .A(n8144), .B(n8145), .Z(n8149) );
  XNOR U8880 ( .A(n8148), .B(n8149), .Z(n8150) );
  XNOR U8881 ( .A(n8151), .B(n8150), .Z(n8154) );
  XNOR U8882 ( .A(sreg[1313]), .B(n8154), .Z(n8155) );
  XOR U8883 ( .A(n8156), .B(n8155), .Z(c[1313]) );
  AND U8884 ( .A(b[2]), .B(a[292]), .Z(n8169) );
  AND U8885 ( .A(a[293]), .B(b[1]), .Z(n8167) );
  AND U8886 ( .A(a[291]), .B(b[3]), .Z(n8166) );
  XOR U8887 ( .A(n8167), .B(n8166), .Z(n8168) );
  XOR U8888 ( .A(n8169), .B(n8168), .Z(n8172) );
  NAND U8889 ( .A(b[0]), .B(a[294]), .Z(n8173) );
  XOR U8890 ( .A(n8172), .B(n8173), .Z(n8175) );
  OR U8891 ( .A(n8137), .B(n8136), .Z(n8141) );
  NANDN U8892 ( .A(n8139), .B(n8138), .Z(n8140) );
  NAND U8893 ( .A(n8141), .B(n8140), .Z(n8174) );
  XNOR U8894 ( .A(n8175), .B(n8174), .Z(n8160) );
  NANDN U8895 ( .A(n8143), .B(n8142), .Z(n8147) );
  NAND U8896 ( .A(n8145), .B(n8144), .Z(n8146) );
  NAND U8897 ( .A(n8147), .B(n8146), .Z(n8161) );
  XNOR U8898 ( .A(n8160), .B(n8161), .Z(n8162) );
  NANDN U8899 ( .A(n8149), .B(n8148), .Z(n8153) );
  NANDN U8900 ( .A(n8151), .B(n8150), .Z(n8152) );
  NAND U8901 ( .A(n8153), .B(n8152), .Z(n8163) );
  XOR U8902 ( .A(n8162), .B(n8163), .Z(n8179) );
  NAND U8903 ( .A(sreg[1313]), .B(n8154), .Z(n8158) );
  OR U8904 ( .A(n8156), .B(n8155), .Z(n8157) );
  NAND U8905 ( .A(n8158), .B(n8157), .Z(n8178) );
  XNOR U8906 ( .A(sreg[1314]), .B(n8178), .Z(n8159) );
  XNOR U8907 ( .A(n8179), .B(n8159), .Z(c[1314]) );
  NANDN U8908 ( .A(n8161), .B(n8160), .Z(n8165) );
  NANDN U8909 ( .A(n8163), .B(n8162), .Z(n8164) );
  NAND U8910 ( .A(n8165), .B(n8164), .Z(n8196) );
  AND U8911 ( .A(b[2]), .B(a[293]), .Z(n8190) );
  AND U8912 ( .A(a[294]), .B(b[1]), .Z(n8188) );
  AND U8913 ( .A(a[292]), .B(b[3]), .Z(n8187) );
  XOR U8914 ( .A(n8188), .B(n8187), .Z(n8189) );
  XOR U8915 ( .A(n8190), .B(n8189), .Z(n8181) );
  NAND U8916 ( .A(b[0]), .B(a[295]), .Z(n8182) );
  XOR U8917 ( .A(n8181), .B(n8182), .Z(n8184) );
  OR U8918 ( .A(n8167), .B(n8166), .Z(n8171) );
  NANDN U8919 ( .A(n8169), .B(n8168), .Z(n8170) );
  NAND U8920 ( .A(n8171), .B(n8170), .Z(n8183) );
  XNOR U8921 ( .A(n8184), .B(n8183), .Z(n8193) );
  NANDN U8922 ( .A(n8173), .B(n8172), .Z(n8177) );
  OR U8923 ( .A(n8175), .B(n8174), .Z(n8176) );
  NAND U8924 ( .A(n8177), .B(n8176), .Z(n8194) );
  XNOR U8925 ( .A(n8193), .B(n8194), .Z(n8195) );
  XOR U8926 ( .A(n8196), .B(n8195), .Z(n8200) );
  XNOR U8927 ( .A(sreg[1315]), .B(n8199), .Z(n8180) );
  XOR U8928 ( .A(n8200), .B(n8180), .Z(c[1315]) );
  NANDN U8929 ( .A(n8182), .B(n8181), .Z(n8186) );
  OR U8930 ( .A(n8184), .B(n8183), .Z(n8185) );
  NAND U8931 ( .A(n8186), .B(n8185), .Z(n8214) );
  AND U8932 ( .A(b[2]), .B(a[294]), .Z(n8205) );
  AND U8933 ( .A(a[295]), .B(b[1]), .Z(n8203) );
  AND U8934 ( .A(a[293]), .B(b[3]), .Z(n8202) );
  XOR U8935 ( .A(n8203), .B(n8202), .Z(n8204) );
  XOR U8936 ( .A(n8205), .B(n8204), .Z(n8208) );
  NAND U8937 ( .A(b[0]), .B(a[296]), .Z(n8209) );
  XNOR U8938 ( .A(n8208), .B(n8209), .Z(n8210) );
  OR U8939 ( .A(n8188), .B(n8187), .Z(n8192) );
  NANDN U8940 ( .A(n8190), .B(n8189), .Z(n8191) );
  AND U8941 ( .A(n8192), .B(n8191), .Z(n8211) );
  XNOR U8942 ( .A(n8210), .B(n8211), .Z(n8215) );
  XNOR U8943 ( .A(n8214), .B(n8215), .Z(n8216) );
  NANDN U8944 ( .A(n8194), .B(n8193), .Z(n8198) );
  NAND U8945 ( .A(n8196), .B(n8195), .Z(n8197) );
  NAND U8946 ( .A(n8198), .B(n8197), .Z(n8217) );
  XOR U8947 ( .A(n8216), .B(n8217), .Z(n8221) );
  XOR U8948 ( .A(n8220), .B(sreg[1316]), .Z(n8201) );
  XNOR U8949 ( .A(n8221), .B(n8201), .Z(c[1316]) );
  AND U8950 ( .A(b[2]), .B(a[295]), .Z(n8232) );
  AND U8951 ( .A(a[296]), .B(b[1]), .Z(n8230) );
  AND U8952 ( .A(a[294]), .B(b[3]), .Z(n8229) );
  XOR U8953 ( .A(n8230), .B(n8229), .Z(n8231) );
  XOR U8954 ( .A(n8232), .B(n8231), .Z(n8235) );
  NAND U8955 ( .A(b[0]), .B(a[297]), .Z(n8236) );
  XOR U8956 ( .A(n8235), .B(n8236), .Z(n8238) );
  OR U8957 ( .A(n8203), .B(n8202), .Z(n8207) );
  NANDN U8958 ( .A(n8205), .B(n8204), .Z(n8206) );
  NAND U8959 ( .A(n8207), .B(n8206), .Z(n8237) );
  XNOR U8960 ( .A(n8238), .B(n8237), .Z(n8223) );
  NANDN U8961 ( .A(n8209), .B(n8208), .Z(n8213) );
  NAND U8962 ( .A(n8211), .B(n8210), .Z(n8212) );
  NAND U8963 ( .A(n8213), .B(n8212), .Z(n8224) );
  XNOR U8964 ( .A(n8223), .B(n8224), .Z(n8225) );
  NANDN U8965 ( .A(n8215), .B(n8214), .Z(n8219) );
  NANDN U8966 ( .A(n8217), .B(n8216), .Z(n8218) );
  AND U8967 ( .A(n8219), .B(n8218), .Z(n8226) );
  XNOR U8968 ( .A(n8225), .B(n8226), .Z(n8242) );
  XOR U8969 ( .A(n8241), .B(sreg[1317]), .Z(n8222) );
  XOR U8970 ( .A(n8242), .B(n8222), .Z(c[1317]) );
  NANDN U8971 ( .A(n8224), .B(n8223), .Z(n8228) );
  NAND U8972 ( .A(n8226), .B(n8225), .Z(n8227) );
  NAND U8973 ( .A(n8228), .B(n8227), .Z(n8261) );
  AND U8974 ( .A(b[2]), .B(a[296]), .Z(n8255) );
  AND U8975 ( .A(a[297]), .B(b[1]), .Z(n8253) );
  AND U8976 ( .A(a[295]), .B(b[3]), .Z(n8252) );
  XOR U8977 ( .A(n8253), .B(n8252), .Z(n8254) );
  XOR U8978 ( .A(n8255), .B(n8254), .Z(n8246) );
  NAND U8979 ( .A(b[0]), .B(a[298]), .Z(n8247) );
  XOR U8980 ( .A(n8246), .B(n8247), .Z(n8249) );
  OR U8981 ( .A(n8230), .B(n8229), .Z(n8234) );
  NANDN U8982 ( .A(n8232), .B(n8231), .Z(n8233) );
  NAND U8983 ( .A(n8234), .B(n8233), .Z(n8248) );
  XNOR U8984 ( .A(n8249), .B(n8248), .Z(n8258) );
  NANDN U8985 ( .A(n8236), .B(n8235), .Z(n8240) );
  OR U8986 ( .A(n8238), .B(n8237), .Z(n8239) );
  NAND U8987 ( .A(n8240), .B(n8239), .Z(n8259) );
  XNOR U8988 ( .A(n8258), .B(n8259), .Z(n8260) );
  XNOR U8989 ( .A(n8261), .B(n8260), .Z(n8245) );
  XOR U8990 ( .A(n8244), .B(sreg[1318]), .Z(n8243) );
  XOR U8991 ( .A(n8245), .B(n8243), .Z(c[1318]) );
  NANDN U8992 ( .A(n8247), .B(n8246), .Z(n8251) );
  OR U8993 ( .A(n8249), .B(n8248), .Z(n8250) );
  NAND U8994 ( .A(n8251), .B(n8250), .Z(n8276) );
  AND U8995 ( .A(b[2]), .B(a[297]), .Z(n8267) );
  AND U8996 ( .A(a[298]), .B(b[1]), .Z(n8265) );
  AND U8997 ( .A(a[296]), .B(b[3]), .Z(n8264) );
  XOR U8998 ( .A(n8265), .B(n8264), .Z(n8266) );
  XOR U8999 ( .A(n8267), .B(n8266), .Z(n8270) );
  NAND U9000 ( .A(b[0]), .B(a[299]), .Z(n8271) );
  XNOR U9001 ( .A(n8270), .B(n8271), .Z(n8272) );
  OR U9002 ( .A(n8253), .B(n8252), .Z(n8257) );
  NANDN U9003 ( .A(n8255), .B(n8254), .Z(n8256) );
  AND U9004 ( .A(n8257), .B(n8256), .Z(n8273) );
  XNOR U9005 ( .A(n8272), .B(n8273), .Z(n8277) );
  XNOR U9006 ( .A(n8276), .B(n8277), .Z(n8278) );
  NANDN U9007 ( .A(n8259), .B(n8258), .Z(n8263) );
  NAND U9008 ( .A(n8261), .B(n8260), .Z(n8262) );
  AND U9009 ( .A(n8263), .B(n8262), .Z(n8279) );
  XOR U9010 ( .A(n8278), .B(n8279), .Z(n8282) );
  XNOR U9011 ( .A(sreg[1319]), .B(n8282), .Z(n8284) );
  XNOR U9012 ( .A(n8283), .B(n8284), .Z(c[1319]) );
  AND U9013 ( .A(b[2]), .B(a[298]), .Z(n8297) );
  AND U9014 ( .A(a[299]), .B(b[1]), .Z(n8295) );
  AND U9015 ( .A(a[297]), .B(b[3]), .Z(n8294) );
  XOR U9016 ( .A(n8295), .B(n8294), .Z(n8296) );
  XOR U9017 ( .A(n8297), .B(n8296), .Z(n8300) );
  NAND U9018 ( .A(b[0]), .B(a[300]), .Z(n8301) );
  XOR U9019 ( .A(n8300), .B(n8301), .Z(n8303) );
  OR U9020 ( .A(n8265), .B(n8264), .Z(n8269) );
  NANDN U9021 ( .A(n8267), .B(n8266), .Z(n8268) );
  NAND U9022 ( .A(n8269), .B(n8268), .Z(n8302) );
  XNOR U9023 ( .A(n8303), .B(n8302), .Z(n8288) );
  NANDN U9024 ( .A(n8271), .B(n8270), .Z(n8275) );
  NAND U9025 ( .A(n8273), .B(n8272), .Z(n8274) );
  NAND U9026 ( .A(n8275), .B(n8274), .Z(n8289) );
  XNOR U9027 ( .A(n8288), .B(n8289), .Z(n8290) );
  NANDN U9028 ( .A(n8277), .B(n8276), .Z(n8281) );
  NAND U9029 ( .A(n8279), .B(n8278), .Z(n8280) );
  NAND U9030 ( .A(n8281), .B(n8280), .Z(n8291) );
  XOR U9031 ( .A(n8290), .B(n8291), .Z(n8307) );
  NAND U9032 ( .A(sreg[1319]), .B(n8282), .Z(n8286) );
  NANDN U9033 ( .A(n8284), .B(n8283), .Z(n8285) );
  NAND U9034 ( .A(n8286), .B(n8285), .Z(n8306) );
  XNOR U9035 ( .A(sreg[1320]), .B(n8306), .Z(n8287) );
  XNOR U9036 ( .A(n8307), .B(n8287), .Z(c[1320]) );
  NANDN U9037 ( .A(n8289), .B(n8288), .Z(n8293) );
  NANDN U9038 ( .A(n8291), .B(n8290), .Z(n8292) );
  NAND U9039 ( .A(n8293), .B(n8292), .Z(n8326) );
  AND U9040 ( .A(b[2]), .B(a[299]), .Z(n8320) );
  AND U9041 ( .A(a[300]), .B(b[1]), .Z(n8318) );
  AND U9042 ( .A(a[298]), .B(b[3]), .Z(n8317) );
  XOR U9043 ( .A(n8318), .B(n8317), .Z(n8319) );
  XOR U9044 ( .A(n8320), .B(n8319), .Z(n8311) );
  NAND U9045 ( .A(b[0]), .B(a[301]), .Z(n8312) );
  XOR U9046 ( .A(n8311), .B(n8312), .Z(n8314) );
  OR U9047 ( .A(n8295), .B(n8294), .Z(n8299) );
  NANDN U9048 ( .A(n8297), .B(n8296), .Z(n8298) );
  NAND U9049 ( .A(n8299), .B(n8298), .Z(n8313) );
  XNOR U9050 ( .A(n8314), .B(n8313), .Z(n8323) );
  NANDN U9051 ( .A(n8301), .B(n8300), .Z(n8305) );
  OR U9052 ( .A(n8303), .B(n8302), .Z(n8304) );
  NAND U9053 ( .A(n8305), .B(n8304), .Z(n8324) );
  XNOR U9054 ( .A(n8323), .B(n8324), .Z(n8325) );
  XOR U9055 ( .A(n8326), .B(n8325), .Z(n8310) );
  XNOR U9056 ( .A(sreg[1321]), .B(n8309), .Z(n8308) );
  XOR U9057 ( .A(n8310), .B(n8308), .Z(c[1321]) );
  NANDN U9058 ( .A(n8312), .B(n8311), .Z(n8316) );
  OR U9059 ( .A(n8314), .B(n8313), .Z(n8315) );
  NAND U9060 ( .A(n8316), .B(n8315), .Z(n8341) );
  AND U9061 ( .A(b[2]), .B(a[300]), .Z(n8332) );
  AND U9062 ( .A(a[301]), .B(b[1]), .Z(n8330) );
  AND U9063 ( .A(a[299]), .B(b[3]), .Z(n8329) );
  XOR U9064 ( .A(n8330), .B(n8329), .Z(n8331) );
  XOR U9065 ( .A(n8332), .B(n8331), .Z(n8335) );
  NAND U9066 ( .A(b[0]), .B(a[302]), .Z(n8336) );
  XNOR U9067 ( .A(n8335), .B(n8336), .Z(n8337) );
  OR U9068 ( .A(n8318), .B(n8317), .Z(n8322) );
  NANDN U9069 ( .A(n8320), .B(n8319), .Z(n8321) );
  AND U9070 ( .A(n8322), .B(n8321), .Z(n8338) );
  XNOR U9071 ( .A(n8337), .B(n8338), .Z(n8342) );
  XNOR U9072 ( .A(n8341), .B(n8342), .Z(n8343) );
  NANDN U9073 ( .A(n8324), .B(n8323), .Z(n8328) );
  NAND U9074 ( .A(n8326), .B(n8325), .Z(n8327) );
  AND U9075 ( .A(n8328), .B(n8327), .Z(n8344) );
  XOR U9076 ( .A(n8343), .B(n8344), .Z(n8347) );
  XNOR U9077 ( .A(sreg[1322]), .B(n8347), .Z(n8348) );
  XOR U9078 ( .A(n8349), .B(n8348), .Z(c[1322]) );
  AND U9079 ( .A(b[2]), .B(a[301]), .Z(n8364) );
  AND U9080 ( .A(a[302]), .B(b[1]), .Z(n8362) );
  AND U9081 ( .A(a[300]), .B(b[3]), .Z(n8361) );
  XOR U9082 ( .A(n8362), .B(n8361), .Z(n8363) );
  XOR U9083 ( .A(n8364), .B(n8363), .Z(n8367) );
  NAND U9084 ( .A(b[0]), .B(a[303]), .Z(n8368) );
  XOR U9085 ( .A(n8367), .B(n8368), .Z(n8370) );
  OR U9086 ( .A(n8330), .B(n8329), .Z(n8334) );
  NANDN U9087 ( .A(n8332), .B(n8331), .Z(n8333) );
  NAND U9088 ( .A(n8334), .B(n8333), .Z(n8369) );
  XNOR U9089 ( .A(n8370), .B(n8369), .Z(n8355) );
  NANDN U9090 ( .A(n8336), .B(n8335), .Z(n8340) );
  NAND U9091 ( .A(n8338), .B(n8337), .Z(n8339) );
  NAND U9092 ( .A(n8340), .B(n8339), .Z(n8356) );
  XNOR U9093 ( .A(n8355), .B(n8356), .Z(n8357) );
  NANDN U9094 ( .A(n8342), .B(n8341), .Z(n8346) );
  NAND U9095 ( .A(n8344), .B(n8343), .Z(n8345) );
  NAND U9096 ( .A(n8346), .B(n8345), .Z(n8358) );
  XOR U9097 ( .A(n8357), .B(n8358), .Z(n8354) );
  NAND U9098 ( .A(sreg[1322]), .B(n8347), .Z(n8351) );
  OR U9099 ( .A(n8349), .B(n8348), .Z(n8350) );
  NAND U9100 ( .A(n8351), .B(n8350), .Z(n8353) );
  XNOR U9101 ( .A(sreg[1323]), .B(n8353), .Z(n8352) );
  XNOR U9102 ( .A(n8354), .B(n8352), .Z(c[1323]) );
  NANDN U9103 ( .A(n8356), .B(n8355), .Z(n8360) );
  NANDN U9104 ( .A(n8358), .B(n8357), .Z(n8359) );
  NAND U9105 ( .A(n8360), .B(n8359), .Z(n8381) );
  AND U9106 ( .A(b[2]), .B(a[302]), .Z(n8387) );
  AND U9107 ( .A(a[303]), .B(b[1]), .Z(n8385) );
  AND U9108 ( .A(a[301]), .B(b[3]), .Z(n8384) );
  XOR U9109 ( .A(n8385), .B(n8384), .Z(n8386) );
  XOR U9110 ( .A(n8387), .B(n8386), .Z(n8390) );
  NAND U9111 ( .A(b[0]), .B(a[304]), .Z(n8391) );
  XOR U9112 ( .A(n8390), .B(n8391), .Z(n8393) );
  OR U9113 ( .A(n8362), .B(n8361), .Z(n8366) );
  NANDN U9114 ( .A(n8364), .B(n8363), .Z(n8365) );
  NAND U9115 ( .A(n8366), .B(n8365), .Z(n8392) );
  XNOR U9116 ( .A(n8393), .B(n8392), .Z(n8378) );
  NANDN U9117 ( .A(n8368), .B(n8367), .Z(n8372) );
  OR U9118 ( .A(n8370), .B(n8369), .Z(n8371) );
  NAND U9119 ( .A(n8372), .B(n8371), .Z(n8379) );
  XNOR U9120 ( .A(n8378), .B(n8379), .Z(n8380) );
  XNOR U9121 ( .A(n8381), .B(n8380), .Z(n8373) );
  XOR U9122 ( .A(sreg[1324]), .B(n8373), .Z(n8375) );
  XNOR U9123 ( .A(n8374), .B(n8375), .Z(c[1324]) );
  OR U9124 ( .A(n8373), .B(sreg[1324]), .Z(n8377) );
  NAND U9125 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U9126 ( .A(n8377), .B(n8376), .Z(n8416) );
  NANDN U9127 ( .A(n8379), .B(n8378), .Z(n8383) );
  NAND U9128 ( .A(n8381), .B(n8380), .Z(n8382) );
  NAND U9129 ( .A(n8383), .B(n8382), .Z(n8400) );
  AND U9130 ( .A(b[2]), .B(a[303]), .Z(n8412) );
  AND U9131 ( .A(a[304]), .B(b[1]), .Z(n8410) );
  AND U9132 ( .A(a[302]), .B(b[3]), .Z(n8409) );
  XOR U9133 ( .A(n8410), .B(n8409), .Z(n8411) );
  XOR U9134 ( .A(n8412), .B(n8411), .Z(n8403) );
  NAND U9135 ( .A(b[0]), .B(a[305]), .Z(n8404) );
  XOR U9136 ( .A(n8403), .B(n8404), .Z(n8406) );
  OR U9137 ( .A(n8385), .B(n8384), .Z(n8389) );
  NANDN U9138 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U9139 ( .A(n8389), .B(n8388), .Z(n8405) );
  XNOR U9140 ( .A(n8406), .B(n8405), .Z(n8397) );
  NANDN U9141 ( .A(n8391), .B(n8390), .Z(n8395) );
  OR U9142 ( .A(n8393), .B(n8392), .Z(n8394) );
  NAND U9143 ( .A(n8395), .B(n8394), .Z(n8398) );
  XNOR U9144 ( .A(n8397), .B(n8398), .Z(n8399) );
  XNOR U9145 ( .A(n8400), .B(n8399), .Z(n8417) );
  XOR U9146 ( .A(sreg[1325]), .B(n8417), .Z(n8396) );
  XOR U9147 ( .A(n8416), .B(n8396), .Z(c[1325]) );
  NANDN U9148 ( .A(n8398), .B(n8397), .Z(n8402) );
  NAND U9149 ( .A(n8400), .B(n8399), .Z(n8401) );
  NAND U9150 ( .A(n8402), .B(n8401), .Z(n8421) );
  NANDN U9151 ( .A(n8404), .B(n8403), .Z(n8408) );
  OR U9152 ( .A(n8406), .B(n8405), .Z(n8407) );
  AND U9153 ( .A(n8408), .B(n8407), .Z(n8420) );
  AND U9154 ( .A(b[2]), .B(a[304]), .Z(n8425) );
  AND U9155 ( .A(a[305]), .B(b[1]), .Z(n8423) );
  AND U9156 ( .A(a[303]), .B(b[3]), .Z(n8422) );
  XOR U9157 ( .A(n8423), .B(n8422), .Z(n8424) );
  XOR U9158 ( .A(n8425), .B(n8424), .Z(n8428) );
  NAND U9159 ( .A(b[0]), .B(a[306]), .Z(n8429) );
  XOR U9160 ( .A(n8428), .B(n8429), .Z(n8431) );
  OR U9161 ( .A(n8410), .B(n8409), .Z(n8414) );
  NANDN U9162 ( .A(n8412), .B(n8411), .Z(n8413) );
  NAND U9163 ( .A(n8414), .B(n8413), .Z(n8430) );
  XOR U9164 ( .A(n8431), .B(n8430), .Z(n8419) );
  XNOR U9165 ( .A(n8420), .B(n8419), .Z(n8415) );
  XNOR U9166 ( .A(n8421), .B(n8415), .Z(n8435) );
  XOR U9167 ( .A(n8434), .B(sreg[1326]), .Z(n8418) );
  XOR U9168 ( .A(n8435), .B(n8418), .Z(c[1326]) );
  AND U9169 ( .A(b[2]), .B(a[305]), .Z(n8448) );
  AND U9170 ( .A(a[306]), .B(b[1]), .Z(n8446) );
  AND U9171 ( .A(a[304]), .B(b[3]), .Z(n8445) );
  XOR U9172 ( .A(n8446), .B(n8445), .Z(n8447) );
  XOR U9173 ( .A(n8448), .B(n8447), .Z(n8451) );
  NAND U9174 ( .A(b[0]), .B(a[307]), .Z(n8452) );
  XOR U9175 ( .A(n8451), .B(n8452), .Z(n8454) );
  OR U9176 ( .A(n8423), .B(n8422), .Z(n8427) );
  NANDN U9177 ( .A(n8425), .B(n8424), .Z(n8426) );
  NAND U9178 ( .A(n8427), .B(n8426), .Z(n8453) );
  XNOR U9179 ( .A(n8454), .B(n8453), .Z(n8439) );
  NANDN U9180 ( .A(n8429), .B(n8428), .Z(n8433) );
  OR U9181 ( .A(n8431), .B(n8430), .Z(n8432) );
  NAND U9182 ( .A(n8433), .B(n8432), .Z(n8440) );
  XNOR U9183 ( .A(n8439), .B(n8440), .Z(n8441) );
  XNOR U9184 ( .A(n8442), .B(n8441), .Z(n8438) );
  XOR U9185 ( .A(n8437), .B(sreg[1327]), .Z(n8436) );
  XNOR U9186 ( .A(n8438), .B(n8436), .Z(c[1327]) );
  NANDN U9187 ( .A(n8440), .B(n8439), .Z(n8444) );
  NANDN U9188 ( .A(n8442), .B(n8441), .Z(n8443) );
  NAND U9189 ( .A(n8444), .B(n8443), .Z(n8460) );
  AND U9190 ( .A(b[2]), .B(a[306]), .Z(n8466) );
  AND U9191 ( .A(a[307]), .B(b[1]), .Z(n8464) );
  AND U9192 ( .A(a[305]), .B(b[3]), .Z(n8463) );
  XOR U9193 ( .A(n8464), .B(n8463), .Z(n8465) );
  XOR U9194 ( .A(n8466), .B(n8465), .Z(n8469) );
  NAND U9195 ( .A(b[0]), .B(a[308]), .Z(n8470) );
  XOR U9196 ( .A(n8469), .B(n8470), .Z(n8472) );
  OR U9197 ( .A(n8446), .B(n8445), .Z(n8450) );
  NANDN U9198 ( .A(n8448), .B(n8447), .Z(n8449) );
  NAND U9199 ( .A(n8450), .B(n8449), .Z(n8471) );
  XNOR U9200 ( .A(n8472), .B(n8471), .Z(n8457) );
  NANDN U9201 ( .A(n8452), .B(n8451), .Z(n8456) );
  OR U9202 ( .A(n8454), .B(n8453), .Z(n8455) );
  NAND U9203 ( .A(n8456), .B(n8455), .Z(n8458) );
  XNOR U9204 ( .A(n8457), .B(n8458), .Z(n8459) );
  XNOR U9205 ( .A(n8460), .B(n8459), .Z(n8476) );
  XNOR U9206 ( .A(n8476), .B(sreg[1328]), .Z(n8478) );
  XNOR U9207 ( .A(n8477), .B(n8478), .Z(c[1328]) );
  NANDN U9208 ( .A(n8458), .B(n8457), .Z(n8462) );
  NAND U9209 ( .A(n8460), .B(n8459), .Z(n8461) );
  NAND U9210 ( .A(n8462), .B(n8461), .Z(n8483) );
  AND U9211 ( .A(b[2]), .B(a[307]), .Z(n8487) );
  AND U9212 ( .A(a[308]), .B(b[1]), .Z(n8485) );
  AND U9213 ( .A(a[306]), .B(b[3]), .Z(n8484) );
  XOR U9214 ( .A(n8485), .B(n8484), .Z(n8486) );
  XOR U9215 ( .A(n8487), .B(n8486), .Z(n8490) );
  NAND U9216 ( .A(b[0]), .B(a[309]), .Z(n8491) );
  XOR U9217 ( .A(n8490), .B(n8491), .Z(n8492) );
  OR U9218 ( .A(n8464), .B(n8463), .Z(n8468) );
  NANDN U9219 ( .A(n8466), .B(n8465), .Z(n8467) );
  AND U9220 ( .A(n8468), .B(n8467), .Z(n8493) );
  XOR U9221 ( .A(n8492), .B(n8493), .Z(n8481) );
  NANDN U9222 ( .A(n8470), .B(n8469), .Z(n8474) );
  OR U9223 ( .A(n8472), .B(n8471), .Z(n8473) );
  AND U9224 ( .A(n8474), .B(n8473), .Z(n8482) );
  XOR U9225 ( .A(n8481), .B(n8482), .Z(n8475) );
  XOR U9226 ( .A(n8483), .B(n8475), .Z(n8494) );
  XOR U9227 ( .A(sreg[1329]), .B(n8494), .Z(n8496) );
  NAND U9228 ( .A(n8476), .B(sreg[1328]), .Z(n8480) );
  NANDN U9229 ( .A(n8478), .B(n8477), .Z(n8479) );
  NAND U9230 ( .A(n8480), .B(n8479), .Z(n8495) );
  XNOR U9231 ( .A(n8496), .B(n8495), .Z(c[1329]) );
  AND U9232 ( .A(b[2]), .B(a[308]), .Z(n8509) );
  AND U9233 ( .A(a[309]), .B(b[1]), .Z(n8507) );
  AND U9234 ( .A(a[307]), .B(b[3]), .Z(n8506) );
  XOR U9235 ( .A(n8507), .B(n8506), .Z(n8508) );
  XOR U9236 ( .A(n8509), .B(n8508), .Z(n8512) );
  NAND U9237 ( .A(b[0]), .B(a[310]), .Z(n8513) );
  XOR U9238 ( .A(n8512), .B(n8513), .Z(n8515) );
  OR U9239 ( .A(n8485), .B(n8484), .Z(n8489) );
  NANDN U9240 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U9241 ( .A(n8489), .B(n8488), .Z(n8514) );
  XNOR U9242 ( .A(n8515), .B(n8514), .Z(n8500) );
  XNOR U9243 ( .A(n8500), .B(n8501), .Z(n8503) );
  XOR U9244 ( .A(n8502), .B(n8503), .Z(n8519) );
  NANDN U9245 ( .A(sreg[1329]), .B(n8494), .Z(n8498) );
  OR U9246 ( .A(n8496), .B(n8495), .Z(n8497) );
  AND U9247 ( .A(n8498), .B(n8497), .Z(n8518) );
  XNOR U9248 ( .A(sreg[1330]), .B(n8518), .Z(n8499) );
  XOR U9249 ( .A(n8519), .B(n8499), .Z(c[1330]) );
  NANDN U9250 ( .A(n8501), .B(n8500), .Z(n8505) );
  NAND U9251 ( .A(n8503), .B(n8502), .Z(n8504) );
  NAND U9252 ( .A(n8505), .B(n8504), .Z(n8536) );
  AND U9253 ( .A(b[2]), .B(a[309]), .Z(n8530) );
  AND U9254 ( .A(a[310]), .B(b[1]), .Z(n8528) );
  AND U9255 ( .A(a[308]), .B(b[3]), .Z(n8527) );
  XOR U9256 ( .A(n8528), .B(n8527), .Z(n8529) );
  XOR U9257 ( .A(n8530), .B(n8529), .Z(n8521) );
  NAND U9258 ( .A(b[0]), .B(a[311]), .Z(n8522) );
  XOR U9259 ( .A(n8521), .B(n8522), .Z(n8524) );
  OR U9260 ( .A(n8507), .B(n8506), .Z(n8511) );
  NANDN U9261 ( .A(n8509), .B(n8508), .Z(n8510) );
  NAND U9262 ( .A(n8511), .B(n8510), .Z(n8523) );
  XNOR U9263 ( .A(n8524), .B(n8523), .Z(n8533) );
  NANDN U9264 ( .A(n8513), .B(n8512), .Z(n8517) );
  OR U9265 ( .A(n8515), .B(n8514), .Z(n8516) );
  NAND U9266 ( .A(n8517), .B(n8516), .Z(n8534) );
  XNOR U9267 ( .A(n8533), .B(n8534), .Z(n8535) );
  XOR U9268 ( .A(n8536), .B(n8535), .Z(n8540) );
  XNOR U9269 ( .A(sreg[1331]), .B(n8539), .Z(n8520) );
  XOR U9270 ( .A(n8540), .B(n8520), .Z(c[1331]) );
  NANDN U9271 ( .A(n8522), .B(n8521), .Z(n8526) );
  OR U9272 ( .A(n8524), .B(n8523), .Z(n8525) );
  NAND U9273 ( .A(n8526), .B(n8525), .Z(n8542) );
  AND U9274 ( .A(b[2]), .B(a[310]), .Z(n8551) );
  AND U9275 ( .A(a[311]), .B(b[1]), .Z(n8549) );
  AND U9276 ( .A(a[309]), .B(b[3]), .Z(n8548) );
  XOR U9277 ( .A(n8549), .B(n8548), .Z(n8550) );
  XOR U9278 ( .A(n8551), .B(n8550), .Z(n8554) );
  NAND U9279 ( .A(b[0]), .B(a[312]), .Z(n8555) );
  XNOR U9280 ( .A(n8554), .B(n8555), .Z(n8556) );
  OR U9281 ( .A(n8528), .B(n8527), .Z(n8532) );
  NANDN U9282 ( .A(n8530), .B(n8529), .Z(n8531) );
  AND U9283 ( .A(n8532), .B(n8531), .Z(n8557) );
  XNOR U9284 ( .A(n8556), .B(n8557), .Z(n8543) );
  XNOR U9285 ( .A(n8542), .B(n8543), .Z(n8544) );
  NANDN U9286 ( .A(n8534), .B(n8533), .Z(n8538) );
  NAND U9287 ( .A(n8536), .B(n8535), .Z(n8537) );
  NAND U9288 ( .A(n8538), .B(n8537), .Z(n8545) );
  XNOR U9289 ( .A(n8544), .B(n8545), .Z(n8561) );
  XNOR U9290 ( .A(sreg[1332]), .B(n8560), .Z(n8541) );
  XOR U9291 ( .A(n8561), .B(n8541), .Z(c[1332]) );
  NANDN U9292 ( .A(n8543), .B(n8542), .Z(n8547) );
  NANDN U9293 ( .A(n8545), .B(n8544), .Z(n8546) );
  NAND U9294 ( .A(n8547), .B(n8546), .Z(n8566) );
  AND U9295 ( .A(b[2]), .B(a[311]), .Z(n8572) );
  AND U9296 ( .A(a[312]), .B(b[1]), .Z(n8570) );
  AND U9297 ( .A(a[310]), .B(b[3]), .Z(n8569) );
  XOR U9298 ( .A(n8570), .B(n8569), .Z(n8571) );
  XOR U9299 ( .A(n8572), .B(n8571), .Z(n8575) );
  NAND U9300 ( .A(b[0]), .B(a[313]), .Z(n8576) );
  XOR U9301 ( .A(n8575), .B(n8576), .Z(n8578) );
  OR U9302 ( .A(n8549), .B(n8548), .Z(n8553) );
  NANDN U9303 ( .A(n8551), .B(n8550), .Z(n8552) );
  NAND U9304 ( .A(n8553), .B(n8552), .Z(n8577) );
  XNOR U9305 ( .A(n8578), .B(n8577), .Z(n8563) );
  NANDN U9306 ( .A(n8555), .B(n8554), .Z(n8559) );
  NAND U9307 ( .A(n8557), .B(n8556), .Z(n8558) );
  NAND U9308 ( .A(n8559), .B(n8558), .Z(n8564) );
  XNOR U9309 ( .A(n8563), .B(n8564), .Z(n8565) );
  XOR U9310 ( .A(n8566), .B(n8565), .Z(n8582) );
  XNOR U9311 ( .A(sreg[1333]), .B(n8581), .Z(n8562) );
  XNOR U9312 ( .A(n8582), .B(n8562), .Z(c[1333]) );
  NANDN U9313 ( .A(n8564), .B(n8563), .Z(n8568) );
  NANDN U9314 ( .A(n8566), .B(n8565), .Z(n8567) );
  NAND U9315 ( .A(n8568), .B(n8567), .Z(n8587) );
  AND U9316 ( .A(b[2]), .B(a[312]), .Z(n8593) );
  AND U9317 ( .A(a[313]), .B(b[1]), .Z(n8591) );
  AND U9318 ( .A(a[311]), .B(b[3]), .Z(n8590) );
  XOR U9319 ( .A(n8591), .B(n8590), .Z(n8592) );
  XOR U9320 ( .A(n8593), .B(n8592), .Z(n8596) );
  NAND U9321 ( .A(b[0]), .B(a[314]), .Z(n8597) );
  XOR U9322 ( .A(n8596), .B(n8597), .Z(n8599) );
  OR U9323 ( .A(n8570), .B(n8569), .Z(n8574) );
  NANDN U9324 ( .A(n8572), .B(n8571), .Z(n8573) );
  NAND U9325 ( .A(n8574), .B(n8573), .Z(n8598) );
  XNOR U9326 ( .A(n8599), .B(n8598), .Z(n8584) );
  NANDN U9327 ( .A(n8576), .B(n8575), .Z(n8580) );
  OR U9328 ( .A(n8578), .B(n8577), .Z(n8579) );
  NAND U9329 ( .A(n8580), .B(n8579), .Z(n8585) );
  XNOR U9330 ( .A(n8584), .B(n8585), .Z(n8586) );
  XNOR U9331 ( .A(n8587), .B(n8586), .Z(n8603) );
  XOR U9332 ( .A(n8602), .B(sreg[1334]), .Z(n8583) );
  XOR U9333 ( .A(n8603), .B(n8583), .Z(c[1334]) );
  NANDN U9334 ( .A(n8585), .B(n8584), .Z(n8589) );
  NAND U9335 ( .A(n8587), .B(n8586), .Z(n8588) );
  NAND U9336 ( .A(n8589), .B(n8588), .Z(n8608) );
  AND U9337 ( .A(b[2]), .B(a[313]), .Z(n8614) );
  AND U9338 ( .A(a[314]), .B(b[1]), .Z(n8612) );
  AND U9339 ( .A(a[312]), .B(b[3]), .Z(n8611) );
  XOR U9340 ( .A(n8612), .B(n8611), .Z(n8613) );
  XOR U9341 ( .A(n8614), .B(n8613), .Z(n8617) );
  NAND U9342 ( .A(b[0]), .B(a[315]), .Z(n8618) );
  XOR U9343 ( .A(n8617), .B(n8618), .Z(n8620) );
  OR U9344 ( .A(n8591), .B(n8590), .Z(n8595) );
  NANDN U9345 ( .A(n8593), .B(n8592), .Z(n8594) );
  NAND U9346 ( .A(n8595), .B(n8594), .Z(n8619) );
  XNOR U9347 ( .A(n8620), .B(n8619), .Z(n8605) );
  NANDN U9348 ( .A(n8597), .B(n8596), .Z(n8601) );
  OR U9349 ( .A(n8599), .B(n8598), .Z(n8600) );
  NAND U9350 ( .A(n8601), .B(n8600), .Z(n8606) );
  XNOR U9351 ( .A(n8605), .B(n8606), .Z(n8607) );
  XNOR U9352 ( .A(n8608), .B(n8607), .Z(n8624) );
  XOR U9353 ( .A(n8623), .B(sreg[1335]), .Z(n8604) );
  XOR U9354 ( .A(n8624), .B(n8604), .Z(c[1335]) );
  NANDN U9355 ( .A(n8606), .B(n8605), .Z(n8610) );
  NAND U9356 ( .A(n8608), .B(n8607), .Z(n8609) );
  NAND U9357 ( .A(n8610), .B(n8609), .Z(n8629) );
  AND U9358 ( .A(b[2]), .B(a[314]), .Z(n8635) );
  AND U9359 ( .A(a[315]), .B(b[1]), .Z(n8633) );
  AND U9360 ( .A(a[313]), .B(b[3]), .Z(n8632) );
  XOR U9361 ( .A(n8633), .B(n8632), .Z(n8634) );
  XOR U9362 ( .A(n8635), .B(n8634), .Z(n8638) );
  NAND U9363 ( .A(b[0]), .B(a[316]), .Z(n8639) );
  XOR U9364 ( .A(n8638), .B(n8639), .Z(n8641) );
  OR U9365 ( .A(n8612), .B(n8611), .Z(n8616) );
  NANDN U9366 ( .A(n8614), .B(n8613), .Z(n8615) );
  NAND U9367 ( .A(n8616), .B(n8615), .Z(n8640) );
  XNOR U9368 ( .A(n8641), .B(n8640), .Z(n8626) );
  NANDN U9369 ( .A(n8618), .B(n8617), .Z(n8622) );
  OR U9370 ( .A(n8620), .B(n8619), .Z(n8621) );
  NAND U9371 ( .A(n8622), .B(n8621), .Z(n8627) );
  XNOR U9372 ( .A(n8626), .B(n8627), .Z(n8628) );
  XOR U9373 ( .A(n8629), .B(n8628), .Z(n8645) );
  XOR U9374 ( .A(sreg[1336]), .B(n8644), .Z(n8625) );
  XOR U9375 ( .A(n8645), .B(n8625), .Z(c[1336]) );
  NANDN U9376 ( .A(n8627), .B(n8626), .Z(n8631) );
  NAND U9377 ( .A(n8629), .B(n8628), .Z(n8630) );
  NAND U9378 ( .A(n8631), .B(n8630), .Z(n8652) );
  AND U9379 ( .A(b[2]), .B(a[315]), .Z(n8658) );
  AND U9380 ( .A(a[316]), .B(b[1]), .Z(n8656) );
  AND U9381 ( .A(a[314]), .B(b[3]), .Z(n8655) );
  XOR U9382 ( .A(n8656), .B(n8655), .Z(n8657) );
  XOR U9383 ( .A(n8658), .B(n8657), .Z(n8661) );
  NAND U9384 ( .A(b[0]), .B(a[317]), .Z(n8662) );
  XOR U9385 ( .A(n8661), .B(n8662), .Z(n8664) );
  OR U9386 ( .A(n8633), .B(n8632), .Z(n8637) );
  NANDN U9387 ( .A(n8635), .B(n8634), .Z(n8636) );
  NAND U9388 ( .A(n8637), .B(n8636), .Z(n8663) );
  XNOR U9389 ( .A(n8664), .B(n8663), .Z(n8649) );
  NANDN U9390 ( .A(n8639), .B(n8638), .Z(n8643) );
  OR U9391 ( .A(n8641), .B(n8640), .Z(n8642) );
  NAND U9392 ( .A(n8643), .B(n8642), .Z(n8650) );
  XNOR U9393 ( .A(n8649), .B(n8650), .Z(n8651) );
  XNOR U9394 ( .A(n8652), .B(n8651), .Z(n8648) );
  XOR U9395 ( .A(n8647), .B(sreg[1337]), .Z(n8646) );
  XOR U9396 ( .A(n8648), .B(n8646), .Z(c[1337]) );
  NANDN U9397 ( .A(n8650), .B(n8649), .Z(n8654) );
  NAND U9398 ( .A(n8652), .B(n8651), .Z(n8653) );
  NAND U9399 ( .A(n8654), .B(n8653), .Z(n8670) );
  AND U9400 ( .A(b[2]), .B(a[316]), .Z(n8676) );
  AND U9401 ( .A(a[317]), .B(b[1]), .Z(n8674) );
  AND U9402 ( .A(a[315]), .B(b[3]), .Z(n8673) );
  XOR U9403 ( .A(n8674), .B(n8673), .Z(n8675) );
  XOR U9404 ( .A(n8676), .B(n8675), .Z(n8679) );
  NAND U9405 ( .A(b[0]), .B(a[318]), .Z(n8680) );
  XOR U9406 ( .A(n8679), .B(n8680), .Z(n8682) );
  OR U9407 ( .A(n8656), .B(n8655), .Z(n8660) );
  NANDN U9408 ( .A(n8658), .B(n8657), .Z(n8659) );
  NAND U9409 ( .A(n8660), .B(n8659), .Z(n8681) );
  XNOR U9410 ( .A(n8682), .B(n8681), .Z(n8667) );
  NANDN U9411 ( .A(n8662), .B(n8661), .Z(n8666) );
  OR U9412 ( .A(n8664), .B(n8663), .Z(n8665) );
  NAND U9413 ( .A(n8666), .B(n8665), .Z(n8668) );
  XNOR U9414 ( .A(n8667), .B(n8668), .Z(n8669) );
  XNOR U9415 ( .A(n8670), .B(n8669), .Z(n8685) );
  XNOR U9416 ( .A(n8685), .B(sreg[1338]), .Z(n8687) );
  XNOR U9417 ( .A(n8686), .B(n8687), .Z(c[1338]) );
  NANDN U9418 ( .A(n8668), .B(n8667), .Z(n8672) );
  NAND U9419 ( .A(n8670), .B(n8669), .Z(n8671) );
  NAND U9420 ( .A(n8672), .B(n8671), .Z(n8693) );
  AND U9421 ( .A(b[2]), .B(a[317]), .Z(n8699) );
  AND U9422 ( .A(a[318]), .B(b[1]), .Z(n8697) );
  AND U9423 ( .A(a[316]), .B(b[3]), .Z(n8696) );
  XOR U9424 ( .A(n8697), .B(n8696), .Z(n8698) );
  XOR U9425 ( .A(n8699), .B(n8698), .Z(n8702) );
  NAND U9426 ( .A(b[0]), .B(a[319]), .Z(n8703) );
  XOR U9427 ( .A(n8702), .B(n8703), .Z(n8705) );
  OR U9428 ( .A(n8674), .B(n8673), .Z(n8678) );
  NANDN U9429 ( .A(n8676), .B(n8675), .Z(n8677) );
  NAND U9430 ( .A(n8678), .B(n8677), .Z(n8704) );
  XNOR U9431 ( .A(n8705), .B(n8704), .Z(n8690) );
  NANDN U9432 ( .A(n8680), .B(n8679), .Z(n8684) );
  OR U9433 ( .A(n8682), .B(n8681), .Z(n8683) );
  NAND U9434 ( .A(n8684), .B(n8683), .Z(n8691) );
  XNOR U9435 ( .A(n8690), .B(n8691), .Z(n8692) );
  XNOR U9436 ( .A(n8693), .B(n8692), .Z(n8708) );
  XOR U9437 ( .A(sreg[1339]), .B(n8708), .Z(n8709) );
  NAND U9438 ( .A(n8685), .B(sreg[1338]), .Z(n8689) );
  NANDN U9439 ( .A(n8687), .B(n8686), .Z(n8688) );
  NAND U9440 ( .A(n8689), .B(n8688), .Z(n8710) );
  XOR U9441 ( .A(n8709), .B(n8710), .Z(c[1339]) );
  NANDN U9442 ( .A(n8691), .B(n8690), .Z(n8695) );
  NAND U9443 ( .A(n8693), .B(n8692), .Z(n8694) );
  NAND U9444 ( .A(n8695), .B(n8694), .Z(n8719) );
  AND U9445 ( .A(b[2]), .B(a[318]), .Z(n8725) );
  AND U9446 ( .A(a[319]), .B(b[1]), .Z(n8723) );
  AND U9447 ( .A(a[317]), .B(b[3]), .Z(n8722) );
  XOR U9448 ( .A(n8723), .B(n8722), .Z(n8724) );
  XOR U9449 ( .A(n8725), .B(n8724), .Z(n8728) );
  NAND U9450 ( .A(b[0]), .B(a[320]), .Z(n8729) );
  XOR U9451 ( .A(n8728), .B(n8729), .Z(n8731) );
  OR U9452 ( .A(n8697), .B(n8696), .Z(n8701) );
  NANDN U9453 ( .A(n8699), .B(n8698), .Z(n8700) );
  NAND U9454 ( .A(n8701), .B(n8700), .Z(n8730) );
  XNOR U9455 ( .A(n8731), .B(n8730), .Z(n8716) );
  NANDN U9456 ( .A(n8703), .B(n8702), .Z(n8707) );
  OR U9457 ( .A(n8705), .B(n8704), .Z(n8706) );
  NAND U9458 ( .A(n8707), .B(n8706), .Z(n8717) );
  XNOR U9459 ( .A(n8716), .B(n8717), .Z(n8718) );
  XOR U9460 ( .A(n8719), .B(n8718), .Z(n8715) );
  OR U9461 ( .A(n8708), .B(sreg[1339]), .Z(n8712) );
  NANDN U9462 ( .A(n8710), .B(n8709), .Z(n8711) );
  AND U9463 ( .A(n8712), .B(n8711), .Z(n8714) );
  XNOR U9464 ( .A(sreg[1340]), .B(n8714), .Z(n8713) );
  XOR U9465 ( .A(n8715), .B(n8713), .Z(c[1340]) );
  NANDN U9466 ( .A(n8717), .B(n8716), .Z(n8721) );
  NAND U9467 ( .A(n8719), .B(n8718), .Z(n8720) );
  NAND U9468 ( .A(n8721), .B(n8720), .Z(n8737) );
  AND U9469 ( .A(b[2]), .B(a[319]), .Z(n8743) );
  AND U9470 ( .A(a[320]), .B(b[1]), .Z(n8741) );
  AND U9471 ( .A(a[318]), .B(b[3]), .Z(n8740) );
  XOR U9472 ( .A(n8741), .B(n8740), .Z(n8742) );
  XOR U9473 ( .A(n8743), .B(n8742), .Z(n8746) );
  NAND U9474 ( .A(b[0]), .B(a[321]), .Z(n8747) );
  XOR U9475 ( .A(n8746), .B(n8747), .Z(n8749) );
  OR U9476 ( .A(n8723), .B(n8722), .Z(n8727) );
  NANDN U9477 ( .A(n8725), .B(n8724), .Z(n8726) );
  NAND U9478 ( .A(n8727), .B(n8726), .Z(n8748) );
  XNOR U9479 ( .A(n8749), .B(n8748), .Z(n8734) );
  NANDN U9480 ( .A(n8729), .B(n8728), .Z(n8733) );
  OR U9481 ( .A(n8731), .B(n8730), .Z(n8732) );
  NAND U9482 ( .A(n8733), .B(n8732), .Z(n8735) );
  XNOR U9483 ( .A(n8734), .B(n8735), .Z(n8736) );
  XNOR U9484 ( .A(n8737), .B(n8736), .Z(n8752) );
  XNOR U9485 ( .A(n8752), .B(sreg[1341]), .Z(n8753) );
  XOR U9486 ( .A(n8754), .B(n8753), .Z(c[1341]) );
  NANDN U9487 ( .A(n8735), .B(n8734), .Z(n8739) );
  NAND U9488 ( .A(n8737), .B(n8736), .Z(n8738) );
  NAND U9489 ( .A(n8739), .B(n8738), .Z(n8763) );
  AND U9490 ( .A(b[2]), .B(a[320]), .Z(n8769) );
  AND U9491 ( .A(a[321]), .B(b[1]), .Z(n8767) );
  AND U9492 ( .A(a[319]), .B(b[3]), .Z(n8766) );
  XOR U9493 ( .A(n8767), .B(n8766), .Z(n8768) );
  XOR U9494 ( .A(n8769), .B(n8768), .Z(n8772) );
  NAND U9495 ( .A(b[0]), .B(a[322]), .Z(n8773) );
  XOR U9496 ( .A(n8772), .B(n8773), .Z(n8775) );
  OR U9497 ( .A(n8741), .B(n8740), .Z(n8745) );
  NANDN U9498 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U9499 ( .A(n8745), .B(n8744), .Z(n8774) );
  XNOR U9500 ( .A(n8775), .B(n8774), .Z(n8760) );
  NANDN U9501 ( .A(n8747), .B(n8746), .Z(n8751) );
  OR U9502 ( .A(n8749), .B(n8748), .Z(n8750) );
  NAND U9503 ( .A(n8751), .B(n8750), .Z(n8761) );
  XNOR U9504 ( .A(n8760), .B(n8761), .Z(n8762) );
  XOR U9505 ( .A(n8763), .B(n8762), .Z(n8759) );
  NAND U9506 ( .A(n8752), .B(sreg[1341]), .Z(n8756) );
  OR U9507 ( .A(n8754), .B(n8753), .Z(n8755) );
  NAND U9508 ( .A(n8756), .B(n8755), .Z(n8758) );
  XNOR U9509 ( .A(sreg[1342]), .B(n8758), .Z(n8757) );
  XOR U9510 ( .A(n8759), .B(n8757), .Z(c[1342]) );
  NANDN U9511 ( .A(n8761), .B(n8760), .Z(n8765) );
  NAND U9512 ( .A(n8763), .B(n8762), .Z(n8764) );
  NAND U9513 ( .A(n8765), .B(n8764), .Z(n8781) );
  AND U9514 ( .A(b[2]), .B(a[321]), .Z(n8787) );
  AND U9515 ( .A(a[322]), .B(b[1]), .Z(n8785) );
  AND U9516 ( .A(a[320]), .B(b[3]), .Z(n8784) );
  XOR U9517 ( .A(n8785), .B(n8784), .Z(n8786) );
  XOR U9518 ( .A(n8787), .B(n8786), .Z(n8790) );
  NAND U9519 ( .A(b[0]), .B(a[323]), .Z(n8791) );
  XOR U9520 ( .A(n8790), .B(n8791), .Z(n8793) );
  OR U9521 ( .A(n8767), .B(n8766), .Z(n8771) );
  NANDN U9522 ( .A(n8769), .B(n8768), .Z(n8770) );
  NAND U9523 ( .A(n8771), .B(n8770), .Z(n8792) );
  XNOR U9524 ( .A(n8793), .B(n8792), .Z(n8778) );
  NANDN U9525 ( .A(n8773), .B(n8772), .Z(n8777) );
  OR U9526 ( .A(n8775), .B(n8774), .Z(n8776) );
  NAND U9527 ( .A(n8777), .B(n8776), .Z(n8779) );
  XNOR U9528 ( .A(n8778), .B(n8779), .Z(n8780) );
  XNOR U9529 ( .A(n8781), .B(n8780), .Z(n8796) );
  XNOR U9530 ( .A(n8796), .B(sreg[1343]), .Z(n8797) );
  XOR U9531 ( .A(n8798), .B(n8797), .Z(c[1343]) );
  NANDN U9532 ( .A(n8779), .B(n8778), .Z(n8783) );
  NAND U9533 ( .A(n8781), .B(n8780), .Z(n8782) );
  NAND U9534 ( .A(n8783), .B(n8782), .Z(n8809) );
  AND U9535 ( .A(b[2]), .B(a[322]), .Z(n8821) );
  AND U9536 ( .A(a[323]), .B(b[1]), .Z(n8819) );
  AND U9537 ( .A(a[321]), .B(b[3]), .Z(n8818) );
  XOR U9538 ( .A(n8819), .B(n8818), .Z(n8820) );
  XOR U9539 ( .A(n8821), .B(n8820), .Z(n8812) );
  NAND U9540 ( .A(b[0]), .B(a[324]), .Z(n8813) );
  XOR U9541 ( .A(n8812), .B(n8813), .Z(n8815) );
  OR U9542 ( .A(n8785), .B(n8784), .Z(n8789) );
  NANDN U9543 ( .A(n8787), .B(n8786), .Z(n8788) );
  NAND U9544 ( .A(n8789), .B(n8788), .Z(n8814) );
  XNOR U9545 ( .A(n8815), .B(n8814), .Z(n8806) );
  NANDN U9546 ( .A(n8791), .B(n8790), .Z(n8795) );
  OR U9547 ( .A(n8793), .B(n8792), .Z(n8794) );
  NAND U9548 ( .A(n8795), .B(n8794), .Z(n8807) );
  XNOR U9549 ( .A(n8806), .B(n8807), .Z(n8808) );
  XNOR U9550 ( .A(n8809), .B(n8808), .Z(n8801) );
  XNOR U9551 ( .A(n8801), .B(sreg[1344]), .Z(n8803) );
  NAND U9552 ( .A(n8796), .B(sreg[1343]), .Z(n8800) );
  OR U9553 ( .A(n8798), .B(n8797), .Z(n8799) );
  AND U9554 ( .A(n8800), .B(n8799), .Z(n8802) );
  XOR U9555 ( .A(n8803), .B(n8802), .Z(c[1344]) );
  NAND U9556 ( .A(n8801), .B(sreg[1344]), .Z(n8805) );
  OR U9557 ( .A(n8803), .B(n8802), .Z(n8804) );
  NAND U9558 ( .A(n8805), .B(n8804), .Z(n8843) );
  NANDN U9559 ( .A(n8807), .B(n8806), .Z(n8811) );
  NAND U9560 ( .A(n8809), .B(n8808), .Z(n8810) );
  NAND U9561 ( .A(n8811), .B(n8810), .Z(n8840) );
  NANDN U9562 ( .A(n8813), .B(n8812), .Z(n8817) );
  OR U9563 ( .A(n8815), .B(n8814), .Z(n8816) );
  NAND U9564 ( .A(n8817), .B(n8816), .Z(n8837) );
  AND U9565 ( .A(b[2]), .B(a[323]), .Z(n8828) );
  AND U9566 ( .A(a[324]), .B(b[1]), .Z(n8826) );
  AND U9567 ( .A(a[322]), .B(b[3]), .Z(n8825) );
  XOR U9568 ( .A(n8826), .B(n8825), .Z(n8827) );
  XOR U9569 ( .A(n8828), .B(n8827), .Z(n8831) );
  NAND U9570 ( .A(b[0]), .B(a[325]), .Z(n8832) );
  XNOR U9571 ( .A(n8831), .B(n8832), .Z(n8833) );
  OR U9572 ( .A(n8819), .B(n8818), .Z(n8823) );
  NANDN U9573 ( .A(n8821), .B(n8820), .Z(n8822) );
  AND U9574 ( .A(n8823), .B(n8822), .Z(n8834) );
  XNOR U9575 ( .A(n8833), .B(n8834), .Z(n8838) );
  XNOR U9576 ( .A(n8837), .B(n8838), .Z(n8839) );
  XNOR U9577 ( .A(n8840), .B(n8839), .Z(n8844) );
  XNOR U9578 ( .A(sreg[1345]), .B(n8844), .Z(n8824) );
  XNOR U9579 ( .A(n8843), .B(n8824), .Z(c[1345]) );
  AND U9580 ( .A(b[2]), .B(a[324]), .Z(n8857) );
  AND U9581 ( .A(a[325]), .B(b[1]), .Z(n8855) );
  AND U9582 ( .A(a[323]), .B(b[3]), .Z(n8854) );
  XOR U9583 ( .A(n8855), .B(n8854), .Z(n8856) );
  XOR U9584 ( .A(n8857), .B(n8856), .Z(n8860) );
  NAND U9585 ( .A(b[0]), .B(a[326]), .Z(n8861) );
  XOR U9586 ( .A(n8860), .B(n8861), .Z(n8863) );
  OR U9587 ( .A(n8826), .B(n8825), .Z(n8830) );
  NANDN U9588 ( .A(n8828), .B(n8827), .Z(n8829) );
  NAND U9589 ( .A(n8830), .B(n8829), .Z(n8862) );
  XNOR U9590 ( .A(n8863), .B(n8862), .Z(n8848) );
  NANDN U9591 ( .A(n8832), .B(n8831), .Z(n8836) );
  NAND U9592 ( .A(n8834), .B(n8833), .Z(n8835) );
  NAND U9593 ( .A(n8836), .B(n8835), .Z(n8849) );
  XNOR U9594 ( .A(n8848), .B(n8849), .Z(n8850) );
  NANDN U9595 ( .A(n8838), .B(n8837), .Z(n8842) );
  NANDN U9596 ( .A(n8840), .B(n8839), .Z(n8841) );
  AND U9597 ( .A(n8842), .B(n8841), .Z(n8851) );
  XNOR U9598 ( .A(n8850), .B(n8851), .Z(n8847) );
  XNOR U9599 ( .A(sreg[1346]), .B(n8846), .Z(n8845) );
  XOR U9600 ( .A(n8847), .B(n8845), .Z(c[1346]) );
  NANDN U9601 ( .A(n8849), .B(n8848), .Z(n8853) );
  NAND U9602 ( .A(n8851), .B(n8850), .Z(n8852) );
  NAND U9603 ( .A(n8853), .B(n8852), .Z(n8881) );
  AND U9604 ( .A(b[2]), .B(a[325]), .Z(n8875) );
  AND U9605 ( .A(a[326]), .B(b[1]), .Z(n8873) );
  AND U9606 ( .A(a[324]), .B(b[3]), .Z(n8872) );
  XOR U9607 ( .A(n8873), .B(n8872), .Z(n8874) );
  XOR U9608 ( .A(n8875), .B(n8874), .Z(n8866) );
  NAND U9609 ( .A(b[0]), .B(a[327]), .Z(n8867) );
  XOR U9610 ( .A(n8866), .B(n8867), .Z(n8869) );
  OR U9611 ( .A(n8855), .B(n8854), .Z(n8859) );
  NANDN U9612 ( .A(n8857), .B(n8856), .Z(n8858) );
  NAND U9613 ( .A(n8859), .B(n8858), .Z(n8868) );
  XNOR U9614 ( .A(n8869), .B(n8868), .Z(n8878) );
  NANDN U9615 ( .A(n8861), .B(n8860), .Z(n8865) );
  OR U9616 ( .A(n8863), .B(n8862), .Z(n8864) );
  NAND U9617 ( .A(n8865), .B(n8864), .Z(n8879) );
  XNOR U9618 ( .A(n8878), .B(n8879), .Z(n8880) );
  XNOR U9619 ( .A(n8881), .B(n8880), .Z(n8884) );
  XNOR U9620 ( .A(n8884), .B(sreg[1347]), .Z(n8885) );
  XOR U9621 ( .A(n8886), .B(n8885), .Z(c[1347]) );
  NANDN U9622 ( .A(n8867), .B(n8866), .Z(n8871) );
  OR U9623 ( .A(n8869), .B(n8868), .Z(n8870) );
  NAND U9624 ( .A(n8871), .B(n8870), .Z(n8892) );
  AND U9625 ( .A(b[2]), .B(a[326]), .Z(n8907) );
  AND U9626 ( .A(a[327]), .B(b[1]), .Z(n8905) );
  AND U9627 ( .A(a[325]), .B(b[3]), .Z(n8904) );
  XOR U9628 ( .A(n8905), .B(n8904), .Z(n8906) );
  XOR U9629 ( .A(n8907), .B(n8906), .Z(n8898) );
  NAND U9630 ( .A(b[0]), .B(a[328]), .Z(n8899) );
  XNOR U9631 ( .A(n8898), .B(n8899), .Z(n8900) );
  OR U9632 ( .A(n8873), .B(n8872), .Z(n8877) );
  NANDN U9633 ( .A(n8875), .B(n8874), .Z(n8876) );
  AND U9634 ( .A(n8877), .B(n8876), .Z(n8901) );
  XNOR U9635 ( .A(n8900), .B(n8901), .Z(n8893) );
  XNOR U9636 ( .A(n8892), .B(n8893), .Z(n8894) );
  NANDN U9637 ( .A(n8879), .B(n8878), .Z(n8883) );
  NAND U9638 ( .A(n8881), .B(n8880), .Z(n8882) );
  NAND U9639 ( .A(n8883), .B(n8882), .Z(n8895) );
  XOR U9640 ( .A(n8894), .B(n8895), .Z(n8891) );
  NAND U9641 ( .A(n8884), .B(sreg[1347]), .Z(n8888) );
  OR U9642 ( .A(n8886), .B(n8885), .Z(n8887) );
  AND U9643 ( .A(n8888), .B(n8887), .Z(n8890) );
  XNOR U9644 ( .A(n8890), .B(sreg[1348]), .Z(n8889) );
  XNOR U9645 ( .A(n8891), .B(n8889), .Z(c[1348]) );
  NANDN U9646 ( .A(n8893), .B(n8892), .Z(n8897) );
  NANDN U9647 ( .A(n8895), .B(n8894), .Z(n8896) );
  NAND U9648 ( .A(n8897), .B(n8896), .Z(n8913) );
  NANDN U9649 ( .A(n8899), .B(n8898), .Z(n8903) );
  NAND U9650 ( .A(n8901), .B(n8900), .Z(n8902) );
  NAND U9651 ( .A(n8903), .B(n8902), .Z(n8910) );
  AND U9652 ( .A(b[2]), .B(a[327]), .Z(n8919) );
  AND U9653 ( .A(a[328]), .B(b[1]), .Z(n8917) );
  AND U9654 ( .A(a[326]), .B(b[3]), .Z(n8916) );
  XOR U9655 ( .A(n8917), .B(n8916), .Z(n8918) );
  XOR U9656 ( .A(n8919), .B(n8918), .Z(n8922) );
  NAND U9657 ( .A(b[0]), .B(a[329]), .Z(n8923) );
  XNOR U9658 ( .A(n8922), .B(n8923), .Z(n8924) );
  OR U9659 ( .A(n8905), .B(n8904), .Z(n8909) );
  NANDN U9660 ( .A(n8907), .B(n8906), .Z(n8908) );
  AND U9661 ( .A(n8909), .B(n8908), .Z(n8925) );
  XNOR U9662 ( .A(n8924), .B(n8925), .Z(n8911) );
  XNOR U9663 ( .A(n8910), .B(n8911), .Z(n8912) );
  XOR U9664 ( .A(n8913), .B(n8912), .Z(n8928) );
  XNOR U9665 ( .A(sreg[1349]), .B(n8928), .Z(n8930) );
  XNOR U9666 ( .A(n8929), .B(n8930), .Z(c[1349]) );
  NANDN U9667 ( .A(n8911), .B(n8910), .Z(n8915) );
  NAND U9668 ( .A(n8913), .B(n8912), .Z(n8914) );
  NAND U9669 ( .A(n8915), .B(n8914), .Z(n8936) );
  AND U9670 ( .A(b[2]), .B(a[328]), .Z(n8942) );
  AND U9671 ( .A(a[329]), .B(b[1]), .Z(n8940) );
  AND U9672 ( .A(a[327]), .B(b[3]), .Z(n8939) );
  XOR U9673 ( .A(n8940), .B(n8939), .Z(n8941) );
  XOR U9674 ( .A(n8942), .B(n8941), .Z(n8945) );
  NAND U9675 ( .A(b[0]), .B(a[330]), .Z(n8946) );
  XOR U9676 ( .A(n8945), .B(n8946), .Z(n8948) );
  OR U9677 ( .A(n8917), .B(n8916), .Z(n8921) );
  NANDN U9678 ( .A(n8919), .B(n8918), .Z(n8920) );
  NAND U9679 ( .A(n8921), .B(n8920), .Z(n8947) );
  XNOR U9680 ( .A(n8948), .B(n8947), .Z(n8933) );
  NANDN U9681 ( .A(n8923), .B(n8922), .Z(n8927) );
  NAND U9682 ( .A(n8925), .B(n8924), .Z(n8926) );
  NAND U9683 ( .A(n8927), .B(n8926), .Z(n8934) );
  XNOR U9684 ( .A(n8933), .B(n8934), .Z(n8935) );
  XOR U9685 ( .A(n8936), .B(n8935), .Z(n8951) );
  XNOR U9686 ( .A(n8951), .B(sreg[1350]), .Z(n8953) );
  NAND U9687 ( .A(sreg[1349]), .B(n8928), .Z(n8932) );
  NANDN U9688 ( .A(n8930), .B(n8929), .Z(n8931) );
  AND U9689 ( .A(n8932), .B(n8931), .Z(n8952) );
  XOR U9690 ( .A(n8953), .B(n8952), .Z(c[1350]) );
  NANDN U9691 ( .A(n8934), .B(n8933), .Z(n8938) );
  NANDN U9692 ( .A(n8936), .B(n8935), .Z(n8937) );
  NAND U9693 ( .A(n8938), .B(n8937), .Z(n8971) );
  AND U9694 ( .A(b[2]), .B(a[329]), .Z(n8965) );
  AND U9695 ( .A(a[330]), .B(b[1]), .Z(n8963) );
  AND U9696 ( .A(a[328]), .B(b[3]), .Z(n8962) );
  XOR U9697 ( .A(n8963), .B(n8962), .Z(n8964) );
  XOR U9698 ( .A(n8965), .B(n8964), .Z(n8956) );
  NAND U9699 ( .A(b[0]), .B(a[331]), .Z(n8957) );
  XOR U9700 ( .A(n8956), .B(n8957), .Z(n8959) );
  OR U9701 ( .A(n8940), .B(n8939), .Z(n8944) );
  NANDN U9702 ( .A(n8942), .B(n8941), .Z(n8943) );
  NAND U9703 ( .A(n8944), .B(n8943), .Z(n8958) );
  XNOR U9704 ( .A(n8959), .B(n8958), .Z(n8968) );
  NANDN U9705 ( .A(n8946), .B(n8945), .Z(n8950) );
  OR U9706 ( .A(n8948), .B(n8947), .Z(n8949) );
  NAND U9707 ( .A(n8950), .B(n8949), .Z(n8969) );
  XNOR U9708 ( .A(n8968), .B(n8969), .Z(n8970) );
  XNOR U9709 ( .A(n8971), .B(n8970), .Z(n8974) );
  XNOR U9710 ( .A(n8974), .B(sreg[1351]), .Z(n8976) );
  NAND U9711 ( .A(n8951), .B(sreg[1350]), .Z(n8955) );
  OR U9712 ( .A(n8953), .B(n8952), .Z(n8954) );
  AND U9713 ( .A(n8955), .B(n8954), .Z(n8975) );
  XOR U9714 ( .A(n8976), .B(n8975), .Z(c[1351]) );
  NANDN U9715 ( .A(n8957), .B(n8956), .Z(n8961) );
  OR U9716 ( .A(n8959), .B(n8958), .Z(n8960) );
  NAND U9717 ( .A(n8961), .B(n8960), .Z(n8979) );
  AND U9718 ( .A(b[2]), .B(a[330]), .Z(n8988) );
  AND U9719 ( .A(a[331]), .B(b[1]), .Z(n8986) );
  AND U9720 ( .A(a[329]), .B(b[3]), .Z(n8985) );
  XOR U9721 ( .A(n8986), .B(n8985), .Z(n8987) );
  XOR U9722 ( .A(n8988), .B(n8987), .Z(n8991) );
  NAND U9723 ( .A(b[0]), .B(a[332]), .Z(n8992) );
  XNOR U9724 ( .A(n8991), .B(n8992), .Z(n8993) );
  OR U9725 ( .A(n8963), .B(n8962), .Z(n8967) );
  NANDN U9726 ( .A(n8965), .B(n8964), .Z(n8966) );
  AND U9727 ( .A(n8967), .B(n8966), .Z(n8994) );
  XNOR U9728 ( .A(n8993), .B(n8994), .Z(n8980) );
  XNOR U9729 ( .A(n8979), .B(n8980), .Z(n8981) );
  NANDN U9730 ( .A(n8969), .B(n8968), .Z(n8973) );
  NAND U9731 ( .A(n8971), .B(n8970), .Z(n8972) );
  AND U9732 ( .A(n8973), .B(n8972), .Z(n8982) );
  XOR U9733 ( .A(n8981), .B(n8982), .Z(n8997) );
  XNOR U9734 ( .A(sreg[1352]), .B(n8997), .Z(n8999) );
  NAND U9735 ( .A(n8974), .B(sreg[1351]), .Z(n8978) );
  OR U9736 ( .A(n8976), .B(n8975), .Z(n8977) );
  AND U9737 ( .A(n8978), .B(n8977), .Z(n8998) );
  XOR U9738 ( .A(n8999), .B(n8998), .Z(c[1352]) );
  NANDN U9739 ( .A(n8980), .B(n8979), .Z(n8984) );
  NAND U9740 ( .A(n8982), .B(n8981), .Z(n8983) );
  NAND U9741 ( .A(n8984), .B(n8983), .Z(n9010) );
  AND U9742 ( .A(b[2]), .B(a[331]), .Z(n9016) );
  AND U9743 ( .A(a[332]), .B(b[1]), .Z(n9014) );
  AND U9744 ( .A(a[330]), .B(b[3]), .Z(n9013) );
  XOR U9745 ( .A(n9014), .B(n9013), .Z(n9015) );
  XOR U9746 ( .A(n9016), .B(n9015), .Z(n9019) );
  NAND U9747 ( .A(b[0]), .B(a[333]), .Z(n9020) );
  XOR U9748 ( .A(n9019), .B(n9020), .Z(n9022) );
  OR U9749 ( .A(n8986), .B(n8985), .Z(n8990) );
  NANDN U9750 ( .A(n8988), .B(n8987), .Z(n8989) );
  NAND U9751 ( .A(n8990), .B(n8989), .Z(n9021) );
  XNOR U9752 ( .A(n9022), .B(n9021), .Z(n9007) );
  NANDN U9753 ( .A(n8992), .B(n8991), .Z(n8996) );
  NAND U9754 ( .A(n8994), .B(n8993), .Z(n8995) );
  NAND U9755 ( .A(n8996), .B(n8995), .Z(n9008) );
  XNOR U9756 ( .A(n9007), .B(n9008), .Z(n9009) );
  XOR U9757 ( .A(n9010), .B(n9009), .Z(n9002) );
  XNOR U9758 ( .A(n9002), .B(sreg[1353]), .Z(n9004) );
  NAND U9759 ( .A(sreg[1352]), .B(n8997), .Z(n9001) );
  OR U9760 ( .A(n8999), .B(n8998), .Z(n9000) );
  AND U9761 ( .A(n9001), .B(n9000), .Z(n9003) );
  XOR U9762 ( .A(n9004), .B(n9003), .Z(c[1353]) );
  NAND U9763 ( .A(n9002), .B(sreg[1353]), .Z(n9006) );
  OR U9764 ( .A(n9004), .B(n9003), .Z(n9005) );
  AND U9765 ( .A(n9006), .B(n9005), .Z(n9045) );
  NANDN U9766 ( .A(n9008), .B(n9007), .Z(n9012) );
  NANDN U9767 ( .A(n9010), .B(n9009), .Z(n9011) );
  NAND U9768 ( .A(n9012), .B(n9011), .Z(n9029) );
  AND U9769 ( .A(b[2]), .B(a[332]), .Z(n9035) );
  AND U9770 ( .A(a[333]), .B(b[1]), .Z(n9033) );
  AND U9771 ( .A(a[331]), .B(b[3]), .Z(n9032) );
  XOR U9772 ( .A(n9033), .B(n9032), .Z(n9034) );
  XOR U9773 ( .A(n9035), .B(n9034), .Z(n9038) );
  NAND U9774 ( .A(b[0]), .B(a[334]), .Z(n9039) );
  XOR U9775 ( .A(n9038), .B(n9039), .Z(n9041) );
  OR U9776 ( .A(n9014), .B(n9013), .Z(n9018) );
  NANDN U9777 ( .A(n9016), .B(n9015), .Z(n9017) );
  NAND U9778 ( .A(n9018), .B(n9017), .Z(n9040) );
  XNOR U9779 ( .A(n9041), .B(n9040), .Z(n9026) );
  NANDN U9780 ( .A(n9020), .B(n9019), .Z(n9024) );
  OR U9781 ( .A(n9022), .B(n9021), .Z(n9023) );
  NAND U9782 ( .A(n9024), .B(n9023), .Z(n9027) );
  XNOR U9783 ( .A(n9026), .B(n9027), .Z(n9028) );
  XNOR U9784 ( .A(n9029), .B(n9028), .Z(n9044) );
  XNOR U9785 ( .A(sreg[1354]), .B(n9044), .Z(n9025) );
  XOR U9786 ( .A(n9045), .B(n9025), .Z(c[1354]) );
  NANDN U9787 ( .A(n9027), .B(n9026), .Z(n9031) );
  NAND U9788 ( .A(n9029), .B(n9028), .Z(n9030) );
  NAND U9789 ( .A(n9031), .B(n9030), .Z(n9052) );
  AND U9790 ( .A(b[2]), .B(a[333]), .Z(n9058) );
  AND U9791 ( .A(a[334]), .B(b[1]), .Z(n9056) );
  AND U9792 ( .A(a[332]), .B(b[3]), .Z(n9055) );
  XOR U9793 ( .A(n9056), .B(n9055), .Z(n9057) );
  XOR U9794 ( .A(n9058), .B(n9057), .Z(n9061) );
  NAND U9795 ( .A(b[0]), .B(a[335]), .Z(n9062) );
  XOR U9796 ( .A(n9061), .B(n9062), .Z(n9064) );
  OR U9797 ( .A(n9033), .B(n9032), .Z(n9037) );
  NANDN U9798 ( .A(n9035), .B(n9034), .Z(n9036) );
  NAND U9799 ( .A(n9037), .B(n9036), .Z(n9063) );
  XNOR U9800 ( .A(n9064), .B(n9063), .Z(n9049) );
  NANDN U9801 ( .A(n9039), .B(n9038), .Z(n9043) );
  OR U9802 ( .A(n9041), .B(n9040), .Z(n9042) );
  NAND U9803 ( .A(n9043), .B(n9042), .Z(n9050) );
  XNOR U9804 ( .A(n9049), .B(n9050), .Z(n9051) );
  XOR U9805 ( .A(n9052), .B(n9051), .Z(n9048) );
  XNOR U9806 ( .A(sreg[1355]), .B(n9047), .Z(n9046) );
  XOR U9807 ( .A(n9048), .B(n9046), .Z(c[1355]) );
  NANDN U9808 ( .A(n9050), .B(n9049), .Z(n9054) );
  NAND U9809 ( .A(n9052), .B(n9051), .Z(n9053) );
  NAND U9810 ( .A(n9054), .B(n9053), .Z(n9070) );
  AND U9811 ( .A(b[2]), .B(a[334]), .Z(n9076) );
  AND U9812 ( .A(a[335]), .B(b[1]), .Z(n9074) );
  AND U9813 ( .A(a[333]), .B(b[3]), .Z(n9073) );
  XOR U9814 ( .A(n9074), .B(n9073), .Z(n9075) );
  XOR U9815 ( .A(n9076), .B(n9075), .Z(n9079) );
  NAND U9816 ( .A(b[0]), .B(a[336]), .Z(n9080) );
  XOR U9817 ( .A(n9079), .B(n9080), .Z(n9082) );
  OR U9818 ( .A(n9056), .B(n9055), .Z(n9060) );
  NANDN U9819 ( .A(n9058), .B(n9057), .Z(n9059) );
  NAND U9820 ( .A(n9060), .B(n9059), .Z(n9081) );
  XNOR U9821 ( .A(n9082), .B(n9081), .Z(n9067) );
  NANDN U9822 ( .A(n9062), .B(n9061), .Z(n9066) );
  OR U9823 ( .A(n9064), .B(n9063), .Z(n9065) );
  NAND U9824 ( .A(n9066), .B(n9065), .Z(n9068) );
  XNOR U9825 ( .A(n9067), .B(n9068), .Z(n9069) );
  XNOR U9826 ( .A(n9070), .B(n9069), .Z(n9085) );
  XNOR U9827 ( .A(n9085), .B(sreg[1356]), .Z(n9086) );
  XOR U9828 ( .A(n9087), .B(n9086), .Z(c[1356]) );
  NANDN U9829 ( .A(n9068), .B(n9067), .Z(n9072) );
  NAND U9830 ( .A(n9070), .B(n9069), .Z(n9071) );
  NAND U9831 ( .A(n9072), .B(n9071), .Z(n9094) );
  AND U9832 ( .A(b[2]), .B(a[335]), .Z(n9100) );
  AND U9833 ( .A(a[336]), .B(b[1]), .Z(n9098) );
  AND U9834 ( .A(a[334]), .B(b[3]), .Z(n9097) );
  XOR U9835 ( .A(n9098), .B(n9097), .Z(n9099) );
  XOR U9836 ( .A(n9100), .B(n9099), .Z(n9103) );
  NAND U9837 ( .A(b[0]), .B(a[337]), .Z(n9104) );
  XOR U9838 ( .A(n9103), .B(n9104), .Z(n9106) );
  OR U9839 ( .A(n9074), .B(n9073), .Z(n9078) );
  NANDN U9840 ( .A(n9076), .B(n9075), .Z(n9077) );
  NAND U9841 ( .A(n9078), .B(n9077), .Z(n9105) );
  XNOR U9842 ( .A(n9106), .B(n9105), .Z(n9091) );
  NANDN U9843 ( .A(n9080), .B(n9079), .Z(n9084) );
  OR U9844 ( .A(n9082), .B(n9081), .Z(n9083) );
  NAND U9845 ( .A(n9084), .B(n9083), .Z(n9092) );
  XNOR U9846 ( .A(n9091), .B(n9092), .Z(n9093) );
  XOR U9847 ( .A(n9094), .B(n9093), .Z(n9110) );
  NAND U9848 ( .A(n9085), .B(sreg[1356]), .Z(n9089) );
  OR U9849 ( .A(n9087), .B(n9086), .Z(n9088) );
  NAND U9850 ( .A(n9089), .B(n9088), .Z(n9109) );
  XNOR U9851 ( .A(sreg[1357]), .B(n9109), .Z(n9090) );
  XOR U9852 ( .A(n9110), .B(n9090), .Z(c[1357]) );
  NANDN U9853 ( .A(n9092), .B(n9091), .Z(n9096) );
  NAND U9854 ( .A(n9094), .B(n9093), .Z(n9095) );
  NAND U9855 ( .A(n9096), .B(n9095), .Z(n9117) );
  AND U9856 ( .A(b[2]), .B(a[336]), .Z(n9123) );
  AND U9857 ( .A(a[337]), .B(b[1]), .Z(n9121) );
  AND U9858 ( .A(a[335]), .B(b[3]), .Z(n9120) );
  XOR U9859 ( .A(n9121), .B(n9120), .Z(n9122) );
  XOR U9860 ( .A(n9123), .B(n9122), .Z(n9126) );
  NAND U9861 ( .A(b[0]), .B(a[338]), .Z(n9127) );
  XOR U9862 ( .A(n9126), .B(n9127), .Z(n9129) );
  OR U9863 ( .A(n9098), .B(n9097), .Z(n9102) );
  NANDN U9864 ( .A(n9100), .B(n9099), .Z(n9101) );
  NAND U9865 ( .A(n9102), .B(n9101), .Z(n9128) );
  XNOR U9866 ( .A(n9129), .B(n9128), .Z(n9114) );
  NANDN U9867 ( .A(n9104), .B(n9103), .Z(n9108) );
  OR U9868 ( .A(n9106), .B(n9105), .Z(n9107) );
  NAND U9869 ( .A(n9108), .B(n9107), .Z(n9115) );
  XNOR U9870 ( .A(n9114), .B(n9115), .Z(n9116) );
  XNOR U9871 ( .A(n9117), .B(n9116), .Z(n9113) );
  XOR U9872 ( .A(n9112), .B(sreg[1358]), .Z(n9111) );
  XOR U9873 ( .A(n9113), .B(n9111), .Z(c[1358]) );
  NANDN U9874 ( .A(n9115), .B(n9114), .Z(n9119) );
  NAND U9875 ( .A(n9117), .B(n9116), .Z(n9118) );
  NAND U9876 ( .A(n9119), .B(n9118), .Z(n9135) );
  AND U9877 ( .A(b[2]), .B(a[337]), .Z(n9141) );
  AND U9878 ( .A(a[338]), .B(b[1]), .Z(n9139) );
  AND U9879 ( .A(a[336]), .B(b[3]), .Z(n9138) );
  XOR U9880 ( .A(n9139), .B(n9138), .Z(n9140) );
  XOR U9881 ( .A(n9141), .B(n9140), .Z(n9144) );
  NAND U9882 ( .A(b[0]), .B(a[339]), .Z(n9145) );
  XOR U9883 ( .A(n9144), .B(n9145), .Z(n9147) );
  OR U9884 ( .A(n9121), .B(n9120), .Z(n9125) );
  NANDN U9885 ( .A(n9123), .B(n9122), .Z(n9124) );
  NAND U9886 ( .A(n9125), .B(n9124), .Z(n9146) );
  XNOR U9887 ( .A(n9147), .B(n9146), .Z(n9132) );
  NANDN U9888 ( .A(n9127), .B(n9126), .Z(n9131) );
  OR U9889 ( .A(n9129), .B(n9128), .Z(n9130) );
  NAND U9890 ( .A(n9131), .B(n9130), .Z(n9133) );
  XNOR U9891 ( .A(n9132), .B(n9133), .Z(n9134) );
  XNOR U9892 ( .A(n9135), .B(n9134), .Z(n9150) );
  XNOR U9893 ( .A(n9150), .B(sreg[1359]), .Z(n9152) );
  XNOR U9894 ( .A(n9151), .B(n9152), .Z(c[1359]) );
  NANDN U9895 ( .A(n9133), .B(n9132), .Z(n9137) );
  NAND U9896 ( .A(n9135), .B(n9134), .Z(n9136) );
  NAND U9897 ( .A(n9137), .B(n9136), .Z(n9161) );
  AND U9898 ( .A(b[2]), .B(a[338]), .Z(n9173) );
  AND U9899 ( .A(a[339]), .B(b[1]), .Z(n9171) );
  AND U9900 ( .A(a[337]), .B(b[3]), .Z(n9170) );
  XOR U9901 ( .A(n9171), .B(n9170), .Z(n9172) );
  XOR U9902 ( .A(n9173), .B(n9172), .Z(n9164) );
  NAND U9903 ( .A(b[0]), .B(a[340]), .Z(n9165) );
  XOR U9904 ( .A(n9164), .B(n9165), .Z(n9167) );
  OR U9905 ( .A(n9139), .B(n9138), .Z(n9143) );
  NANDN U9906 ( .A(n9141), .B(n9140), .Z(n9142) );
  NAND U9907 ( .A(n9143), .B(n9142), .Z(n9166) );
  XNOR U9908 ( .A(n9167), .B(n9166), .Z(n9158) );
  NANDN U9909 ( .A(n9145), .B(n9144), .Z(n9149) );
  OR U9910 ( .A(n9147), .B(n9146), .Z(n9148) );
  NAND U9911 ( .A(n9149), .B(n9148), .Z(n9159) );
  XNOR U9912 ( .A(n9158), .B(n9159), .Z(n9160) );
  XOR U9913 ( .A(n9161), .B(n9160), .Z(n9157) );
  NAND U9914 ( .A(n9150), .B(sreg[1359]), .Z(n9154) );
  NANDN U9915 ( .A(n9152), .B(n9151), .Z(n9153) );
  NAND U9916 ( .A(n9154), .B(n9153), .Z(n9156) );
  XNOR U9917 ( .A(sreg[1360]), .B(n9156), .Z(n9155) );
  XOR U9918 ( .A(n9157), .B(n9155), .Z(c[1360]) );
  NANDN U9919 ( .A(n9159), .B(n9158), .Z(n9163) );
  NAND U9920 ( .A(n9161), .B(n9160), .Z(n9162) );
  NAND U9921 ( .A(n9163), .B(n9162), .Z(n9191) );
  NANDN U9922 ( .A(n9165), .B(n9164), .Z(n9169) );
  OR U9923 ( .A(n9167), .B(n9166), .Z(n9168) );
  NAND U9924 ( .A(n9169), .B(n9168), .Z(n9188) );
  AND U9925 ( .A(b[2]), .B(a[339]), .Z(n9179) );
  AND U9926 ( .A(a[340]), .B(b[1]), .Z(n9177) );
  AND U9927 ( .A(a[338]), .B(b[3]), .Z(n9176) );
  XOR U9928 ( .A(n9177), .B(n9176), .Z(n9178) );
  XOR U9929 ( .A(n9179), .B(n9178), .Z(n9182) );
  NAND U9930 ( .A(b[0]), .B(a[341]), .Z(n9183) );
  XNOR U9931 ( .A(n9182), .B(n9183), .Z(n9184) );
  OR U9932 ( .A(n9171), .B(n9170), .Z(n9175) );
  NANDN U9933 ( .A(n9173), .B(n9172), .Z(n9174) );
  AND U9934 ( .A(n9175), .B(n9174), .Z(n9185) );
  XNOR U9935 ( .A(n9184), .B(n9185), .Z(n9189) );
  XNOR U9936 ( .A(n9188), .B(n9189), .Z(n9190) );
  XNOR U9937 ( .A(n9191), .B(n9190), .Z(n9194) );
  XNOR U9938 ( .A(sreg[1361]), .B(n9194), .Z(n9195) );
  XOR U9939 ( .A(n9196), .B(n9195), .Z(c[1361]) );
  AND U9940 ( .A(b[2]), .B(a[340]), .Z(n9209) );
  AND U9941 ( .A(a[341]), .B(b[1]), .Z(n9207) );
  AND U9942 ( .A(a[339]), .B(b[3]), .Z(n9206) );
  XOR U9943 ( .A(n9207), .B(n9206), .Z(n9208) );
  XOR U9944 ( .A(n9209), .B(n9208), .Z(n9212) );
  NAND U9945 ( .A(b[0]), .B(a[342]), .Z(n9213) );
  XOR U9946 ( .A(n9212), .B(n9213), .Z(n9215) );
  OR U9947 ( .A(n9177), .B(n9176), .Z(n9181) );
  NANDN U9948 ( .A(n9179), .B(n9178), .Z(n9180) );
  NAND U9949 ( .A(n9181), .B(n9180), .Z(n9214) );
  XNOR U9950 ( .A(n9215), .B(n9214), .Z(n9200) );
  NANDN U9951 ( .A(n9183), .B(n9182), .Z(n9187) );
  NAND U9952 ( .A(n9185), .B(n9184), .Z(n9186) );
  NAND U9953 ( .A(n9187), .B(n9186), .Z(n9201) );
  XNOR U9954 ( .A(n9200), .B(n9201), .Z(n9202) );
  NANDN U9955 ( .A(n9189), .B(n9188), .Z(n9193) );
  NANDN U9956 ( .A(n9191), .B(n9190), .Z(n9192) );
  NAND U9957 ( .A(n9193), .B(n9192), .Z(n9203) );
  XOR U9958 ( .A(n9202), .B(n9203), .Z(n9219) );
  NAND U9959 ( .A(sreg[1361]), .B(n9194), .Z(n9198) );
  OR U9960 ( .A(n9196), .B(n9195), .Z(n9197) );
  NAND U9961 ( .A(n9198), .B(n9197), .Z(n9218) );
  XNOR U9962 ( .A(sreg[1362]), .B(n9218), .Z(n9199) );
  XNOR U9963 ( .A(n9219), .B(n9199), .Z(c[1362]) );
  NANDN U9964 ( .A(n9201), .B(n9200), .Z(n9205) );
  NANDN U9965 ( .A(n9203), .B(n9202), .Z(n9204) );
  NAND U9966 ( .A(n9205), .B(n9204), .Z(n9236) );
  AND U9967 ( .A(b[2]), .B(a[341]), .Z(n9230) );
  AND U9968 ( .A(a[342]), .B(b[1]), .Z(n9228) );
  AND U9969 ( .A(a[340]), .B(b[3]), .Z(n9227) );
  XOR U9970 ( .A(n9228), .B(n9227), .Z(n9229) );
  XOR U9971 ( .A(n9230), .B(n9229), .Z(n9221) );
  NAND U9972 ( .A(b[0]), .B(a[343]), .Z(n9222) );
  XOR U9973 ( .A(n9221), .B(n9222), .Z(n9224) );
  OR U9974 ( .A(n9207), .B(n9206), .Z(n9211) );
  NANDN U9975 ( .A(n9209), .B(n9208), .Z(n9210) );
  NAND U9976 ( .A(n9211), .B(n9210), .Z(n9223) );
  XNOR U9977 ( .A(n9224), .B(n9223), .Z(n9233) );
  NANDN U9978 ( .A(n9213), .B(n9212), .Z(n9217) );
  OR U9979 ( .A(n9215), .B(n9214), .Z(n9216) );
  NAND U9980 ( .A(n9217), .B(n9216), .Z(n9234) );
  XNOR U9981 ( .A(n9233), .B(n9234), .Z(n9235) );
  XNOR U9982 ( .A(n9236), .B(n9235), .Z(n9240) );
  XOR U9983 ( .A(n9239), .B(sreg[1363]), .Z(n9220) );
  XOR U9984 ( .A(n9240), .B(n9220), .Z(c[1363]) );
  NANDN U9985 ( .A(n9222), .B(n9221), .Z(n9226) );
  OR U9986 ( .A(n9224), .B(n9223), .Z(n9225) );
  NAND U9987 ( .A(n9226), .B(n9225), .Z(n9256) );
  AND U9988 ( .A(b[2]), .B(a[342]), .Z(n9247) );
  AND U9989 ( .A(a[343]), .B(b[1]), .Z(n9245) );
  AND U9990 ( .A(a[341]), .B(b[3]), .Z(n9244) );
  XOR U9991 ( .A(n9245), .B(n9244), .Z(n9246) );
  XOR U9992 ( .A(n9247), .B(n9246), .Z(n9250) );
  NAND U9993 ( .A(b[0]), .B(a[344]), .Z(n9251) );
  XNOR U9994 ( .A(n9250), .B(n9251), .Z(n9252) );
  OR U9995 ( .A(n9228), .B(n9227), .Z(n9232) );
  NANDN U9996 ( .A(n9230), .B(n9229), .Z(n9231) );
  AND U9997 ( .A(n9232), .B(n9231), .Z(n9253) );
  XNOR U9998 ( .A(n9252), .B(n9253), .Z(n9257) );
  XNOR U9999 ( .A(n9256), .B(n9257), .Z(n9258) );
  NANDN U10000 ( .A(n9234), .B(n9233), .Z(n9238) );
  NAND U10001 ( .A(n9236), .B(n9235), .Z(n9237) );
  AND U10002 ( .A(n9238), .B(n9237), .Z(n9259) );
  XNOR U10003 ( .A(n9258), .B(n9259), .Z(n9243) );
  XOR U10004 ( .A(sreg[1364]), .B(n9242), .Z(n9241) );
  XOR U10005 ( .A(n9243), .B(n9241), .Z(c[1364]) );
  AND U10006 ( .A(b[2]), .B(a[343]), .Z(n9271) );
  AND U10007 ( .A(a[344]), .B(b[1]), .Z(n9269) );
  AND U10008 ( .A(a[342]), .B(b[3]), .Z(n9268) );
  XOR U10009 ( .A(n9269), .B(n9268), .Z(n9270) );
  XOR U10010 ( .A(n9271), .B(n9270), .Z(n9274) );
  NAND U10011 ( .A(b[0]), .B(a[345]), .Z(n9275) );
  XOR U10012 ( .A(n9274), .B(n9275), .Z(n9277) );
  OR U10013 ( .A(n9245), .B(n9244), .Z(n9249) );
  NANDN U10014 ( .A(n9247), .B(n9246), .Z(n9248) );
  NAND U10015 ( .A(n9249), .B(n9248), .Z(n9276) );
  XNOR U10016 ( .A(n9277), .B(n9276), .Z(n9262) );
  NANDN U10017 ( .A(n9251), .B(n9250), .Z(n9255) );
  NAND U10018 ( .A(n9253), .B(n9252), .Z(n9254) );
  NAND U10019 ( .A(n9255), .B(n9254), .Z(n9263) );
  XNOR U10020 ( .A(n9262), .B(n9263), .Z(n9264) );
  NANDN U10021 ( .A(n9257), .B(n9256), .Z(n9261) );
  NAND U10022 ( .A(n9259), .B(n9258), .Z(n9260) );
  NAND U10023 ( .A(n9261), .B(n9260), .Z(n9265) );
  XOR U10024 ( .A(n9264), .B(n9265), .Z(n9280) );
  XNOR U10025 ( .A(n9280), .B(sreg[1365]), .Z(n9281) );
  XOR U10026 ( .A(n9282), .B(n9281), .Z(c[1365]) );
  NANDN U10027 ( .A(n9263), .B(n9262), .Z(n9267) );
  NANDN U10028 ( .A(n9265), .B(n9264), .Z(n9266) );
  NAND U10029 ( .A(n9267), .B(n9266), .Z(n9300) );
  AND U10030 ( .A(b[2]), .B(a[344]), .Z(n9294) );
  AND U10031 ( .A(a[345]), .B(b[1]), .Z(n9292) );
  AND U10032 ( .A(a[343]), .B(b[3]), .Z(n9291) );
  XOR U10033 ( .A(n9292), .B(n9291), .Z(n9293) );
  XOR U10034 ( .A(n9294), .B(n9293), .Z(n9285) );
  NAND U10035 ( .A(b[0]), .B(a[346]), .Z(n9286) );
  XOR U10036 ( .A(n9285), .B(n9286), .Z(n9288) );
  OR U10037 ( .A(n9269), .B(n9268), .Z(n9273) );
  NANDN U10038 ( .A(n9271), .B(n9270), .Z(n9272) );
  NAND U10039 ( .A(n9273), .B(n9272), .Z(n9287) );
  XNOR U10040 ( .A(n9288), .B(n9287), .Z(n9297) );
  NANDN U10041 ( .A(n9275), .B(n9274), .Z(n9279) );
  OR U10042 ( .A(n9277), .B(n9276), .Z(n9278) );
  NAND U10043 ( .A(n9279), .B(n9278), .Z(n9298) );
  XNOR U10044 ( .A(n9297), .B(n9298), .Z(n9299) );
  XNOR U10045 ( .A(n9300), .B(n9299), .Z(n9303) );
  XOR U10046 ( .A(sreg[1366]), .B(n9303), .Z(n9304) );
  NAND U10047 ( .A(n9280), .B(sreg[1365]), .Z(n9284) );
  OR U10048 ( .A(n9282), .B(n9281), .Z(n9283) );
  NAND U10049 ( .A(n9284), .B(n9283), .Z(n9305) );
  XOR U10050 ( .A(n9304), .B(n9305), .Z(c[1366]) );
  NANDN U10051 ( .A(n9286), .B(n9285), .Z(n9290) );
  OR U10052 ( .A(n9288), .B(n9287), .Z(n9289) );
  NAND U10053 ( .A(n9290), .B(n9289), .Z(n9309) );
  AND U10054 ( .A(b[2]), .B(a[345]), .Z(n9318) );
  AND U10055 ( .A(a[346]), .B(b[1]), .Z(n9316) );
  AND U10056 ( .A(a[344]), .B(b[3]), .Z(n9315) );
  XOR U10057 ( .A(n9316), .B(n9315), .Z(n9317) );
  XOR U10058 ( .A(n9318), .B(n9317), .Z(n9321) );
  NAND U10059 ( .A(b[0]), .B(a[347]), .Z(n9322) );
  XNOR U10060 ( .A(n9321), .B(n9322), .Z(n9323) );
  OR U10061 ( .A(n9292), .B(n9291), .Z(n9296) );
  NANDN U10062 ( .A(n9294), .B(n9293), .Z(n9295) );
  AND U10063 ( .A(n9296), .B(n9295), .Z(n9324) );
  XNOR U10064 ( .A(n9323), .B(n9324), .Z(n9310) );
  XNOR U10065 ( .A(n9309), .B(n9310), .Z(n9311) );
  NANDN U10066 ( .A(n9298), .B(n9297), .Z(n9302) );
  NAND U10067 ( .A(n9300), .B(n9299), .Z(n9301) );
  AND U10068 ( .A(n9302), .B(n9301), .Z(n9312) );
  XNOR U10069 ( .A(n9311), .B(n9312), .Z(n9328) );
  OR U10070 ( .A(n9303), .B(sreg[1366]), .Z(n9307) );
  NANDN U10071 ( .A(n9305), .B(n9304), .Z(n9306) );
  AND U10072 ( .A(n9307), .B(n9306), .Z(n9327) );
  XNOR U10073 ( .A(sreg[1367]), .B(n9327), .Z(n9308) );
  XOR U10074 ( .A(n9328), .B(n9308), .Z(c[1367]) );
  NANDN U10075 ( .A(n9310), .B(n9309), .Z(n9314) );
  NAND U10076 ( .A(n9312), .B(n9311), .Z(n9313) );
  NAND U10077 ( .A(n9314), .B(n9313), .Z(n9335) );
  AND U10078 ( .A(b[2]), .B(a[346]), .Z(n9341) );
  AND U10079 ( .A(a[347]), .B(b[1]), .Z(n9339) );
  AND U10080 ( .A(a[345]), .B(b[3]), .Z(n9338) );
  XOR U10081 ( .A(n9339), .B(n9338), .Z(n9340) );
  XOR U10082 ( .A(n9341), .B(n9340), .Z(n9344) );
  NAND U10083 ( .A(b[0]), .B(a[348]), .Z(n9345) );
  XOR U10084 ( .A(n9344), .B(n9345), .Z(n9347) );
  OR U10085 ( .A(n9316), .B(n9315), .Z(n9320) );
  NANDN U10086 ( .A(n9318), .B(n9317), .Z(n9319) );
  NAND U10087 ( .A(n9320), .B(n9319), .Z(n9346) );
  XNOR U10088 ( .A(n9347), .B(n9346), .Z(n9332) );
  NANDN U10089 ( .A(n9322), .B(n9321), .Z(n9326) );
  NAND U10090 ( .A(n9324), .B(n9323), .Z(n9325) );
  NAND U10091 ( .A(n9326), .B(n9325), .Z(n9333) );
  XNOR U10092 ( .A(n9332), .B(n9333), .Z(n9334) );
  XNOR U10093 ( .A(n9335), .B(n9334), .Z(n9331) );
  XOR U10094 ( .A(n9330), .B(sreg[1368]), .Z(n9329) );
  XNOR U10095 ( .A(n9331), .B(n9329), .Z(c[1368]) );
  NANDN U10096 ( .A(n9333), .B(n9332), .Z(n9337) );
  NANDN U10097 ( .A(n9335), .B(n9334), .Z(n9336) );
  NAND U10098 ( .A(n9337), .B(n9336), .Z(n9370) );
  AND U10099 ( .A(b[2]), .B(a[347]), .Z(n9364) );
  AND U10100 ( .A(a[348]), .B(b[1]), .Z(n9362) );
  AND U10101 ( .A(a[346]), .B(b[3]), .Z(n9361) );
  XOR U10102 ( .A(n9362), .B(n9361), .Z(n9363) );
  XOR U10103 ( .A(n9364), .B(n9363), .Z(n9355) );
  NAND U10104 ( .A(b[0]), .B(a[349]), .Z(n9356) );
  XOR U10105 ( .A(n9355), .B(n9356), .Z(n9358) );
  OR U10106 ( .A(n9339), .B(n9338), .Z(n9343) );
  NANDN U10107 ( .A(n9341), .B(n9340), .Z(n9342) );
  NAND U10108 ( .A(n9343), .B(n9342), .Z(n9357) );
  XNOR U10109 ( .A(n9358), .B(n9357), .Z(n9367) );
  NANDN U10110 ( .A(n9345), .B(n9344), .Z(n9349) );
  OR U10111 ( .A(n9347), .B(n9346), .Z(n9348) );
  NAND U10112 ( .A(n9349), .B(n9348), .Z(n9368) );
  XNOR U10113 ( .A(n9367), .B(n9368), .Z(n9369) );
  XNOR U10114 ( .A(n9370), .B(n9369), .Z(n9350) );
  XNOR U10115 ( .A(n9350), .B(sreg[1369]), .Z(n9352) );
  XNOR U10116 ( .A(n9351), .B(n9352), .Z(c[1369]) );
  NAND U10117 ( .A(n9350), .B(sreg[1369]), .Z(n9354) );
  NANDN U10118 ( .A(n9352), .B(n9351), .Z(n9353) );
  NAND U10119 ( .A(n9354), .B(n9353), .Z(n9374) );
  NANDN U10120 ( .A(n9356), .B(n9355), .Z(n9360) );
  OR U10121 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U10122 ( .A(n9360), .B(n9359), .Z(n9376) );
  AND U10123 ( .A(b[2]), .B(a[348]), .Z(n9385) );
  AND U10124 ( .A(a[349]), .B(b[1]), .Z(n9383) );
  AND U10125 ( .A(a[347]), .B(b[3]), .Z(n9382) );
  XOR U10126 ( .A(n9383), .B(n9382), .Z(n9384) );
  XOR U10127 ( .A(n9385), .B(n9384), .Z(n9388) );
  NAND U10128 ( .A(b[0]), .B(a[350]), .Z(n9389) );
  XNOR U10129 ( .A(n9388), .B(n9389), .Z(n9390) );
  OR U10130 ( .A(n9362), .B(n9361), .Z(n9366) );
  NANDN U10131 ( .A(n9364), .B(n9363), .Z(n9365) );
  AND U10132 ( .A(n9366), .B(n9365), .Z(n9391) );
  XNOR U10133 ( .A(n9390), .B(n9391), .Z(n9377) );
  XNOR U10134 ( .A(n9376), .B(n9377), .Z(n9378) );
  NANDN U10135 ( .A(n9368), .B(n9367), .Z(n9372) );
  NAND U10136 ( .A(n9370), .B(n9369), .Z(n9371) );
  AND U10137 ( .A(n9372), .B(n9371), .Z(n9379) );
  XNOR U10138 ( .A(n9378), .B(n9379), .Z(n9375) );
  XOR U10139 ( .A(sreg[1370]), .B(n9375), .Z(n9373) );
  XNOR U10140 ( .A(n9374), .B(n9373), .Z(c[1370]) );
  NANDN U10141 ( .A(n9377), .B(n9376), .Z(n9381) );
  NAND U10142 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND U10143 ( .A(n9381), .B(n9380), .Z(n9397) );
  AND U10144 ( .A(b[2]), .B(a[349]), .Z(n9403) );
  AND U10145 ( .A(a[350]), .B(b[1]), .Z(n9401) );
  AND U10146 ( .A(a[348]), .B(b[3]), .Z(n9400) );
  XOR U10147 ( .A(n9401), .B(n9400), .Z(n9402) );
  XOR U10148 ( .A(n9403), .B(n9402), .Z(n9406) );
  NAND U10149 ( .A(b[0]), .B(a[351]), .Z(n9407) );
  XOR U10150 ( .A(n9406), .B(n9407), .Z(n9409) );
  OR U10151 ( .A(n9383), .B(n9382), .Z(n9387) );
  NANDN U10152 ( .A(n9385), .B(n9384), .Z(n9386) );
  NAND U10153 ( .A(n9387), .B(n9386), .Z(n9408) );
  XNOR U10154 ( .A(n9409), .B(n9408), .Z(n9394) );
  NANDN U10155 ( .A(n9389), .B(n9388), .Z(n9393) );
  NAND U10156 ( .A(n9391), .B(n9390), .Z(n9392) );
  NAND U10157 ( .A(n9393), .B(n9392), .Z(n9395) );
  XNOR U10158 ( .A(n9394), .B(n9395), .Z(n9396) );
  XOR U10159 ( .A(n9397), .B(n9396), .Z(n9412) );
  XNOR U10160 ( .A(n9412), .B(sreg[1371]), .Z(n9413) );
  XOR U10161 ( .A(n9414), .B(n9413), .Z(c[1371]) );
  NANDN U10162 ( .A(n9395), .B(n9394), .Z(n9399) );
  NANDN U10163 ( .A(n9397), .B(n9396), .Z(n9398) );
  NAND U10164 ( .A(n9399), .B(n9398), .Z(n9432) );
  AND U10165 ( .A(b[2]), .B(a[350]), .Z(n9426) );
  AND U10166 ( .A(a[351]), .B(b[1]), .Z(n9424) );
  AND U10167 ( .A(a[349]), .B(b[3]), .Z(n9423) );
  XOR U10168 ( .A(n9424), .B(n9423), .Z(n9425) );
  XOR U10169 ( .A(n9426), .B(n9425), .Z(n9417) );
  NAND U10170 ( .A(b[0]), .B(a[352]), .Z(n9418) );
  XOR U10171 ( .A(n9417), .B(n9418), .Z(n9420) );
  OR U10172 ( .A(n9401), .B(n9400), .Z(n9405) );
  NANDN U10173 ( .A(n9403), .B(n9402), .Z(n9404) );
  NAND U10174 ( .A(n9405), .B(n9404), .Z(n9419) );
  XNOR U10175 ( .A(n9420), .B(n9419), .Z(n9429) );
  NANDN U10176 ( .A(n9407), .B(n9406), .Z(n9411) );
  OR U10177 ( .A(n9409), .B(n9408), .Z(n9410) );
  NAND U10178 ( .A(n9411), .B(n9410), .Z(n9430) );
  XNOR U10179 ( .A(n9429), .B(n9430), .Z(n9431) );
  XNOR U10180 ( .A(n9432), .B(n9431), .Z(n9435) );
  XOR U10181 ( .A(sreg[1372]), .B(n9435), .Z(n9436) );
  NAND U10182 ( .A(n9412), .B(sreg[1371]), .Z(n9416) );
  OR U10183 ( .A(n9414), .B(n9413), .Z(n9415) );
  NAND U10184 ( .A(n9416), .B(n9415), .Z(n9437) );
  XOR U10185 ( .A(n9436), .B(n9437), .Z(c[1372]) );
  NANDN U10186 ( .A(n9418), .B(n9417), .Z(n9422) );
  OR U10187 ( .A(n9420), .B(n9419), .Z(n9421) );
  NAND U10188 ( .A(n9422), .B(n9421), .Z(n9441) );
  AND U10189 ( .A(b[2]), .B(a[351]), .Z(n9450) );
  AND U10190 ( .A(a[352]), .B(b[1]), .Z(n9448) );
  AND U10191 ( .A(a[350]), .B(b[3]), .Z(n9447) );
  XOR U10192 ( .A(n9448), .B(n9447), .Z(n9449) );
  XOR U10193 ( .A(n9450), .B(n9449), .Z(n9453) );
  NAND U10194 ( .A(b[0]), .B(a[353]), .Z(n9454) );
  XNOR U10195 ( .A(n9453), .B(n9454), .Z(n9455) );
  OR U10196 ( .A(n9424), .B(n9423), .Z(n9428) );
  NANDN U10197 ( .A(n9426), .B(n9425), .Z(n9427) );
  AND U10198 ( .A(n9428), .B(n9427), .Z(n9456) );
  XNOR U10199 ( .A(n9455), .B(n9456), .Z(n9442) );
  XNOR U10200 ( .A(n9441), .B(n9442), .Z(n9443) );
  NANDN U10201 ( .A(n9430), .B(n9429), .Z(n9434) );
  NAND U10202 ( .A(n9432), .B(n9431), .Z(n9433) );
  AND U10203 ( .A(n9434), .B(n9433), .Z(n9444) );
  XNOR U10204 ( .A(n9443), .B(n9444), .Z(n9460) );
  OR U10205 ( .A(n9435), .B(sreg[1372]), .Z(n9439) );
  NANDN U10206 ( .A(n9437), .B(n9436), .Z(n9438) );
  AND U10207 ( .A(n9439), .B(n9438), .Z(n9459) );
  XNOR U10208 ( .A(sreg[1373]), .B(n9459), .Z(n9440) );
  XOR U10209 ( .A(n9460), .B(n9440), .Z(c[1373]) );
  NANDN U10210 ( .A(n9442), .B(n9441), .Z(n9446) );
  NAND U10211 ( .A(n9444), .B(n9443), .Z(n9445) );
  NAND U10212 ( .A(n9446), .B(n9445), .Z(n9465) );
  AND U10213 ( .A(b[2]), .B(a[352]), .Z(n9471) );
  AND U10214 ( .A(a[353]), .B(b[1]), .Z(n9469) );
  AND U10215 ( .A(a[351]), .B(b[3]), .Z(n9468) );
  XOR U10216 ( .A(n9469), .B(n9468), .Z(n9470) );
  XOR U10217 ( .A(n9471), .B(n9470), .Z(n9474) );
  NAND U10218 ( .A(b[0]), .B(a[354]), .Z(n9475) );
  XOR U10219 ( .A(n9474), .B(n9475), .Z(n9477) );
  OR U10220 ( .A(n9448), .B(n9447), .Z(n9452) );
  NANDN U10221 ( .A(n9450), .B(n9449), .Z(n9451) );
  NAND U10222 ( .A(n9452), .B(n9451), .Z(n9476) );
  XNOR U10223 ( .A(n9477), .B(n9476), .Z(n9462) );
  NANDN U10224 ( .A(n9454), .B(n9453), .Z(n9458) );
  NAND U10225 ( .A(n9456), .B(n9455), .Z(n9457) );
  NAND U10226 ( .A(n9458), .B(n9457), .Z(n9463) );
  XNOR U10227 ( .A(n9462), .B(n9463), .Z(n9464) );
  XNOR U10228 ( .A(n9465), .B(n9464), .Z(n9481) );
  XOR U10229 ( .A(n9480), .B(sreg[1374]), .Z(n9461) );
  XNOR U10230 ( .A(n9481), .B(n9461), .Z(c[1374]) );
  NANDN U10231 ( .A(n9463), .B(n9462), .Z(n9467) );
  NANDN U10232 ( .A(n9465), .B(n9464), .Z(n9466) );
  NAND U10233 ( .A(n9467), .B(n9466), .Z(n9486) );
  AND U10234 ( .A(b[2]), .B(a[353]), .Z(n9492) );
  AND U10235 ( .A(a[354]), .B(b[1]), .Z(n9490) );
  AND U10236 ( .A(a[352]), .B(b[3]), .Z(n9489) );
  XOR U10237 ( .A(n9490), .B(n9489), .Z(n9491) );
  XOR U10238 ( .A(n9492), .B(n9491), .Z(n9495) );
  NAND U10239 ( .A(b[0]), .B(a[355]), .Z(n9496) );
  XOR U10240 ( .A(n9495), .B(n9496), .Z(n9498) );
  OR U10241 ( .A(n9469), .B(n9468), .Z(n9473) );
  NANDN U10242 ( .A(n9471), .B(n9470), .Z(n9472) );
  NAND U10243 ( .A(n9473), .B(n9472), .Z(n9497) );
  XNOR U10244 ( .A(n9498), .B(n9497), .Z(n9483) );
  NANDN U10245 ( .A(n9475), .B(n9474), .Z(n9479) );
  OR U10246 ( .A(n9477), .B(n9476), .Z(n9478) );
  NAND U10247 ( .A(n9479), .B(n9478), .Z(n9484) );
  XNOR U10248 ( .A(n9483), .B(n9484), .Z(n9485) );
  XNOR U10249 ( .A(n9486), .B(n9485), .Z(n9502) );
  XNOR U10250 ( .A(sreg[1375]), .B(n9503), .Z(n9482) );
  XNOR U10251 ( .A(n9502), .B(n9482), .Z(c[1375]) );
  NANDN U10252 ( .A(n9484), .B(n9483), .Z(n9488) );
  NAND U10253 ( .A(n9486), .B(n9485), .Z(n9487) );
  NAND U10254 ( .A(n9488), .B(n9487), .Z(n9509) );
  AND U10255 ( .A(b[2]), .B(a[354]), .Z(n9513) );
  AND U10256 ( .A(a[355]), .B(b[1]), .Z(n9511) );
  AND U10257 ( .A(a[353]), .B(b[3]), .Z(n9510) );
  XOR U10258 ( .A(n9511), .B(n9510), .Z(n9512) );
  XOR U10259 ( .A(n9513), .B(n9512), .Z(n9516) );
  NAND U10260 ( .A(b[0]), .B(a[356]), .Z(n9517) );
  XOR U10261 ( .A(n9516), .B(n9517), .Z(n9518) );
  OR U10262 ( .A(n9490), .B(n9489), .Z(n9494) );
  NANDN U10263 ( .A(n9492), .B(n9491), .Z(n9493) );
  AND U10264 ( .A(n9494), .B(n9493), .Z(n9519) );
  XOR U10265 ( .A(n9518), .B(n9519), .Z(n9507) );
  NANDN U10266 ( .A(n9496), .B(n9495), .Z(n9500) );
  OR U10267 ( .A(n9498), .B(n9497), .Z(n9499) );
  AND U10268 ( .A(n9500), .B(n9499), .Z(n9508) );
  XOR U10269 ( .A(n9507), .B(n9508), .Z(n9501) );
  XOR U10270 ( .A(n9509), .B(n9501), .Z(n9506) );
  XOR U10271 ( .A(n9505), .B(sreg[1376]), .Z(n9504) );
  XNOR U10272 ( .A(n9506), .B(n9504), .Z(c[1376]) );
  AND U10273 ( .A(b[2]), .B(a[355]), .Z(n9529) );
  AND U10274 ( .A(a[356]), .B(b[1]), .Z(n9527) );
  AND U10275 ( .A(a[354]), .B(b[3]), .Z(n9526) );
  XOR U10276 ( .A(n9527), .B(n9526), .Z(n9528) );
  XOR U10277 ( .A(n9529), .B(n9528), .Z(n9532) );
  NAND U10278 ( .A(b[0]), .B(a[357]), .Z(n9533) );
  XOR U10279 ( .A(n9532), .B(n9533), .Z(n9535) );
  OR U10280 ( .A(n9511), .B(n9510), .Z(n9515) );
  NANDN U10281 ( .A(n9513), .B(n9512), .Z(n9514) );
  NAND U10282 ( .A(n9515), .B(n9514), .Z(n9534) );
  XNOR U10283 ( .A(n9535), .B(n9534), .Z(n9520) );
  XNOR U10284 ( .A(n9520), .B(n9521), .Z(n9523) );
  XOR U10285 ( .A(n9522), .B(n9523), .Z(n9538) );
  XOR U10286 ( .A(n9538), .B(sreg[1377]), .Z(n9540) );
  XNOR U10287 ( .A(n9539), .B(n9540), .Z(c[1377]) );
  NANDN U10288 ( .A(n9521), .B(n9520), .Z(n9525) );
  NAND U10289 ( .A(n9523), .B(n9522), .Z(n9524) );
  NAND U10290 ( .A(n9525), .B(n9524), .Z(n9547) );
  AND U10291 ( .A(b[2]), .B(a[356]), .Z(n9553) );
  AND U10292 ( .A(a[357]), .B(b[1]), .Z(n9551) );
  AND U10293 ( .A(a[355]), .B(b[3]), .Z(n9550) );
  XOR U10294 ( .A(n9551), .B(n9550), .Z(n9552) );
  XOR U10295 ( .A(n9553), .B(n9552), .Z(n9556) );
  NAND U10296 ( .A(b[0]), .B(a[358]), .Z(n9557) );
  XOR U10297 ( .A(n9556), .B(n9557), .Z(n9559) );
  OR U10298 ( .A(n9527), .B(n9526), .Z(n9531) );
  NANDN U10299 ( .A(n9529), .B(n9528), .Z(n9530) );
  NAND U10300 ( .A(n9531), .B(n9530), .Z(n9558) );
  XNOR U10301 ( .A(n9559), .B(n9558), .Z(n9544) );
  NANDN U10302 ( .A(n9533), .B(n9532), .Z(n9537) );
  OR U10303 ( .A(n9535), .B(n9534), .Z(n9536) );
  NAND U10304 ( .A(n9537), .B(n9536), .Z(n9545) );
  XNOR U10305 ( .A(n9544), .B(n9545), .Z(n9546) );
  XOR U10306 ( .A(n9547), .B(n9546), .Z(n9563) );
  NANDN U10307 ( .A(n9538), .B(sreg[1377]), .Z(n9542) );
  NANDN U10308 ( .A(n9540), .B(n9539), .Z(n9541) );
  NAND U10309 ( .A(n9542), .B(n9541), .Z(n9562) );
  XNOR U10310 ( .A(sreg[1378]), .B(n9562), .Z(n9543) );
  XOR U10311 ( .A(n9563), .B(n9543), .Z(c[1378]) );
  NANDN U10312 ( .A(n9545), .B(n9544), .Z(n9549) );
  NAND U10313 ( .A(n9547), .B(n9546), .Z(n9548) );
  NAND U10314 ( .A(n9549), .B(n9548), .Z(n9568) );
  AND U10315 ( .A(b[2]), .B(a[357]), .Z(n9574) );
  AND U10316 ( .A(a[358]), .B(b[1]), .Z(n9572) );
  AND U10317 ( .A(a[356]), .B(b[3]), .Z(n9571) );
  XOR U10318 ( .A(n9572), .B(n9571), .Z(n9573) );
  XOR U10319 ( .A(n9574), .B(n9573), .Z(n9577) );
  NAND U10320 ( .A(b[0]), .B(a[359]), .Z(n9578) );
  XOR U10321 ( .A(n9577), .B(n9578), .Z(n9580) );
  OR U10322 ( .A(n9551), .B(n9550), .Z(n9555) );
  NANDN U10323 ( .A(n9553), .B(n9552), .Z(n9554) );
  NAND U10324 ( .A(n9555), .B(n9554), .Z(n9579) );
  XNOR U10325 ( .A(n9580), .B(n9579), .Z(n9565) );
  NANDN U10326 ( .A(n9557), .B(n9556), .Z(n9561) );
  OR U10327 ( .A(n9559), .B(n9558), .Z(n9560) );
  NAND U10328 ( .A(n9561), .B(n9560), .Z(n9566) );
  XNOR U10329 ( .A(n9565), .B(n9566), .Z(n9567) );
  XNOR U10330 ( .A(n9568), .B(n9567), .Z(n9584) );
  XOR U10331 ( .A(n9583), .B(sreg[1379]), .Z(n9564) );
  XOR U10332 ( .A(n9584), .B(n9564), .Z(c[1379]) );
  NANDN U10333 ( .A(n9566), .B(n9565), .Z(n9570) );
  NAND U10334 ( .A(n9568), .B(n9567), .Z(n9569) );
  NAND U10335 ( .A(n9570), .B(n9569), .Z(n9589) );
  AND U10336 ( .A(b[2]), .B(a[358]), .Z(n9595) );
  AND U10337 ( .A(a[359]), .B(b[1]), .Z(n9593) );
  AND U10338 ( .A(a[357]), .B(b[3]), .Z(n9592) );
  XOR U10339 ( .A(n9593), .B(n9592), .Z(n9594) );
  XOR U10340 ( .A(n9595), .B(n9594), .Z(n9598) );
  NAND U10341 ( .A(b[0]), .B(a[360]), .Z(n9599) );
  XOR U10342 ( .A(n9598), .B(n9599), .Z(n9601) );
  OR U10343 ( .A(n9572), .B(n9571), .Z(n9576) );
  NANDN U10344 ( .A(n9574), .B(n9573), .Z(n9575) );
  NAND U10345 ( .A(n9576), .B(n9575), .Z(n9600) );
  XNOR U10346 ( .A(n9601), .B(n9600), .Z(n9586) );
  NANDN U10347 ( .A(n9578), .B(n9577), .Z(n9582) );
  OR U10348 ( .A(n9580), .B(n9579), .Z(n9581) );
  NAND U10349 ( .A(n9582), .B(n9581), .Z(n9587) );
  XNOR U10350 ( .A(n9586), .B(n9587), .Z(n9588) );
  XOR U10351 ( .A(n9589), .B(n9588), .Z(n9605) );
  XOR U10352 ( .A(sreg[1380]), .B(n9604), .Z(n9585) );
  XOR U10353 ( .A(n9605), .B(n9585), .Z(c[1380]) );
  NANDN U10354 ( .A(n9587), .B(n9586), .Z(n9591) );
  NAND U10355 ( .A(n9589), .B(n9588), .Z(n9590) );
  NAND U10356 ( .A(n9591), .B(n9590), .Z(n9610) );
  AND U10357 ( .A(b[2]), .B(a[359]), .Z(n9616) );
  AND U10358 ( .A(a[360]), .B(b[1]), .Z(n9614) );
  AND U10359 ( .A(a[358]), .B(b[3]), .Z(n9613) );
  XOR U10360 ( .A(n9614), .B(n9613), .Z(n9615) );
  XOR U10361 ( .A(n9616), .B(n9615), .Z(n9619) );
  NAND U10362 ( .A(b[0]), .B(a[361]), .Z(n9620) );
  XOR U10363 ( .A(n9619), .B(n9620), .Z(n9622) );
  OR U10364 ( .A(n9593), .B(n9592), .Z(n9597) );
  NANDN U10365 ( .A(n9595), .B(n9594), .Z(n9596) );
  NAND U10366 ( .A(n9597), .B(n9596), .Z(n9621) );
  XNOR U10367 ( .A(n9622), .B(n9621), .Z(n9607) );
  NANDN U10368 ( .A(n9599), .B(n9598), .Z(n9603) );
  OR U10369 ( .A(n9601), .B(n9600), .Z(n9602) );
  NAND U10370 ( .A(n9603), .B(n9602), .Z(n9608) );
  XNOR U10371 ( .A(n9607), .B(n9608), .Z(n9609) );
  XOR U10372 ( .A(n9610), .B(n9609), .Z(n9626) );
  XNOR U10373 ( .A(sreg[1381]), .B(n9625), .Z(n9606) );
  XOR U10374 ( .A(n9626), .B(n9606), .Z(c[1381]) );
  NANDN U10375 ( .A(n9608), .B(n9607), .Z(n9612) );
  NAND U10376 ( .A(n9610), .B(n9609), .Z(n9611) );
  NAND U10377 ( .A(n9612), .B(n9611), .Z(n9631) );
  AND U10378 ( .A(b[2]), .B(a[360]), .Z(n9637) );
  AND U10379 ( .A(a[361]), .B(b[1]), .Z(n9635) );
  AND U10380 ( .A(a[359]), .B(b[3]), .Z(n9634) );
  XOR U10381 ( .A(n9635), .B(n9634), .Z(n9636) );
  XOR U10382 ( .A(n9637), .B(n9636), .Z(n9640) );
  NAND U10383 ( .A(b[0]), .B(a[362]), .Z(n9641) );
  XOR U10384 ( .A(n9640), .B(n9641), .Z(n9643) );
  OR U10385 ( .A(n9614), .B(n9613), .Z(n9618) );
  NANDN U10386 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U10387 ( .A(n9618), .B(n9617), .Z(n9642) );
  XNOR U10388 ( .A(n9643), .B(n9642), .Z(n9628) );
  NANDN U10389 ( .A(n9620), .B(n9619), .Z(n9624) );
  OR U10390 ( .A(n9622), .B(n9621), .Z(n9623) );
  NAND U10391 ( .A(n9624), .B(n9623), .Z(n9629) );
  XNOR U10392 ( .A(n9628), .B(n9629), .Z(n9630) );
  XNOR U10393 ( .A(n9631), .B(n9630), .Z(n9647) );
  XOR U10394 ( .A(n9646), .B(sreg[1382]), .Z(n9627) );
  XOR U10395 ( .A(n9647), .B(n9627), .Z(c[1382]) );
  NANDN U10396 ( .A(n9629), .B(n9628), .Z(n9633) );
  NAND U10397 ( .A(n9631), .B(n9630), .Z(n9632) );
  NAND U10398 ( .A(n9633), .B(n9632), .Z(n9654) );
  AND U10399 ( .A(b[2]), .B(a[361]), .Z(n9660) );
  AND U10400 ( .A(a[362]), .B(b[1]), .Z(n9658) );
  AND U10401 ( .A(a[360]), .B(b[3]), .Z(n9657) );
  XOR U10402 ( .A(n9658), .B(n9657), .Z(n9659) );
  XOR U10403 ( .A(n9660), .B(n9659), .Z(n9663) );
  NAND U10404 ( .A(b[0]), .B(a[363]), .Z(n9664) );
  XOR U10405 ( .A(n9663), .B(n9664), .Z(n9666) );
  OR U10406 ( .A(n9635), .B(n9634), .Z(n9639) );
  NANDN U10407 ( .A(n9637), .B(n9636), .Z(n9638) );
  NAND U10408 ( .A(n9639), .B(n9638), .Z(n9665) );
  XNOR U10409 ( .A(n9666), .B(n9665), .Z(n9651) );
  NANDN U10410 ( .A(n9641), .B(n9640), .Z(n9645) );
  OR U10411 ( .A(n9643), .B(n9642), .Z(n9644) );
  NAND U10412 ( .A(n9645), .B(n9644), .Z(n9652) );
  XNOR U10413 ( .A(n9651), .B(n9652), .Z(n9653) );
  XOR U10414 ( .A(n9654), .B(n9653), .Z(n9650) );
  XOR U10415 ( .A(sreg[1383]), .B(n9649), .Z(n9648) );
  XOR U10416 ( .A(n9650), .B(n9648), .Z(c[1383]) );
  NANDN U10417 ( .A(n9652), .B(n9651), .Z(n9656) );
  NAND U10418 ( .A(n9654), .B(n9653), .Z(n9655) );
  NAND U10419 ( .A(n9656), .B(n9655), .Z(n9672) );
  AND U10420 ( .A(b[2]), .B(a[362]), .Z(n9678) );
  AND U10421 ( .A(a[363]), .B(b[1]), .Z(n9676) );
  AND U10422 ( .A(a[361]), .B(b[3]), .Z(n9675) );
  XOR U10423 ( .A(n9676), .B(n9675), .Z(n9677) );
  XOR U10424 ( .A(n9678), .B(n9677), .Z(n9681) );
  NAND U10425 ( .A(b[0]), .B(a[364]), .Z(n9682) );
  XOR U10426 ( .A(n9681), .B(n9682), .Z(n9684) );
  OR U10427 ( .A(n9658), .B(n9657), .Z(n9662) );
  NANDN U10428 ( .A(n9660), .B(n9659), .Z(n9661) );
  NAND U10429 ( .A(n9662), .B(n9661), .Z(n9683) );
  XNOR U10430 ( .A(n9684), .B(n9683), .Z(n9669) );
  NANDN U10431 ( .A(n9664), .B(n9663), .Z(n9668) );
  OR U10432 ( .A(n9666), .B(n9665), .Z(n9667) );
  NAND U10433 ( .A(n9668), .B(n9667), .Z(n9670) );
  XNOR U10434 ( .A(n9669), .B(n9670), .Z(n9671) );
  XNOR U10435 ( .A(n9672), .B(n9671), .Z(n9687) );
  XNOR U10436 ( .A(n9687), .B(sreg[1384]), .Z(n9688) );
  XOR U10437 ( .A(n9689), .B(n9688), .Z(c[1384]) );
  NANDN U10438 ( .A(n9670), .B(n9669), .Z(n9674) );
  NAND U10439 ( .A(n9672), .B(n9671), .Z(n9673) );
  NAND U10440 ( .A(n9674), .B(n9673), .Z(n9695) );
  AND U10441 ( .A(b[2]), .B(a[363]), .Z(n9701) );
  AND U10442 ( .A(a[364]), .B(b[1]), .Z(n9699) );
  AND U10443 ( .A(a[362]), .B(b[3]), .Z(n9698) );
  XOR U10444 ( .A(n9699), .B(n9698), .Z(n9700) );
  XOR U10445 ( .A(n9701), .B(n9700), .Z(n9704) );
  NAND U10446 ( .A(b[0]), .B(a[365]), .Z(n9705) );
  XOR U10447 ( .A(n9704), .B(n9705), .Z(n9707) );
  OR U10448 ( .A(n9676), .B(n9675), .Z(n9680) );
  NANDN U10449 ( .A(n9678), .B(n9677), .Z(n9679) );
  NAND U10450 ( .A(n9680), .B(n9679), .Z(n9706) );
  XNOR U10451 ( .A(n9707), .B(n9706), .Z(n9692) );
  NANDN U10452 ( .A(n9682), .B(n9681), .Z(n9686) );
  OR U10453 ( .A(n9684), .B(n9683), .Z(n9685) );
  NAND U10454 ( .A(n9686), .B(n9685), .Z(n9693) );
  XNOR U10455 ( .A(n9692), .B(n9693), .Z(n9694) );
  XNOR U10456 ( .A(n9695), .B(n9694), .Z(n9710) );
  XNOR U10457 ( .A(n9710), .B(sreg[1385]), .Z(n9712) );
  NAND U10458 ( .A(n9687), .B(sreg[1384]), .Z(n9691) );
  OR U10459 ( .A(n9689), .B(n9688), .Z(n9690) );
  AND U10460 ( .A(n9691), .B(n9690), .Z(n9711) );
  XOR U10461 ( .A(n9712), .B(n9711), .Z(c[1385]) );
  NANDN U10462 ( .A(n9693), .B(n9692), .Z(n9697) );
  NAND U10463 ( .A(n9695), .B(n9694), .Z(n9696) );
  NAND U10464 ( .A(n9697), .B(n9696), .Z(n9718) );
  AND U10465 ( .A(b[2]), .B(a[364]), .Z(n9724) );
  AND U10466 ( .A(a[365]), .B(b[1]), .Z(n9722) );
  AND U10467 ( .A(a[363]), .B(b[3]), .Z(n9721) );
  XOR U10468 ( .A(n9722), .B(n9721), .Z(n9723) );
  XOR U10469 ( .A(n9724), .B(n9723), .Z(n9727) );
  NAND U10470 ( .A(b[0]), .B(a[366]), .Z(n9728) );
  XOR U10471 ( .A(n9727), .B(n9728), .Z(n9730) );
  OR U10472 ( .A(n9699), .B(n9698), .Z(n9703) );
  NANDN U10473 ( .A(n9701), .B(n9700), .Z(n9702) );
  NAND U10474 ( .A(n9703), .B(n9702), .Z(n9729) );
  XNOR U10475 ( .A(n9730), .B(n9729), .Z(n9715) );
  NANDN U10476 ( .A(n9705), .B(n9704), .Z(n9709) );
  OR U10477 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U10478 ( .A(n9709), .B(n9708), .Z(n9716) );
  XNOR U10479 ( .A(n9715), .B(n9716), .Z(n9717) );
  XNOR U10480 ( .A(n9718), .B(n9717), .Z(n9733) );
  XOR U10481 ( .A(sreg[1386]), .B(n9733), .Z(n9734) );
  NAND U10482 ( .A(n9710), .B(sreg[1385]), .Z(n9714) );
  OR U10483 ( .A(n9712), .B(n9711), .Z(n9713) );
  NAND U10484 ( .A(n9714), .B(n9713), .Z(n9735) );
  XOR U10485 ( .A(n9734), .B(n9735), .Z(c[1386]) );
  NANDN U10486 ( .A(n9716), .B(n9715), .Z(n9720) );
  NAND U10487 ( .A(n9718), .B(n9717), .Z(n9719) );
  NAND U10488 ( .A(n9720), .B(n9719), .Z(n9744) );
  AND U10489 ( .A(b[2]), .B(a[365]), .Z(n9750) );
  AND U10490 ( .A(a[366]), .B(b[1]), .Z(n9748) );
  AND U10491 ( .A(a[364]), .B(b[3]), .Z(n9747) );
  XOR U10492 ( .A(n9748), .B(n9747), .Z(n9749) );
  XOR U10493 ( .A(n9750), .B(n9749), .Z(n9753) );
  NAND U10494 ( .A(b[0]), .B(a[367]), .Z(n9754) );
  XOR U10495 ( .A(n9753), .B(n9754), .Z(n9756) );
  OR U10496 ( .A(n9722), .B(n9721), .Z(n9726) );
  NANDN U10497 ( .A(n9724), .B(n9723), .Z(n9725) );
  NAND U10498 ( .A(n9726), .B(n9725), .Z(n9755) );
  XNOR U10499 ( .A(n9756), .B(n9755), .Z(n9741) );
  NANDN U10500 ( .A(n9728), .B(n9727), .Z(n9732) );
  OR U10501 ( .A(n9730), .B(n9729), .Z(n9731) );
  NAND U10502 ( .A(n9732), .B(n9731), .Z(n9742) );
  XNOR U10503 ( .A(n9741), .B(n9742), .Z(n9743) );
  XOR U10504 ( .A(n9744), .B(n9743), .Z(n9740) );
  OR U10505 ( .A(n9733), .B(sreg[1386]), .Z(n9737) );
  NANDN U10506 ( .A(n9735), .B(n9734), .Z(n9736) );
  AND U10507 ( .A(n9737), .B(n9736), .Z(n9739) );
  XNOR U10508 ( .A(sreg[1387]), .B(n9739), .Z(n9738) );
  XOR U10509 ( .A(n9740), .B(n9738), .Z(c[1387]) );
  NANDN U10510 ( .A(n9742), .B(n9741), .Z(n9746) );
  NAND U10511 ( .A(n9744), .B(n9743), .Z(n9745) );
  NAND U10512 ( .A(n9746), .B(n9745), .Z(n9763) );
  AND U10513 ( .A(b[2]), .B(a[366]), .Z(n9769) );
  AND U10514 ( .A(a[367]), .B(b[1]), .Z(n9767) );
  AND U10515 ( .A(a[365]), .B(b[3]), .Z(n9766) );
  XOR U10516 ( .A(n9767), .B(n9766), .Z(n9768) );
  XOR U10517 ( .A(n9769), .B(n9768), .Z(n9772) );
  NAND U10518 ( .A(b[0]), .B(a[368]), .Z(n9773) );
  XOR U10519 ( .A(n9772), .B(n9773), .Z(n9775) );
  OR U10520 ( .A(n9748), .B(n9747), .Z(n9752) );
  NANDN U10521 ( .A(n9750), .B(n9749), .Z(n9751) );
  NAND U10522 ( .A(n9752), .B(n9751), .Z(n9774) );
  XNOR U10523 ( .A(n9775), .B(n9774), .Z(n9760) );
  NANDN U10524 ( .A(n9754), .B(n9753), .Z(n9758) );
  OR U10525 ( .A(n9756), .B(n9755), .Z(n9757) );
  NAND U10526 ( .A(n9758), .B(n9757), .Z(n9761) );
  XNOR U10527 ( .A(n9760), .B(n9761), .Z(n9762) );
  XNOR U10528 ( .A(n9763), .B(n9762), .Z(n9779) );
  XNOR U10529 ( .A(sreg[1388]), .B(n9779), .Z(n9759) );
  XOR U10530 ( .A(n9778), .B(n9759), .Z(c[1388]) );
  NANDN U10531 ( .A(n9761), .B(n9760), .Z(n9765) );
  NAND U10532 ( .A(n9763), .B(n9762), .Z(n9764) );
  NAND U10533 ( .A(n9765), .B(n9764), .Z(n9786) );
  AND U10534 ( .A(b[2]), .B(a[367]), .Z(n9792) );
  AND U10535 ( .A(a[368]), .B(b[1]), .Z(n9790) );
  AND U10536 ( .A(a[366]), .B(b[3]), .Z(n9789) );
  XOR U10537 ( .A(n9790), .B(n9789), .Z(n9791) );
  XOR U10538 ( .A(n9792), .B(n9791), .Z(n9795) );
  NAND U10539 ( .A(b[0]), .B(a[369]), .Z(n9796) );
  XOR U10540 ( .A(n9795), .B(n9796), .Z(n9798) );
  OR U10541 ( .A(n9767), .B(n9766), .Z(n9771) );
  NANDN U10542 ( .A(n9769), .B(n9768), .Z(n9770) );
  NAND U10543 ( .A(n9771), .B(n9770), .Z(n9797) );
  XNOR U10544 ( .A(n9798), .B(n9797), .Z(n9783) );
  NANDN U10545 ( .A(n9773), .B(n9772), .Z(n9777) );
  OR U10546 ( .A(n9775), .B(n9774), .Z(n9776) );
  NAND U10547 ( .A(n9777), .B(n9776), .Z(n9784) );
  XNOR U10548 ( .A(n9783), .B(n9784), .Z(n9785) );
  XOR U10549 ( .A(n9786), .B(n9785), .Z(n9782) );
  XNOR U10550 ( .A(sreg[1389]), .B(n9781), .Z(n9780) );
  XOR U10551 ( .A(n9782), .B(n9780), .Z(c[1389]) );
  NANDN U10552 ( .A(n9784), .B(n9783), .Z(n9788) );
  NAND U10553 ( .A(n9786), .B(n9785), .Z(n9787) );
  NAND U10554 ( .A(n9788), .B(n9787), .Z(n9804) );
  AND U10555 ( .A(b[2]), .B(a[368]), .Z(n9810) );
  AND U10556 ( .A(a[369]), .B(b[1]), .Z(n9808) );
  AND U10557 ( .A(a[367]), .B(b[3]), .Z(n9807) );
  XOR U10558 ( .A(n9808), .B(n9807), .Z(n9809) );
  XOR U10559 ( .A(n9810), .B(n9809), .Z(n9813) );
  NAND U10560 ( .A(b[0]), .B(a[370]), .Z(n9814) );
  XOR U10561 ( .A(n9813), .B(n9814), .Z(n9816) );
  OR U10562 ( .A(n9790), .B(n9789), .Z(n9794) );
  NANDN U10563 ( .A(n9792), .B(n9791), .Z(n9793) );
  NAND U10564 ( .A(n9794), .B(n9793), .Z(n9815) );
  XNOR U10565 ( .A(n9816), .B(n9815), .Z(n9801) );
  NANDN U10566 ( .A(n9796), .B(n9795), .Z(n9800) );
  OR U10567 ( .A(n9798), .B(n9797), .Z(n9799) );
  NAND U10568 ( .A(n9800), .B(n9799), .Z(n9802) );
  XNOR U10569 ( .A(n9801), .B(n9802), .Z(n9803) );
  XNOR U10570 ( .A(n9804), .B(n9803), .Z(n9819) );
  XNOR U10571 ( .A(n9819), .B(sreg[1390]), .Z(n9820) );
  XOR U10572 ( .A(n9821), .B(n9820), .Z(c[1390]) );
  NANDN U10573 ( .A(n9802), .B(n9801), .Z(n9806) );
  NAND U10574 ( .A(n9804), .B(n9803), .Z(n9805) );
  NAND U10575 ( .A(n9806), .B(n9805), .Z(n9827) );
  AND U10576 ( .A(b[2]), .B(a[369]), .Z(n9833) );
  AND U10577 ( .A(a[370]), .B(b[1]), .Z(n9831) );
  AND U10578 ( .A(a[368]), .B(b[3]), .Z(n9830) );
  XOR U10579 ( .A(n9831), .B(n9830), .Z(n9832) );
  XOR U10580 ( .A(n9833), .B(n9832), .Z(n9836) );
  NAND U10581 ( .A(b[0]), .B(a[371]), .Z(n9837) );
  XOR U10582 ( .A(n9836), .B(n9837), .Z(n9839) );
  OR U10583 ( .A(n9808), .B(n9807), .Z(n9812) );
  NANDN U10584 ( .A(n9810), .B(n9809), .Z(n9811) );
  NAND U10585 ( .A(n9812), .B(n9811), .Z(n9838) );
  XNOR U10586 ( .A(n9839), .B(n9838), .Z(n9824) );
  NANDN U10587 ( .A(n9814), .B(n9813), .Z(n9818) );
  OR U10588 ( .A(n9816), .B(n9815), .Z(n9817) );
  NAND U10589 ( .A(n9818), .B(n9817), .Z(n9825) );
  XNOR U10590 ( .A(n9824), .B(n9825), .Z(n9826) );
  XNOR U10591 ( .A(n9827), .B(n9826), .Z(n9842) );
  XNOR U10592 ( .A(n9842), .B(sreg[1391]), .Z(n9844) );
  NAND U10593 ( .A(n9819), .B(sreg[1390]), .Z(n9823) );
  OR U10594 ( .A(n9821), .B(n9820), .Z(n9822) );
  AND U10595 ( .A(n9823), .B(n9822), .Z(n9843) );
  XOR U10596 ( .A(n9844), .B(n9843), .Z(c[1391]) );
  NANDN U10597 ( .A(n9825), .B(n9824), .Z(n9829) );
  NAND U10598 ( .A(n9827), .B(n9826), .Z(n9828) );
  NAND U10599 ( .A(n9829), .B(n9828), .Z(n9853) );
  AND U10600 ( .A(b[2]), .B(a[370]), .Z(n9865) );
  AND U10601 ( .A(a[371]), .B(b[1]), .Z(n9863) );
  AND U10602 ( .A(a[369]), .B(b[3]), .Z(n9862) );
  XOR U10603 ( .A(n9863), .B(n9862), .Z(n9864) );
  XOR U10604 ( .A(n9865), .B(n9864), .Z(n9856) );
  NAND U10605 ( .A(b[0]), .B(a[372]), .Z(n9857) );
  XOR U10606 ( .A(n9856), .B(n9857), .Z(n9859) );
  OR U10607 ( .A(n9831), .B(n9830), .Z(n9835) );
  NANDN U10608 ( .A(n9833), .B(n9832), .Z(n9834) );
  NAND U10609 ( .A(n9835), .B(n9834), .Z(n9858) );
  XNOR U10610 ( .A(n9859), .B(n9858), .Z(n9850) );
  NANDN U10611 ( .A(n9837), .B(n9836), .Z(n9841) );
  OR U10612 ( .A(n9839), .B(n9838), .Z(n9840) );
  NAND U10613 ( .A(n9841), .B(n9840), .Z(n9851) );
  XNOR U10614 ( .A(n9850), .B(n9851), .Z(n9852) );
  XOR U10615 ( .A(n9853), .B(n9852), .Z(n9849) );
  NAND U10616 ( .A(n9842), .B(sreg[1391]), .Z(n9846) );
  OR U10617 ( .A(n9844), .B(n9843), .Z(n9845) );
  NAND U10618 ( .A(n9846), .B(n9845), .Z(n9848) );
  XNOR U10619 ( .A(sreg[1392]), .B(n9848), .Z(n9847) );
  XOR U10620 ( .A(n9849), .B(n9847), .Z(c[1392]) );
  NANDN U10621 ( .A(n9851), .B(n9850), .Z(n9855) );
  NAND U10622 ( .A(n9853), .B(n9852), .Z(n9854) );
  AND U10623 ( .A(n9855), .B(n9854), .Z(n9871) );
  NANDN U10624 ( .A(n9857), .B(n9856), .Z(n9861) );
  OR U10625 ( .A(n9859), .B(n9858), .Z(n9860) );
  AND U10626 ( .A(n9861), .B(n9860), .Z(n9870) );
  AND U10627 ( .A(b[2]), .B(a[371]), .Z(n9875) );
  AND U10628 ( .A(a[372]), .B(b[1]), .Z(n9873) );
  AND U10629 ( .A(a[370]), .B(b[3]), .Z(n9872) );
  XOR U10630 ( .A(n9873), .B(n9872), .Z(n9874) );
  XOR U10631 ( .A(n9875), .B(n9874), .Z(n9878) );
  NAND U10632 ( .A(b[0]), .B(a[373]), .Z(n9879) );
  XOR U10633 ( .A(n9878), .B(n9879), .Z(n9881) );
  OR U10634 ( .A(n9863), .B(n9862), .Z(n9867) );
  NANDN U10635 ( .A(n9865), .B(n9864), .Z(n9866) );
  NAND U10636 ( .A(n9867), .B(n9866), .Z(n9880) );
  XOR U10637 ( .A(n9881), .B(n9880), .Z(n9869) );
  XNOR U10638 ( .A(n9870), .B(n9869), .Z(n9868) );
  XOR U10639 ( .A(n9871), .B(n9868), .Z(n9884) );
  XNOR U10640 ( .A(sreg[1393]), .B(n9884), .Z(n9885) );
  XOR U10641 ( .A(n9886), .B(n9885), .Z(c[1393]) );
  AND U10642 ( .A(b[2]), .B(a[372]), .Z(n9901) );
  AND U10643 ( .A(a[373]), .B(b[1]), .Z(n9899) );
  AND U10644 ( .A(a[371]), .B(b[3]), .Z(n9898) );
  XOR U10645 ( .A(n9899), .B(n9898), .Z(n9900) );
  XOR U10646 ( .A(n9901), .B(n9900), .Z(n9904) );
  NAND U10647 ( .A(b[0]), .B(a[374]), .Z(n9905) );
  XOR U10648 ( .A(n9904), .B(n9905), .Z(n9907) );
  OR U10649 ( .A(n9873), .B(n9872), .Z(n9877) );
  NANDN U10650 ( .A(n9875), .B(n9874), .Z(n9876) );
  NAND U10651 ( .A(n9877), .B(n9876), .Z(n9906) );
  XNOR U10652 ( .A(n9907), .B(n9906), .Z(n9892) );
  NANDN U10653 ( .A(n9879), .B(n9878), .Z(n9883) );
  OR U10654 ( .A(n9881), .B(n9880), .Z(n9882) );
  NAND U10655 ( .A(n9883), .B(n9882), .Z(n9893) );
  XNOR U10656 ( .A(n9892), .B(n9893), .Z(n9894) );
  XNOR U10657 ( .A(n9895), .B(n9894), .Z(n9891) );
  NAND U10658 ( .A(sreg[1393]), .B(n9884), .Z(n9888) );
  OR U10659 ( .A(n9886), .B(n9885), .Z(n9887) );
  AND U10660 ( .A(n9888), .B(n9887), .Z(n9890) );
  XNOR U10661 ( .A(n9890), .B(sreg[1394]), .Z(n9889) );
  XNOR U10662 ( .A(n9891), .B(n9889), .Z(c[1394]) );
  NANDN U10663 ( .A(n9893), .B(n9892), .Z(n9897) );
  NANDN U10664 ( .A(n9895), .B(n9894), .Z(n9896) );
  NAND U10665 ( .A(n9897), .B(n9896), .Z(n9913) );
  AND U10666 ( .A(b[2]), .B(a[373]), .Z(n9919) );
  AND U10667 ( .A(a[374]), .B(b[1]), .Z(n9917) );
  AND U10668 ( .A(a[372]), .B(b[3]), .Z(n9916) );
  XOR U10669 ( .A(n9917), .B(n9916), .Z(n9918) );
  XOR U10670 ( .A(n9919), .B(n9918), .Z(n9922) );
  NAND U10671 ( .A(b[0]), .B(a[375]), .Z(n9923) );
  XOR U10672 ( .A(n9922), .B(n9923), .Z(n9925) );
  OR U10673 ( .A(n9899), .B(n9898), .Z(n9903) );
  NANDN U10674 ( .A(n9901), .B(n9900), .Z(n9902) );
  NAND U10675 ( .A(n9903), .B(n9902), .Z(n9924) );
  XNOR U10676 ( .A(n9925), .B(n9924), .Z(n9910) );
  NANDN U10677 ( .A(n9905), .B(n9904), .Z(n9909) );
  OR U10678 ( .A(n9907), .B(n9906), .Z(n9908) );
  NAND U10679 ( .A(n9909), .B(n9908), .Z(n9911) );
  XNOR U10680 ( .A(n9910), .B(n9911), .Z(n9912) );
  XNOR U10681 ( .A(n9913), .B(n9912), .Z(n9929) );
  XNOR U10682 ( .A(n9929), .B(sreg[1395]), .Z(n9931) );
  XNOR U10683 ( .A(n9930), .B(n9931), .Z(c[1395]) );
  NANDN U10684 ( .A(n9911), .B(n9910), .Z(n9915) );
  NAND U10685 ( .A(n9913), .B(n9912), .Z(n9914) );
  AND U10686 ( .A(n9915), .B(n9914), .Z(n9936) );
  AND U10687 ( .A(b[2]), .B(a[374]), .Z(n9940) );
  AND U10688 ( .A(a[375]), .B(b[1]), .Z(n9938) );
  AND U10689 ( .A(a[373]), .B(b[3]), .Z(n9937) );
  XOR U10690 ( .A(n9938), .B(n9937), .Z(n9939) );
  XOR U10691 ( .A(n9940), .B(n9939), .Z(n9943) );
  NAND U10692 ( .A(b[0]), .B(a[376]), .Z(n9944) );
  XOR U10693 ( .A(n9943), .B(n9944), .Z(n9945) );
  OR U10694 ( .A(n9917), .B(n9916), .Z(n9921) );
  NANDN U10695 ( .A(n9919), .B(n9918), .Z(n9920) );
  AND U10696 ( .A(n9921), .B(n9920), .Z(n9946) );
  XOR U10697 ( .A(n9945), .B(n9946), .Z(n9934) );
  NANDN U10698 ( .A(n9923), .B(n9922), .Z(n9927) );
  OR U10699 ( .A(n9925), .B(n9924), .Z(n9926) );
  AND U10700 ( .A(n9927), .B(n9926), .Z(n9935) );
  XOR U10701 ( .A(n9934), .B(n9935), .Z(n9928) );
  XOR U10702 ( .A(n9936), .B(n9928), .Z(n9947) );
  XNOR U10703 ( .A(sreg[1396]), .B(n9947), .Z(n9949) );
  NAND U10704 ( .A(n9929), .B(sreg[1395]), .Z(n9933) );
  NANDN U10705 ( .A(n9931), .B(n9930), .Z(n9932) );
  AND U10706 ( .A(n9933), .B(n9932), .Z(n9948) );
  XOR U10707 ( .A(n9949), .B(n9948), .Z(c[1396]) );
  AND U10708 ( .A(b[2]), .B(a[375]), .Z(n9964) );
  AND U10709 ( .A(a[376]), .B(b[1]), .Z(n9962) );
  AND U10710 ( .A(a[374]), .B(b[3]), .Z(n9961) );
  XOR U10711 ( .A(n9962), .B(n9961), .Z(n9963) );
  XOR U10712 ( .A(n9964), .B(n9963), .Z(n9967) );
  NAND U10713 ( .A(b[0]), .B(a[377]), .Z(n9968) );
  XOR U10714 ( .A(n9967), .B(n9968), .Z(n9970) );
  OR U10715 ( .A(n9938), .B(n9937), .Z(n9942) );
  NANDN U10716 ( .A(n9940), .B(n9939), .Z(n9941) );
  NAND U10717 ( .A(n9942), .B(n9941), .Z(n9969) );
  XNOR U10718 ( .A(n9970), .B(n9969), .Z(n9955) );
  XNOR U10719 ( .A(n9955), .B(n9956), .Z(n9958) );
  XOR U10720 ( .A(n9957), .B(n9958), .Z(n9954) );
  NAND U10721 ( .A(sreg[1396]), .B(n9947), .Z(n9951) );
  OR U10722 ( .A(n9949), .B(n9948), .Z(n9950) );
  AND U10723 ( .A(n9951), .B(n9950), .Z(n9953) );
  XNOR U10724 ( .A(n9953), .B(sreg[1397]), .Z(n9952) );
  XNOR U10725 ( .A(n9954), .B(n9952), .Z(c[1397]) );
  NANDN U10726 ( .A(n9956), .B(n9955), .Z(n9960) );
  NAND U10727 ( .A(n9958), .B(n9957), .Z(n9959) );
  NAND U10728 ( .A(n9960), .B(n9959), .Z(n9976) );
  AND U10729 ( .A(b[2]), .B(a[376]), .Z(n9988) );
  AND U10730 ( .A(a[377]), .B(b[1]), .Z(n9986) );
  AND U10731 ( .A(a[375]), .B(b[3]), .Z(n9985) );
  XOR U10732 ( .A(n9986), .B(n9985), .Z(n9987) );
  XOR U10733 ( .A(n9988), .B(n9987), .Z(n9979) );
  NAND U10734 ( .A(b[0]), .B(a[378]), .Z(n9980) );
  XOR U10735 ( .A(n9979), .B(n9980), .Z(n9982) );
  OR U10736 ( .A(n9962), .B(n9961), .Z(n9966) );
  NANDN U10737 ( .A(n9964), .B(n9963), .Z(n9965) );
  NAND U10738 ( .A(n9966), .B(n9965), .Z(n9981) );
  XNOR U10739 ( .A(n9982), .B(n9981), .Z(n9973) );
  NANDN U10740 ( .A(n9968), .B(n9967), .Z(n9972) );
  OR U10741 ( .A(n9970), .B(n9969), .Z(n9971) );
  NAND U10742 ( .A(n9972), .B(n9971), .Z(n9974) );
  XNOR U10743 ( .A(n9973), .B(n9974), .Z(n9975) );
  XNOR U10744 ( .A(n9976), .B(n9975), .Z(n9992) );
  XNOR U10745 ( .A(n9992), .B(sreg[1398]), .Z(n9994) );
  XNOR U10746 ( .A(n9993), .B(n9994), .Z(c[1398]) );
  NANDN U10747 ( .A(n9974), .B(n9973), .Z(n9978) );
  NAND U10748 ( .A(n9976), .B(n9975), .Z(n9977) );
  AND U10749 ( .A(n9978), .B(n9977), .Z(n9999) );
  NANDN U10750 ( .A(n9980), .B(n9979), .Z(n9984) );
  OR U10751 ( .A(n9982), .B(n9981), .Z(n9983) );
  AND U10752 ( .A(n9984), .B(n9983), .Z(n9998) );
  AND U10753 ( .A(b[2]), .B(a[377]), .Z(n10003) );
  AND U10754 ( .A(a[378]), .B(b[1]), .Z(n10001) );
  AND U10755 ( .A(a[376]), .B(b[3]), .Z(n10000) );
  XOR U10756 ( .A(n10001), .B(n10000), .Z(n10002) );
  XOR U10757 ( .A(n10003), .B(n10002), .Z(n10006) );
  NAND U10758 ( .A(b[0]), .B(a[379]), .Z(n10007) );
  XOR U10759 ( .A(n10006), .B(n10007), .Z(n10009) );
  OR U10760 ( .A(n9986), .B(n9985), .Z(n9990) );
  NANDN U10761 ( .A(n9988), .B(n9987), .Z(n9989) );
  NAND U10762 ( .A(n9990), .B(n9989), .Z(n10008) );
  XOR U10763 ( .A(n10009), .B(n10008), .Z(n9997) );
  XNOR U10764 ( .A(n9998), .B(n9997), .Z(n9991) );
  XOR U10765 ( .A(n9999), .B(n9991), .Z(n10012) );
  XNOR U10766 ( .A(sreg[1399]), .B(n10012), .Z(n10014) );
  NAND U10767 ( .A(n9992), .B(sreg[1398]), .Z(n9996) );
  NANDN U10768 ( .A(n9994), .B(n9993), .Z(n9995) );
  AND U10769 ( .A(n9996), .B(n9995), .Z(n10013) );
  XOR U10770 ( .A(n10014), .B(n10013), .Z(c[1399]) );
  AND U10771 ( .A(b[2]), .B(a[378]), .Z(n10026) );
  AND U10772 ( .A(a[379]), .B(b[1]), .Z(n10024) );
  AND U10773 ( .A(a[377]), .B(b[3]), .Z(n10023) );
  XOR U10774 ( .A(n10024), .B(n10023), .Z(n10025) );
  XOR U10775 ( .A(n10026), .B(n10025), .Z(n10029) );
  NAND U10776 ( .A(b[0]), .B(a[380]), .Z(n10030) );
  XOR U10777 ( .A(n10029), .B(n10030), .Z(n10032) );
  OR U10778 ( .A(n10001), .B(n10000), .Z(n10005) );
  NANDN U10779 ( .A(n10003), .B(n10002), .Z(n10004) );
  NAND U10780 ( .A(n10005), .B(n10004), .Z(n10031) );
  XNOR U10781 ( .A(n10032), .B(n10031), .Z(n10017) );
  NANDN U10782 ( .A(n10007), .B(n10006), .Z(n10011) );
  OR U10783 ( .A(n10009), .B(n10008), .Z(n10010) );
  NAND U10784 ( .A(n10011), .B(n10010), .Z(n10018) );
  XNOR U10785 ( .A(n10017), .B(n10018), .Z(n10019) );
  XOR U10786 ( .A(n10020), .B(n10019), .Z(n10035) );
  XNOR U10787 ( .A(n10035), .B(sreg[1400]), .Z(n10037) );
  NAND U10788 ( .A(sreg[1399]), .B(n10012), .Z(n10016) );
  OR U10789 ( .A(n10014), .B(n10013), .Z(n10015) );
  AND U10790 ( .A(n10016), .B(n10015), .Z(n10036) );
  XOR U10791 ( .A(n10037), .B(n10036), .Z(c[1400]) );
  NANDN U10792 ( .A(n10018), .B(n10017), .Z(n10022) );
  NANDN U10793 ( .A(n10020), .B(n10019), .Z(n10021) );
  NAND U10794 ( .A(n10022), .B(n10021), .Z(n10046) );
  AND U10795 ( .A(b[2]), .B(a[379]), .Z(n10052) );
  AND U10796 ( .A(a[380]), .B(b[1]), .Z(n10050) );
  AND U10797 ( .A(a[378]), .B(b[3]), .Z(n10049) );
  XOR U10798 ( .A(n10050), .B(n10049), .Z(n10051) );
  XOR U10799 ( .A(n10052), .B(n10051), .Z(n10055) );
  NAND U10800 ( .A(b[0]), .B(a[381]), .Z(n10056) );
  XOR U10801 ( .A(n10055), .B(n10056), .Z(n10058) );
  OR U10802 ( .A(n10024), .B(n10023), .Z(n10028) );
  NANDN U10803 ( .A(n10026), .B(n10025), .Z(n10027) );
  NAND U10804 ( .A(n10028), .B(n10027), .Z(n10057) );
  XNOR U10805 ( .A(n10058), .B(n10057), .Z(n10043) );
  NANDN U10806 ( .A(n10030), .B(n10029), .Z(n10034) );
  OR U10807 ( .A(n10032), .B(n10031), .Z(n10033) );
  NAND U10808 ( .A(n10034), .B(n10033), .Z(n10044) );
  XNOR U10809 ( .A(n10043), .B(n10044), .Z(n10045) );
  XOR U10810 ( .A(n10046), .B(n10045), .Z(n10042) );
  NAND U10811 ( .A(n10035), .B(sreg[1400]), .Z(n10039) );
  OR U10812 ( .A(n10037), .B(n10036), .Z(n10038) );
  NAND U10813 ( .A(n10039), .B(n10038), .Z(n10041) );
  XNOR U10814 ( .A(sreg[1401]), .B(n10041), .Z(n10040) );
  XOR U10815 ( .A(n10042), .B(n10040), .Z(c[1401]) );
  NANDN U10816 ( .A(n10044), .B(n10043), .Z(n10048) );
  NAND U10817 ( .A(n10046), .B(n10045), .Z(n10047) );
  AND U10818 ( .A(n10048), .B(n10047), .Z(n10065) );
  AND U10819 ( .A(b[2]), .B(a[380]), .Z(n10069) );
  AND U10820 ( .A(a[381]), .B(b[1]), .Z(n10067) );
  AND U10821 ( .A(a[379]), .B(b[3]), .Z(n10066) );
  XOR U10822 ( .A(n10067), .B(n10066), .Z(n10068) );
  XOR U10823 ( .A(n10069), .B(n10068), .Z(n10072) );
  NAND U10824 ( .A(b[0]), .B(a[382]), .Z(n10073) );
  XOR U10825 ( .A(n10072), .B(n10073), .Z(n10074) );
  OR U10826 ( .A(n10050), .B(n10049), .Z(n10054) );
  NANDN U10827 ( .A(n10052), .B(n10051), .Z(n10053) );
  AND U10828 ( .A(n10054), .B(n10053), .Z(n10075) );
  XOR U10829 ( .A(n10074), .B(n10075), .Z(n10063) );
  NANDN U10830 ( .A(n10056), .B(n10055), .Z(n10060) );
  OR U10831 ( .A(n10058), .B(n10057), .Z(n10059) );
  AND U10832 ( .A(n10060), .B(n10059), .Z(n10064) );
  XOR U10833 ( .A(n10063), .B(n10064), .Z(n10061) );
  XOR U10834 ( .A(n10065), .B(n10061), .Z(n10076) );
  XNOR U10835 ( .A(sreg[1402]), .B(n10076), .Z(n10062) );
  XOR U10836 ( .A(n10077), .B(n10062), .Z(c[1402]) );
  AND U10837 ( .A(b[2]), .B(a[381]), .Z(n10090) );
  AND U10838 ( .A(a[382]), .B(b[1]), .Z(n10088) );
  AND U10839 ( .A(a[380]), .B(b[3]), .Z(n10087) );
  XOR U10840 ( .A(n10088), .B(n10087), .Z(n10089) );
  XOR U10841 ( .A(n10090), .B(n10089), .Z(n10093) );
  NAND U10842 ( .A(b[0]), .B(a[383]), .Z(n10094) );
  XOR U10843 ( .A(n10093), .B(n10094), .Z(n10096) );
  OR U10844 ( .A(n10067), .B(n10066), .Z(n10071) );
  NANDN U10845 ( .A(n10069), .B(n10068), .Z(n10070) );
  NAND U10846 ( .A(n10071), .B(n10070), .Z(n10095) );
  XNOR U10847 ( .A(n10096), .B(n10095), .Z(n10081) );
  XNOR U10848 ( .A(n10081), .B(n10082), .Z(n10084) );
  XOR U10849 ( .A(n10083), .B(n10084), .Z(n10080) );
  XNOR U10850 ( .A(sreg[1403]), .B(n10079), .Z(n10078) );
  XOR U10851 ( .A(n10080), .B(n10078), .Z(c[1403]) );
  NANDN U10852 ( .A(n10082), .B(n10081), .Z(n10086) );
  NAND U10853 ( .A(n10084), .B(n10083), .Z(n10085) );
  NAND U10854 ( .A(n10086), .B(n10085), .Z(n10102) );
  AND U10855 ( .A(b[2]), .B(a[382]), .Z(n10114) );
  AND U10856 ( .A(a[383]), .B(b[1]), .Z(n10112) );
  AND U10857 ( .A(a[381]), .B(b[3]), .Z(n10111) );
  XOR U10858 ( .A(n10112), .B(n10111), .Z(n10113) );
  XOR U10859 ( .A(n10114), .B(n10113), .Z(n10105) );
  NAND U10860 ( .A(b[0]), .B(a[384]), .Z(n10106) );
  XOR U10861 ( .A(n10105), .B(n10106), .Z(n10108) );
  OR U10862 ( .A(n10088), .B(n10087), .Z(n10092) );
  NANDN U10863 ( .A(n10090), .B(n10089), .Z(n10091) );
  NAND U10864 ( .A(n10092), .B(n10091), .Z(n10107) );
  XNOR U10865 ( .A(n10108), .B(n10107), .Z(n10099) );
  NANDN U10866 ( .A(n10094), .B(n10093), .Z(n10098) );
  OR U10867 ( .A(n10096), .B(n10095), .Z(n10097) );
  NAND U10868 ( .A(n10098), .B(n10097), .Z(n10100) );
  XNOR U10869 ( .A(n10099), .B(n10100), .Z(n10101) );
  XNOR U10870 ( .A(n10102), .B(n10101), .Z(n10118) );
  XNOR U10871 ( .A(n10118), .B(sreg[1404]), .Z(n10119) );
  XOR U10872 ( .A(n10120), .B(n10119), .Z(c[1404]) );
  NANDN U10873 ( .A(n10100), .B(n10099), .Z(n10104) );
  NAND U10874 ( .A(n10102), .B(n10101), .Z(n10103) );
  NAND U10875 ( .A(n10104), .B(n10103), .Z(n10125) );
  NANDN U10876 ( .A(n10106), .B(n10105), .Z(n10110) );
  OR U10877 ( .A(n10108), .B(n10107), .Z(n10109) );
  AND U10878 ( .A(n10110), .B(n10109), .Z(n10124) );
  AND U10879 ( .A(b[2]), .B(a[383]), .Z(n10129) );
  AND U10880 ( .A(a[384]), .B(b[1]), .Z(n10127) );
  AND U10881 ( .A(a[382]), .B(b[3]), .Z(n10126) );
  XOR U10882 ( .A(n10127), .B(n10126), .Z(n10128) );
  XOR U10883 ( .A(n10129), .B(n10128), .Z(n10132) );
  NAND U10884 ( .A(b[0]), .B(a[385]), .Z(n10133) );
  XOR U10885 ( .A(n10132), .B(n10133), .Z(n10135) );
  OR U10886 ( .A(n10112), .B(n10111), .Z(n10116) );
  NANDN U10887 ( .A(n10114), .B(n10113), .Z(n10115) );
  NAND U10888 ( .A(n10116), .B(n10115), .Z(n10134) );
  XOR U10889 ( .A(n10135), .B(n10134), .Z(n10123) );
  XNOR U10890 ( .A(n10124), .B(n10123), .Z(n10117) );
  XNOR U10891 ( .A(n10125), .B(n10117), .Z(n10138) );
  XOR U10892 ( .A(sreg[1405]), .B(n10138), .Z(n10139) );
  NAND U10893 ( .A(n10118), .B(sreg[1404]), .Z(n10122) );
  OR U10894 ( .A(n10120), .B(n10119), .Z(n10121) );
  NAND U10895 ( .A(n10122), .B(n10121), .Z(n10140) );
  XOR U10896 ( .A(n10139), .B(n10140), .Z(c[1405]) );
  AND U10897 ( .A(b[2]), .B(a[384]), .Z(n10152) );
  AND U10898 ( .A(a[385]), .B(b[1]), .Z(n10150) );
  AND U10899 ( .A(a[383]), .B(b[3]), .Z(n10149) );
  XOR U10900 ( .A(n10150), .B(n10149), .Z(n10151) );
  XOR U10901 ( .A(n10152), .B(n10151), .Z(n10155) );
  NAND U10902 ( .A(b[0]), .B(a[386]), .Z(n10156) );
  XOR U10903 ( .A(n10155), .B(n10156), .Z(n10158) );
  OR U10904 ( .A(n10127), .B(n10126), .Z(n10131) );
  NANDN U10905 ( .A(n10129), .B(n10128), .Z(n10130) );
  NAND U10906 ( .A(n10131), .B(n10130), .Z(n10157) );
  XNOR U10907 ( .A(n10158), .B(n10157), .Z(n10143) );
  NANDN U10908 ( .A(n10133), .B(n10132), .Z(n10137) );
  OR U10909 ( .A(n10135), .B(n10134), .Z(n10136) );
  NAND U10910 ( .A(n10137), .B(n10136), .Z(n10144) );
  XNOR U10911 ( .A(n10143), .B(n10144), .Z(n10145) );
  XNOR U10912 ( .A(n10146), .B(n10145), .Z(n10161) );
  XOR U10913 ( .A(sreg[1406]), .B(n10161), .Z(n10163) );
  OR U10914 ( .A(n10138), .B(sreg[1405]), .Z(n10142) );
  NANDN U10915 ( .A(n10140), .B(n10139), .Z(n10141) );
  AND U10916 ( .A(n10142), .B(n10141), .Z(n10162) );
  XNOR U10917 ( .A(n10163), .B(n10162), .Z(c[1406]) );
  NANDN U10918 ( .A(n10144), .B(n10143), .Z(n10148) );
  NANDN U10919 ( .A(n10146), .B(n10145), .Z(n10147) );
  NAND U10920 ( .A(n10148), .B(n10147), .Z(n10172) );
  AND U10921 ( .A(b[2]), .B(a[385]), .Z(n10178) );
  AND U10922 ( .A(a[386]), .B(b[1]), .Z(n10176) );
  AND U10923 ( .A(a[384]), .B(b[3]), .Z(n10175) );
  XOR U10924 ( .A(n10176), .B(n10175), .Z(n10177) );
  XOR U10925 ( .A(n10178), .B(n10177), .Z(n10181) );
  NAND U10926 ( .A(b[0]), .B(a[387]), .Z(n10182) );
  XOR U10927 ( .A(n10181), .B(n10182), .Z(n10184) );
  OR U10928 ( .A(n10150), .B(n10149), .Z(n10154) );
  NANDN U10929 ( .A(n10152), .B(n10151), .Z(n10153) );
  NAND U10930 ( .A(n10154), .B(n10153), .Z(n10183) );
  XNOR U10931 ( .A(n10184), .B(n10183), .Z(n10169) );
  NANDN U10932 ( .A(n10156), .B(n10155), .Z(n10160) );
  OR U10933 ( .A(n10158), .B(n10157), .Z(n10159) );
  NAND U10934 ( .A(n10160), .B(n10159), .Z(n10170) );
  XNOR U10935 ( .A(n10169), .B(n10170), .Z(n10171) );
  XOR U10936 ( .A(n10172), .B(n10171), .Z(n10168) );
  NANDN U10937 ( .A(sreg[1406]), .B(n10161), .Z(n10165) );
  OR U10938 ( .A(n10163), .B(n10162), .Z(n10164) );
  AND U10939 ( .A(n10165), .B(n10164), .Z(n10167) );
  XNOR U10940 ( .A(sreg[1407]), .B(n10167), .Z(n10166) );
  XOR U10941 ( .A(n10168), .B(n10166), .Z(c[1407]) );
  NANDN U10942 ( .A(n10170), .B(n10169), .Z(n10174) );
  NAND U10943 ( .A(n10172), .B(n10171), .Z(n10173) );
  AND U10944 ( .A(n10174), .B(n10173), .Z(n10190) );
  AND U10945 ( .A(b[2]), .B(a[386]), .Z(n10194) );
  AND U10946 ( .A(a[387]), .B(b[1]), .Z(n10192) );
  AND U10947 ( .A(a[385]), .B(b[3]), .Z(n10191) );
  XOR U10948 ( .A(n10192), .B(n10191), .Z(n10193) );
  XOR U10949 ( .A(n10194), .B(n10193), .Z(n10197) );
  NAND U10950 ( .A(b[0]), .B(a[388]), .Z(n10198) );
  XOR U10951 ( .A(n10197), .B(n10198), .Z(n10199) );
  OR U10952 ( .A(n10176), .B(n10175), .Z(n10180) );
  NANDN U10953 ( .A(n10178), .B(n10177), .Z(n10179) );
  AND U10954 ( .A(n10180), .B(n10179), .Z(n10200) );
  XOR U10955 ( .A(n10199), .B(n10200), .Z(n10188) );
  NANDN U10956 ( .A(n10182), .B(n10181), .Z(n10186) );
  OR U10957 ( .A(n10184), .B(n10183), .Z(n10185) );
  AND U10958 ( .A(n10186), .B(n10185), .Z(n10189) );
  XOR U10959 ( .A(n10188), .B(n10189), .Z(n10187) );
  XOR U10960 ( .A(n10190), .B(n10187), .Z(n10201) );
  XNOR U10961 ( .A(sreg[1408]), .B(n10201), .Z(n10202) );
  XOR U10962 ( .A(n10203), .B(n10202), .Z(c[1408]) );
  AND U10963 ( .A(b[2]), .B(a[387]), .Z(n10220) );
  AND U10964 ( .A(a[388]), .B(b[1]), .Z(n10218) );
  AND U10965 ( .A(a[386]), .B(b[3]), .Z(n10217) );
  XOR U10966 ( .A(n10218), .B(n10217), .Z(n10219) );
  XOR U10967 ( .A(n10220), .B(n10219), .Z(n10223) );
  NAND U10968 ( .A(b[0]), .B(a[389]), .Z(n10224) );
  XOR U10969 ( .A(n10223), .B(n10224), .Z(n10226) );
  OR U10970 ( .A(n10192), .B(n10191), .Z(n10196) );
  NANDN U10971 ( .A(n10194), .B(n10193), .Z(n10195) );
  NAND U10972 ( .A(n10196), .B(n10195), .Z(n10225) );
  XNOR U10973 ( .A(n10226), .B(n10225), .Z(n10211) );
  XNOR U10974 ( .A(n10211), .B(n10212), .Z(n10214) );
  XOR U10975 ( .A(n10213), .B(n10214), .Z(n10206) );
  XOR U10976 ( .A(sreg[1409]), .B(n10206), .Z(n10208) );
  NAND U10977 ( .A(sreg[1408]), .B(n10201), .Z(n10205) );
  OR U10978 ( .A(n10203), .B(n10202), .Z(n10204) );
  NAND U10979 ( .A(n10205), .B(n10204), .Z(n10207) );
  XNOR U10980 ( .A(n10208), .B(n10207), .Z(c[1409]) );
  NANDN U10981 ( .A(sreg[1409]), .B(n10206), .Z(n10210) );
  OR U10982 ( .A(n10208), .B(n10207), .Z(n10209) );
  AND U10983 ( .A(n10210), .B(n10209), .Z(n10230) );
  NANDN U10984 ( .A(n10212), .B(n10211), .Z(n10216) );
  NAND U10985 ( .A(n10214), .B(n10213), .Z(n10215) );
  NAND U10986 ( .A(n10216), .B(n10215), .Z(n10235) );
  AND U10987 ( .A(b[2]), .B(a[388]), .Z(n10241) );
  AND U10988 ( .A(a[389]), .B(b[1]), .Z(n10239) );
  AND U10989 ( .A(a[387]), .B(b[3]), .Z(n10238) );
  XOR U10990 ( .A(n10239), .B(n10238), .Z(n10240) );
  XOR U10991 ( .A(n10241), .B(n10240), .Z(n10244) );
  NAND U10992 ( .A(b[0]), .B(a[390]), .Z(n10245) );
  XOR U10993 ( .A(n10244), .B(n10245), .Z(n10247) );
  OR U10994 ( .A(n10218), .B(n10217), .Z(n10222) );
  NANDN U10995 ( .A(n10220), .B(n10219), .Z(n10221) );
  NAND U10996 ( .A(n10222), .B(n10221), .Z(n10246) );
  XNOR U10997 ( .A(n10247), .B(n10246), .Z(n10232) );
  NANDN U10998 ( .A(n10224), .B(n10223), .Z(n10228) );
  OR U10999 ( .A(n10226), .B(n10225), .Z(n10227) );
  NAND U11000 ( .A(n10228), .B(n10227), .Z(n10233) );
  XNOR U11001 ( .A(n10232), .B(n10233), .Z(n10234) );
  XNOR U11002 ( .A(n10235), .B(n10234), .Z(n10231) );
  XOR U11003 ( .A(sreg[1410]), .B(n10231), .Z(n10229) );
  XOR U11004 ( .A(n10230), .B(n10229), .Z(c[1410]) );
  NANDN U11005 ( .A(n10233), .B(n10232), .Z(n10237) );
  NAND U11006 ( .A(n10235), .B(n10234), .Z(n10236) );
  NAND U11007 ( .A(n10237), .B(n10236), .Z(n10253) );
  AND U11008 ( .A(b[2]), .B(a[389]), .Z(n10259) );
  AND U11009 ( .A(a[390]), .B(b[1]), .Z(n10257) );
  AND U11010 ( .A(a[388]), .B(b[3]), .Z(n10256) );
  XOR U11011 ( .A(n10257), .B(n10256), .Z(n10258) );
  XOR U11012 ( .A(n10259), .B(n10258), .Z(n10262) );
  NAND U11013 ( .A(b[0]), .B(a[391]), .Z(n10263) );
  XOR U11014 ( .A(n10262), .B(n10263), .Z(n10265) );
  OR U11015 ( .A(n10239), .B(n10238), .Z(n10243) );
  NANDN U11016 ( .A(n10241), .B(n10240), .Z(n10242) );
  NAND U11017 ( .A(n10243), .B(n10242), .Z(n10264) );
  XNOR U11018 ( .A(n10265), .B(n10264), .Z(n10250) );
  NANDN U11019 ( .A(n10245), .B(n10244), .Z(n10249) );
  OR U11020 ( .A(n10247), .B(n10246), .Z(n10248) );
  NAND U11021 ( .A(n10249), .B(n10248), .Z(n10251) );
  XNOR U11022 ( .A(n10250), .B(n10251), .Z(n10252) );
  XNOR U11023 ( .A(n10253), .B(n10252), .Z(n10268) );
  XNOR U11024 ( .A(n10268), .B(sreg[1411]), .Z(n10270) );
  XNOR U11025 ( .A(n10269), .B(n10270), .Z(c[1411]) );
  NANDN U11026 ( .A(n10251), .B(n10250), .Z(n10255) );
  NAND U11027 ( .A(n10253), .B(n10252), .Z(n10254) );
  NAND U11028 ( .A(n10255), .B(n10254), .Z(n10276) );
  AND U11029 ( .A(b[2]), .B(a[390]), .Z(n10282) );
  AND U11030 ( .A(a[391]), .B(b[1]), .Z(n10280) );
  AND U11031 ( .A(a[389]), .B(b[3]), .Z(n10279) );
  XOR U11032 ( .A(n10280), .B(n10279), .Z(n10281) );
  XOR U11033 ( .A(n10282), .B(n10281), .Z(n10285) );
  NAND U11034 ( .A(b[0]), .B(a[392]), .Z(n10286) );
  XOR U11035 ( .A(n10285), .B(n10286), .Z(n10288) );
  OR U11036 ( .A(n10257), .B(n10256), .Z(n10261) );
  NANDN U11037 ( .A(n10259), .B(n10258), .Z(n10260) );
  NAND U11038 ( .A(n10261), .B(n10260), .Z(n10287) );
  XNOR U11039 ( .A(n10288), .B(n10287), .Z(n10273) );
  NANDN U11040 ( .A(n10263), .B(n10262), .Z(n10267) );
  OR U11041 ( .A(n10265), .B(n10264), .Z(n10266) );
  NAND U11042 ( .A(n10267), .B(n10266), .Z(n10274) );
  XNOR U11043 ( .A(n10273), .B(n10274), .Z(n10275) );
  XNOR U11044 ( .A(n10276), .B(n10275), .Z(n10291) );
  XOR U11045 ( .A(sreg[1412]), .B(n10291), .Z(n10292) );
  NAND U11046 ( .A(n10268), .B(sreg[1411]), .Z(n10272) );
  NANDN U11047 ( .A(n10270), .B(n10269), .Z(n10271) );
  NAND U11048 ( .A(n10272), .B(n10271), .Z(n10293) );
  XOR U11049 ( .A(n10292), .B(n10293), .Z(c[1412]) );
  NANDN U11050 ( .A(n10274), .B(n10273), .Z(n10278) );
  NAND U11051 ( .A(n10276), .B(n10275), .Z(n10277) );
  NAND U11052 ( .A(n10278), .B(n10277), .Z(n10302) );
  AND U11053 ( .A(b[2]), .B(a[391]), .Z(n10308) );
  AND U11054 ( .A(a[392]), .B(b[1]), .Z(n10306) );
  AND U11055 ( .A(a[390]), .B(b[3]), .Z(n10305) );
  XOR U11056 ( .A(n10306), .B(n10305), .Z(n10307) );
  XOR U11057 ( .A(n10308), .B(n10307), .Z(n10311) );
  NAND U11058 ( .A(b[0]), .B(a[393]), .Z(n10312) );
  XOR U11059 ( .A(n10311), .B(n10312), .Z(n10314) );
  OR U11060 ( .A(n10280), .B(n10279), .Z(n10284) );
  NANDN U11061 ( .A(n10282), .B(n10281), .Z(n10283) );
  NAND U11062 ( .A(n10284), .B(n10283), .Z(n10313) );
  XNOR U11063 ( .A(n10314), .B(n10313), .Z(n10299) );
  NANDN U11064 ( .A(n10286), .B(n10285), .Z(n10290) );
  OR U11065 ( .A(n10288), .B(n10287), .Z(n10289) );
  NAND U11066 ( .A(n10290), .B(n10289), .Z(n10300) );
  XNOR U11067 ( .A(n10299), .B(n10300), .Z(n10301) );
  XOR U11068 ( .A(n10302), .B(n10301), .Z(n10298) );
  OR U11069 ( .A(n10291), .B(sreg[1412]), .Z(n10295) );
  NANDN U11070 ( .A(n10293), .B(n10292), .Z(n10294) );
  AND U11071 ( .A(n10295), .B(n10294), .Z(n10297) );
  XNOR U11072 ( .A(sreg[1413]), .B(n10297), .Z(n10296) );
  XOR U11073 ( .A(n10298), .B(n10296), .Z(c[1413]) );
  NANDN U11074 ( .A(n10300), .B(n10299), .Z(n10304) );
  NAND U11075 ( .A(n10302), .B(n10301), .Z(n10303) );
  NAND U11076 ( .A(n10304), .B(n10303), .Z(n10320) );
  AND U11077 ( .A(b[2]), .B(a[392]), .Z(n10326) );
  AND U11078 ( .A(a[393]), .B(b[1]), .Z(n10324) );
  AND U11079 ( .A(a[391]), .B(b[3]), .Z(n10323) );
  XOR U11080 ( .A(n10324), .B(n10323), .Z(n10325) );
  XOR U11081 ( .A(n10326), .B(n10325), .Z(n10329) );
  NAND U11082 ( .A(b[0]), .B(a[394]), .Z(n10330) );
  XOR U11083 ( .A(n10329), .B(n10330), .Z(n10332) );
  OR U11084 ( .A(n10306), .B(n10305), .Z(n10310) );
  NANDN U11085 ( .A(n10308), .B(n10307), .Z(n10309) );
  NAND U11086 ( .A(n10310), .B(n10309), .Z(n10331) );
  XNOR U11087 ( .A(n10332), .B(n10331), .Z(n10317) );
  NANDN U11088 ( .A(n10312), .B(n10311), .Z(n10316) );
  OR U11089 ( .A(n10314), .B(n10313), .Z(n10315) );
  NAND U11090 ( .A(n10316), .B(n10315), .Z(n10318) );
  XNOR U11091 ( .A(n10317), .B(n10318), .Z(n10319) );
  XNOR U11092 ( .A(n10320), .B(n10319), .Z(n10335) );
  XNOR U11093 ( .A(n10335), .B(sreg[1414]), .Z(n10336) );
  XOR U11094 ( .A(n10337), .B(n10336), .Z(c[1414]) );
  NANDN U11095 ( .A(n10318), .B(n10317), .Z(n10322) );
  NAND U11096 ( .A(n10320), .B(n10319), .Z(n10321) );
  NAND U11097 ( .A(n10322), .B(n10321), .Z(n10348) );
  AND U11098 ( .A(b[2]), .B(a[393]), .Z(n10354) );
  AND U11099 ( .A(a[394]), .B(b[1]), .Z(n10352) );
  AND U11100 ( .A(a[392]), .B(b[3]), .Z(n10351) );
  XOR U11101 ( .A(n10352), .B(n10351), .Z(n10353) );
  XOR U11102 ( .A(n10354), .B(n10353), .Z(n10357) );
  NAND U11103 ( .A(b[0]), .B(a[395]), .Z(n10358) );
  XOR U11104 ( .A(n10357), .B(n10358), .Z(n10360) );
  OR U11105 ( .A(n10324), .B(n10323), .Z(n10328) );
  NANDN U11106 ( .A(n10326), .B(n10325), .Z(n10327) );
  NAND U11107 ( .A(n10328), .B(n10327), .Z(n10359) );
  XNOR U11108 ( .A(n10360), .B(n10359), .Z(n10345) );
  NANDN U11109 ( .A(n10330), .B(n10329), .Z(n10334) );
  OR U11110 ( .A(n10332), .B(n10331), .Z(n10333) );
  NAND U11111 ( .A(n10334), .B(n10333), .Z(n10346) );
  XNOR U11112 ( .A(n10345), .B(n10346), .Z(n10347) );
  XNOR U11113 ( .A(n10348), .B(n10347), .Z(n10340) );
  XOR U11114 ( .A(sreg[1415]), .B(n10340), .Z(n10341) );
  NAND U11115 ( .A(n10335), .B(sreg[1414]), .Z(n10339) );
  OR U11116 ( .A(n10337), .B(n10336), .Z(n10338) );
  NAND U11117 ( .A(n10339), .B(n10338), .Z(n10342) );
  XOR U11118 ( .A(n10341), .B(n10342), .Z(c[1415]) );
  OR U11119 ( .A(n10340), .B(sreg[1415]), .Z(n10344) );
  NANDN U11120 ( .A(n10342), .B(n10341), .Z(n10343) );
  AND U11121 ( .A(n10344), .B(n10343), .Z(n10364) );
  NANDN U11122 ( .A(n10346), .B(n10345), .Z(n10350) );
  NAND U11123 ( .A(n10348), .B(n10347), .Z(n10349) );
  NAND U11124 ( .A(n10350), .B(n10349), .Z(n10369) );
  AND U11125 ( .A(b[2]), .B(a[394]), .Z(n10375) );
  AND U11126 ( .A(a[395]), .B(b[1]), .Z(n10373) );
  AND U11127 ( .A(a[393]), .B(b[3]), .Z(n10372) );
  XOR U11128 ( .A(n10373), .B(n10372), .Z(n10374) );
  XOR U11129 ( .A(n10375), .B(n10374), .Z(n10378) );
  NAND U11130 ( .A(b[0]), .B(a[396]), .Z(n10379) );
  XOR U11131 ( .A(n10378), .B(n10379), .Z(n10381) );
  OR U11132 ( .A(n10352), .B(n10351), .Z(n10356) );
  NANDN U11133 ( .A(n10354), .B(n10353), .Z(n10355) );
  NAND U11134 ( .A(n10356), .B(n10355), .Z(n10380) );
  XNOR U11135 ( .A(n10381), .B(n10380), .Z(n10366) );
  NANDN U11136 ( .A(n10358), .B(n10357), .Z(n10362) );
  OR U11137 ( .A(n10360), .B(n10359), .Z(n10361) );
  NAND U11138 ( .A(n10362), .B(n10361), .Z(n10367) );
  XNOR U11139 ( .A(n10366), .B(n10367), .Z(n10368) );
  XNOR U11140 ( .A(n10369), .B(n10368), .Z(n10365) );
  XOR U11141 ( .A(sreg[1416]), .B(n10365), .Z(n10363) );
  XOR U11142 ( .A(n10364), .B(n10363), .Z(c[1416]) );
  NANDN U11143 ( .A(n10367), .B(n10366), .Z(n10371) );
  NAND U11144 ( .A(n10369), .B(n10368), .Z(n10370) );
  NAND U11145 ( .A(n10371), .B(n10370), .Z(n10387) );
  AND U11146 ( .A(b[2]), .B(a[395]), .Z(n10393) );
  AND U11147 ( .A(a[396]), .B(b[1]), .Z(n10391) );
  AND U11148 ( .A(a[394]), .B(b[3]), .Z(n10390) );
  XOR U11149 ( .A(n10391), .B(n10390), .Z(n10392) );
  XOR U11150 ( .A(n10393), .B(n10392), .Z(n10396) );
  NAND U11151 ( .A(b[0]), .B(a[397]), .Z(n10397) );
  XOR U11152 ( .A(n10396), .B(n10397), .Z(n10399) );
  OR U11153 ( .A(n10373), .B(n10372), .Z(n10377) );
  NANDN U11154 ( .A(n10375), .B(n10374), .Z(n10376) );
  NAND U11155 ( .A(n10377), .B(n10376), .Z(n10398) );
  XNOR U11156 ( .A(n10399), .B(n10398), .Z(n10384) );
  NANDN U11157 ( .A(n10379), .B(n10378), .Z(n10383) );
  OR U11158 ( .A(n10381), .B(n10380), .Z(n10382) );
  NAND U11159 ( .A(n10383), .B(n10382), .Z(n10385) );
  XNOR U11160 ( .A(n10384), .B(n10385), .Z(n10386) );
  XNOR U11161 ( .A(n10387), .B(n10386), .Z(n10402) );
  XNOR U11162 ( .A(n10402), .B(sreg[1417]), .Z(n10404) );
  XNOR U11163 ( .A(n10403), .B(n10404), .Z(c[1417]) );
  NANDN U11164 ( .A(n10385), .B(n10384), .Z(n10389) );
  NAND U11165 ( .A(n10387), .B(n10386), .Z(n10388) );
  NAND U11166 ( .A(n10389), .B(n10388), .Z(n10410) );
  AND U11167 ( .A(b[2]), .B(a[396]), .Z(n10416) );
  AND U11168 ( .A(a[397]), .B(b[1]), .Z(n10414) );
  AND U11169 ( .A(a[395]), .B(b[3]), .Z(n10413) );
  XOR U11170 ( .A(n10414), .B(n10413), .Z(n10415) );
  XOR U11171 ( .A(n10416), .B(n10415), .Z(n10419) );
  NAND U11172 ( .A(b[0]), .B(a[398]), .Z(n10420) );
  XOR U11173 ( .A(n10419), .B(n10420), .Z(n10422) );
  OR U11174 ( .A(n10391), .B(n10390), .Z(n10395) );
  NANDN U11175 ( .A(n10393), .B(n10392), .Z(n10394) );
  NAND U11176 ( .A(n10395), .B(n10394), .Z(n10421) );
  XNOR U11177 ( .A(n10422), .B(n10421), .Z(n10407) );
  NANDN U11178 ( .A(n10397), .B(n10396), .Z(n10401) );
  OR U11179 ( .A(n10399), .B(n10398), .Z(n10400) );
  NAND U11180 ( .A(n10401), .B(n10400), .Z(n10408) );
  XNOR U11181 ( .A(n10407), .B(n10408), .Z(n10409) );
  XNOR U11182 ( .A(n10410), .B(n10409), .Z(n10425) );
  XNOR U11183 ( .A(n10425), .B(sreg[1418]), .Z(n10427) );
  NAND U11184 ( .A(n10402), .B(sreg[1417]), .Z(n10406) );
  NANDN U11185 ( .A(n10404), .B(n10403), .Z(n10405) );
  AND U11186 ( .A(n10406), .B(n10405), .Z(n10426) );
  XOR U11187 ( .A(n10427), .B(n10426), .Z(c[1418]) );
  NANDN U11188 ( .A(n10408), .B(n10407), .Z(n10412) );
  NAND U11189 ( .A(n10410), .B(n10409), .Z(n10411) );
  NAND U11190 ( .A(n10412), .B(n10411), .Z(n10433) );
  AND U11191 ( .A(b[2]), .B(a[397]), .Z(n10439) );
  AND U11192 ( .A(a[398]), .B(b[1]), .Z(n10437) );
  AND U11193 ( .A(a[396]), .B(b[3]), .Z(n10436) );
  XOR U11194 ( .A(n10437), .B(n10436), .Z(n10438) );
  XOR U11195 ( .A(n10439), .B(n10438), .Z(n10442) );
  NAND U11196 ( .A(b[0]), .B(a[399]), .Z(n10443) );
  XOR U11197 ( .A(n10442), .B(n10443), .Z(n10445) );
  OR U11198 ( .A(n10414), .B(n10413), .Z(n10418) );
  NANDN U11199 ( .A(n10416), .B(n10415), .Z(n10417) );
  NAND U11200 ( .A(n10418), .B(n10417), .Z(n10444) );
  XNOR U11201 ( .A(n10445), .B(n10444), .Z(n10430) );
  NANDN U11202 ( .A(n10420), .B(n10419), .Z(n10424) );
  OR U11203 ( .A(n10422), .B(n10421), .Z(n10423) );
  NAND U11204 ( .A(n10424), .B(n10423), .Z(n10431) );
  XNOR U11205 ( .A(n10430), .B(n10431), .Z(n10432) );
  XNOR U11206 ( .A(n10433), .B(n10432), .Z(n10448) );
  XNOR U11207 ( .A(n10448), .B(sreg[1419]), .Z(n10450) );
  NAND U11208 ( .A(n10425), .B(sreg[1418]), .Z(n10429) );
  OR U11209 ( .A(n10427), .B(n10426), .Z(n10428) );
  AND U11210 ( .A(n10429), .B(n10428), .Z(n10449) );
  XOR U11211 ( .A(n10450), .B(n10449), .Z(c[1419]) );
  NANDN U11212 ( .A(n10431), .B(n10430), .Z(n10435) );
  NAND U11213 ( .A(n10433), .B(n10432), .Z(n10434) );
  NAND U11214 ( .A(n10435), .B(n10434), .Z(n10459) );
  AND U11215 ( .A(b[2]), .B(a[398]), .Z(n10465) );
  AND U11216 ( .A(a[399]), .B(b[1]), .Z(n10463) );
  AND U11217 ( .A(a[397]), .B(b[3]), .Z(n10462) );
  XOR U11218 ( .A(n10463), .B(n10462), .Z(n10464) );
  XOR U11219 ( .A(n10465), .B(n10464), .Z(n10468) );
  NAND U11220 ( .A(b[0]), .B(a[400]), .Z(n10469) );
  XOR U11221 ( .A(n10468), .B(n10469), .Z(n10471) );
  OR U11222 ( .A(n10437), .B(n10436), .Z(n10441) );
  NANDN U11223 ( .A(n10439), .B(n10438), .Z(n10440) );
  NAND U11224 ( .A(n10441), .B(n10440), .Z(n10470) );
  XNOR U11225 ( .A(n10471), .B(n10470), .Z(n10456) );
  NANDN U11226 ( .A(n10443), .B(n10442), .Z(n10447) );
  OR U11227 ( .A(n10445), .B(n10444), .Z(n10446) );
  NAND U11228 ( .A(n10447), .B(n10446), .Z(n10457) );
  XNOR U11229 ( .A(n10456), .B(n10457), .Z(n10458) );
  XOR U11230 ( .A(n10459), .B(n10458), .Z(n10455) );
  NAND U11231 ( .A(n10448), .B(sreg[1419]), .Z(n10452) );
  OR U11232 ( .A(n10450), .B(n10449), .Z(n10451) );
  NAND U11233 ( .A(n10452), .B(n10451), .Z(n10454) );
  XNOR U11234 ( .A(sreg[1420]), .B(n10454), .Z(n10453) );
  XOR U11235 ( .A(n10455), .B(n10453), .Z(c[1420]) );
  NANDN U11236 ( .A(n10457), .B(n10456), .Z(n10461) );
  NAND U11237 ( .A(n10459), .B(n10458), .Z(n10460) );
  NAND U11238 ( .A(n10461), .B(n10460), .Z(n10477) );
  AND U11239 ( .A(b[2]), .B(a[399]), .Z(n10483) );
  AND U11240 ( .A(a[400]), .B(b[1]), .Z(n10481) );
  AND U11241 ( .A(a[398]), .B(b[3]), .Z(n10480) );
  XOR U11242 ( .A(n10481), .B(n10480), .Z(n10482) );
  XOR U11243 ( .A(n10483), .B(n10482), .Z(n10486) );
  NAND U11244 ( .A(b[0]), .B(a[401]), .Z(n10487) );
  XOR U11245 ( .A(n10486), .B(n10487), .Z(n10489) );
  OR U11246 ( .A(n10463), .B(n10462), .Z(n10467) );
  NANDN U11247 ( .A(n10465), .B(n10464), .Z(n10466) );
  NAND U11248 ( .A(n10467), .B(n10466), .Z(n10488) );
  XNOR U11249 ( .A(n10489), .B(n10488), .Z(n10474) );
  NANDN U11250 ( .A(n10469), .B(n10468), .Z(n10473) );
  OR U11251 ( .A(n10471), .B(n10470), .Z(n10472) );
  NAND U11252 ( .A(n10473), .B(n10472), .Z(n10475) );
  XNOR U11253 ( .A(n10474), .B(n10475), .Z(n10476) );
  XNOR U11254 ( .A(n10477), .B(n10476), .Z(n10492) );
  XNOR U11255 ( .A(n10492), .B(sreg[1421]), .Z(n10493) );
  XOR U11256 ( .A(n10494), .B(n10493), .Z(c[1421]) );
  NANDN U11257 ( .A(n10475), .B(n10474), .Z(n10479) );
  NAND U11258 ( .A(n10477), .B(n10476), .Z(n10478) );
  NAND U11259 ( .A(n10479), .B(n10478), .Z(n10503) );
  AND U11260 ( .A(b[2]), .B(a[400]), .Z(n10509) );
  AND U11261 ( .A(a[401]), .B(b[1]), .Z(n10507) );
  AND U11262 ( .A(a[399]), .B(b[3]), .Z(n10506) );
  XOR U11263 ( .A(n10507), .B(n10506), .Z(n10508) );
  XOR U11264 ( .A(n10509), .B(n10508), .Z(n10512) );
  NAND U11265 ( .A(b[0]), .B(a[402]), .Z(n10513) );
  XOR U11266 ( .A(n10512), .B(n10513), .Z(n10515) );
  OR U11267 ( .A(n10481), .B(n10480), .Z(n10485) );
  NANDN U11268 ( .A(n10483), .B(n10482), .Z(n10484) );
  NAND U11269 ( .A(n10485), .B(n10484), .Z(n10514) );
  XNOR U11270 ( .A(n10515), .B(n10514), .Z(n10500) );
  NANDN U11271 ( .A(n10487), .B(n10486), .Z(n10491) );
  OR U11272 ( .A(n10489), .B(n10488), .Z(n10490) );
  NAND U11273 ( .A(n10491), .B(n10490), .Z(n10501) );
  XNOR U11274 ( .A(n10500), .B(n10501), .Z(n10502) );
  XOR U11275 ( .A(n10503), .B(n10502), .Z(n10499) );
  NAND U11276 ( .A(n10492), .B(sreg[1421]), .Z(n10496) );
  OR U11277 ( .A(n10494), .B(n10493), .Z(n10495) );
  NAND U11278 ( .A(n10496), .B(n10495), .Z(n10498) );
  XNOR U11279 ( .A(sreg[1422]), .B(n10498), .Z(n10497) );
  XOR U11280 ( .A(n10499), .B(n10497), .Z(c[1422]) );
  NANDN U11281 ( .A(n10501), .B(n10500), .Z(n10505) );
  NAND U11282 ( .A(n10503), .B(n10502), .Z(n10504) );
  NAND U11283 ( .A(n10505), .B(n10504), .Z(n10521) );
  AND U11284 ( .A(b[2]), .B(a[401]), .Z(n10527) );
  AND U11285 ( .A(a[402]), .B(b[1]), .Z(n10525) );
  AND U11286 ( .A(a[400]), .B(b[3]), .Z(n10524) );
  XOR U11287 ( .A(n10525), .B(n10524), .Z(n10526) );
  XOR U11288 ( .A(n10527), .B(n10526), .Z(n10530) );
  NAND U11289 ( .A(b[0]), .B(a[403]), .Z(n10531) );
  XOR U11290 ( .A(n10530), .B(n10531), .Z(n10533) );
  OR U11291 ( .A(n10507), .B(n10506), .Z(n10511) );
  NANDN U11292 ( .A(n10509), .B(n10508), .Z(n10510) );
  NAND U11293 ( .A(n10511), .B(n10510), .Z(n10532) );
  XNOR U11294 ( .A(n10533), .B(n10532), .Z(n10518) );
  NANDN U11295 ( .A(n10513), .B(n10512), .Z(n10517) );
  OR U11296 ( .A(n10515), .B(n10514), .Z(n10516) );
  NAND U11297 ( .A(n10517), .B(n10516), .Z(n10519) );
  XNOR U11298 ( .A(n10518), .B(n10519), .Z(n10520) );
  XNOR U11299 ( .A(n10521), .B(n10520), .Z(n10536) );
  XOR U11300 ( .A(sreg[1423]), .B(n10536), .Z(n10538) );
  XNOR U11301 ( .A(n10537), .B(n10538), .Z(c[1423]) );
  NANDN U11302 ( .A(n10519), .B(n10518), .Z(n10523) );
  NAND U11303 ( .A(n10521), .B(n10520), .Z(n10522) );
  NAND U11304 ( .A(n10523), .B(n10522), .Z(n10547) );
  AND U11305 ( .A(b[2]), .B(a[402]), .Z(n10559) );
  AND U11306 ( .A(a[403]), .B(b[1]), .Z(n10557) );
  AND U11307 ( .A(a[401]), .B(b[3]), .Z(n10556) );
  XOR U11308 ( .A(n10557), .B(n10556), .Z(n10558) );
  XOR U11309 ( .A(n10559), .B(n10558), .Z(n10550) );
  NAND U11310 ( .A(b[0]), .B(a[404]), .Z(n10551) );
  XOR U11311 ( .A(n10550), .B(n10551), .Z(n10553) );
  OR U11312 ( .A(n10525), .B(n10524), .Z(n10529) );
  NANDN U11313 ( .A(n10527), .B(n10526), .Z(n10528) );
  NAND U11314 ( .A(n10529), .B(n10528), .Z(n10552) );
  XNOR U11315 ( .A(n10553), .B(n10552), .Z(n10544) );
  NANDN U11316 ( .A(n10531), .B(n10530), .Z(n10535) );
  OR U11317 ( .A(n10533), .B(n10532), .Z(n10534) );
  NAND U11318 ( .A(n10535), .B(n10534), .Z(n10545) );
  XNOR U11319 ( .A(n10544), .B(n10545), .Z(n10546) );
  XOR U11320 ( .A(n10547), .B(n10546), .Z(n10543) );
  OR U11321 ( .A(n10536), .B(sreg[1423]), .Z(n10540) );
  NAND U11322 ( .A(n10538), .B(n10537), .Z(n10539) );
  AND U11323 ( .A(n10540), .B(n10539), .Z(n10542) );
  XNOR U11324 ( .A(sreg[1424]), .B(n10542), .Z(n10541) );
  XOR U11325 ( .A(n10543), .B(n10541), .Z(c[1424]) );
  NANDN U11326 ( .A(n10545), .B(n10544), .Z(n10549) );
  NAND U11327 ( .A(n10547), .B(n10546), .Z(n10548) );
  NAND U11328 ( .A(n10549), .B(n10548), .Z(n10577) );
  NANDN U11329 ( .A(n10551), .B(n10550), .Z(n10555) );
  OR U11330 ( .A(n10553), .B(n10552), .Z(n10554) );
  NAND U11331 ( .A(n10555), .B(n10554), .Z(n10574) );
  AND U11332 ( .A(b[2]), .B(a[403]), .Z(n10565) );
  AND U11333 ( .A(a[404]), .B(b[1]), .Z(n10563) );
  AND U11334 ( .A(a[402]), .B(b[3]), .Z(n10562) );
  XOR U11335 ( .A(n10563), .B(n10562), .Z(n10564) );
  XOR U11336 ( .A(n10565), .B(n10564), .Z(n10568) );
  NAND U11337 ( .A(b[0]), .B(a[405]), .Z(n10569) );
  XNOR U11338 ( .A(n10568), .B(n10569), .Z(n10570) );
  OR U11339 ( .A(n10557), .B(n10556), .Z(n10561) );
  NANDN U11340 ( .A(n10559), .B(n10558), .Z(n10560) );
  AND U11341 ( .A(n10561), .B(n10560), .Z(n10571) );
  XNOR U11342 ( .A(n10570), .B(n10571), .Z(n10575) );
  XNOR U11343 ( .A(n10574), .B(n10575), .Z(n10576) );
  XNOR U11344 ( .A(n10577), .B(n10576), .Z(n10580) );
  XNOR U11345 ( .A(sreg[1425]), .B(n10580), .Z(n10581) );
  XOR U11346 ( .A(n10582), .B(n10581), .Z(c[1425]) );
  AND U11347 ( .A(b[2]), .B(a[404]), .Z(n10595) );
  AND U11348 ( .A(a[405]), .B(b[1]), .Z(n10593) );
  AND U11349 ( .A(a[403]), .B(b[3]), .Z(n10592) );
  XOR U11350 ( .A(n10593), .B(n10592), .Z(n10594) );
  XOR U11351 ( .A(n10595), .B(n10594), .Z(n10598) );
  NAND U11352 ( .A(b[0]), .B(a[406]), .Z(n10599) );
  XOR U11353 ( .A(n10598), .B(n10599), .Z(n10601) );
  OR U11354 ( .A(n10563), .B(n10562), .Z(n10567) );
  NANDN U11355 ( .A(n10565), .B(n10564), .Z(n10566) );
  NAND U11356 ( .A(n10567), .B(n10566), .Z(n10600) );
  XNOR U11357 ( .A(n10601), .B(n10600), .Z(n10586) );
  NANDN U11358 ( .A(n10569), .B(n10568), .Z(n10573) );
  NAND U11359 ( .A(n10571), .B(n10570), .Z(n10572) );
  NAND U11360 ( .A(n10573), .B(n10572), .Z(n10587) );
  XNOR U11361 ( .A(n10586), .B(n10587), .Z(n10588) );
  NANDN U11362 ( .A(n10575), .B(n10574), .Z(n10579) );
  NANDN U11363 ( .A(n10577), .B(n10576), .Z(n10578) );
  NAND U11364 ( .A(n10579), .B(n10578), .Z(n10589) );
  XOR U11365 ( .A(n10588), .B(n10589), .Z(n10605) );
  NAND U11366 ( .A(sreg[1425]), .B(n10580), .Z(n10584) );
  OR U11367 ( .A(n10582), .B(n10581), .Z(n10583) );
  NAND U11368 ( .A(n10584), .B(n10583), .Z(n10604) );
  XNOR U11369 ( .A(sreg[1426]), .B(n10604), .Z(n10585) );
  XNOR U11370 ( .A(n10605), .B(n10585), .Z(c[1426]) );
  NANDN U11371 ( .A(n10587), .B(n10586), .Z(n10591) );
  NANDN U11372 ( .A(n10589), .B(n10588), .Z(n10590) );
  NAND U11373 ( .A(n10591), .B(n10590), .Z(n10624) );
  AND U11374 ( .A(b[2]), .B(a[405]), .Z(n10618) );
  AND U11375 ( .A(a[406]), .B(b[1]), .Z(n10616) );
  AND U11376 ( .A(a[404]), .B(b[3]), .Z(n10615) );
  XOR U11377 ( .A(n10616), .B(n10615), .Z(n10617) );
  XOR U11378 ( .A(n10618), .B(n10617), .Z(n10609) );
  NAND U11379 ( .A(b[0]), .B(a[407]), .Z(n10610) );
  XOR U11380 ( .A(n10609), .B(n10610), .Z(n10612) );
  OR U11381 ( .A(n10593), .B(n10592), .Z(n10597) );
  NANDN U11382 ( .A(n10595), .B(n10594), .Z(n10596) );
  NAND U11383 ( .A(n10597), .B(n10596), .Z(n10611) );
  XNOR U11384 ( .A(n10612), .B(n10611), .Z(n10621) );
  NANDN U11385 ( .A(n10599), .B(n10598), .Z(n10603) );
  OR U11386 ( .A(n10601), .B(n10600), .Z(n10602) );
  NAND U11387 ( .A(n10603), .B(n10602), .Z(n10622) );
  XNOR U11388 ( .A(n10621), .B(n10622), .Z(n10623) );
  XOR U11389 ( .A(n10624), .B(n10623), .Z(n10608) );
  XNOR U11390 ( .A(sreg[1427]), .B(n10607), .Z(n10606) );
  XOR U11391 ( .A(n10608), .B(n10606), .Z(c[1427]) );
  NANDN U11392 ( .A(n10610), .B(n10609), .Z(n10614) );
  OR U11393 ( .A(n10612), .B(n10611), .Z(n10613) );
  NAND U11394 ( .A(n10614), .B(n10613), .Z(n10639) );
  AND U11395 ( .A(b[2]), .B(a[406]), .Z(n10630) );
  AND U11396 ( .A(a[407]), .B(b[1]), .Z(n10628) );
  AND U11397 ( .A(a[405]), .B(b[3]), .Z(n10627) );
  XOR U11398 ( .A(n10628), .B(n10627), .Z(n10629) );
  XOR U11399 ( .A(n10630), .B(n10629), .Z(n10633) );
  NAND U11400 ( .A(b[0]), .B(a[408]), .Z(n10634) );
  XNOR U11401 ( .A(n10633), .B(n10634), .Z(n10635) );
  OR U11402 ( .A(n10616), .B(n10615), .Z(n10620) );
  NANDN U11403 ( .A(n10618), .B(n10617), .Z(n10619) );
  AND U11404 ( .A(n10620), .B(n10619), .Z(n10636) );
  XNOR U11405 ( .A(n10635), .B(n10636), .Z(n10640) );
  XNOR U11406 ( .A(n10639), .B(n10640), .Z(n10641) );
  NANDN U11407 ( .A(n10622), .B(n10621), .Z(n10626) );
  NAND U11408 ( .A(n10624), .B(n10623), .Z(n10625) );
  AND U11409 ( .A(n10626), .B(n10625), .Z(n10642) );
  XOR U11410 ( .A(n10641), .B(n10642), .Z(n10645) );
  XNOR U11411 ( .A(sreg[1428]), .B(n10645), .Z(n10646) );
  XOR U11412 ( .A(n10647), .B(n10646), .Z(c[1428]) );
  AND U11413 ( .A(b[2]), .B(a[407]), .Z(n10662) );
  AND U11414 ( .A(a[408]), .B(b[1]), .Z(n10660) );
  AND U11415 ( .A(a[406]), .B(b[3]), .Z(n10659) );
  XOR U11416 ( .A(n10660), .B(n10659), .Z(n10661) );
  XOR U11417 ( .A(n10662), .B(n10661), .Z(n10665) );
  NAND U11418 ( .A(b[0]), .B(a[409]), .Z(n10666) );
  XOR U11419 ( .A(n10665), .B(n10666), .Z(n10668) );
  OR U11420 ( .A(n10628), .B(n10627), .Z(n10632) );
  NANDN U11421 ( .A(n10630), .B(n10629), .Z(n10631) );
  NAND U11422 ( .A(n10632), .B(n10631), .Z(n10667) );
  XNOR U11423 ( .A(n10668), .B(n10667), .Z(n10653) );
  NANDN U11424 ( .A(n10634), .B(n10633), .Z(n10638) );
  NAND U11425 ( .A(n10636), .B(n10635), .Z(n10637) );
  NAND U11426 ( .A(n10638), .B(n10637), .Z(n10654) );
  XNOR U11427 ( .A(n10653), .B(n10654), .Z(n10655) );
  NANDN U11428 ( .A(n10640), .B(n10639), .Z(n10644) );
  NAND U11429 ( .A(n10642), .B(n10641), .Z(n10643) );
  AND U11430 ( .A(n10644), .B(n10643), .Z(n10656) );
  XNOR U11431 ( .A(n10655), .B(n10656), .Z(n10652) );
  NAND U11432 ( .A(sreg[1428]), .B(n10645), .Z(n10649) );
  OR U11433 ( .A(n10647), .B(n10646), .Z(n10648) );
  AND U11434 ( .A(n10649), .B(n10648), .Z(n10651) );
  XNOR U11435 ( .A(n10651), .B(sreg[1429]), .Z(n10650) );
  XOR U11436 ( .A(n10652), .B(n10650), .Z(c[1429]) );
  NANDN U11437 ( .A(n10654), .B(n10653), .Z(n10658) );
  NAND U11438 ( .A(n10656), .B(n10655), .Z(n10657) );
  NAND U11439 ( .A(n10658), .B(n10657), .Z(n10686) );
  AND U11440 ( .A(b[2]), .B(a[408]), .Z(n10680) );
  AND U11441 ( .A(a[409]), .B(b[1]), .Z(n10678) );
  AND U11442 ( .A(a[407]), .B(b[3]), .Z(n10677) );
  XOR U11443 ( .A(n10678), .B(n10677), .Z(n10679) );
  XOR U11444 ( .A(n10680), .B(n10679), .Z(n10671) );
  NAND U11445 ( .A(b[0]), .B(a[410]), .Z(n10672) );
  XOR U11446 ( .A(n10671), .B(n10672), .Z(n10674) );
  OR U11447 ( .A(n10660), .B(n10659), .Z(n10664) );
  NANDN U11448 ( .A(n10662), .B(n10661), .Z(n10663) );
  NAND U11449 ( .A(n10664), .B(n10663), .Z(n10673) );
  XNOR U11450 ( .A(n10674), .B(n10673), .Z(n10683) );
  NANDN U11451 ( .A(n10666), .B(n10665), .Z(n10670) );
  OR U11452 ( .A(n10668), .B(n10667), .Z(n10669) );
  NAND U11453 ( .A(n10670), .B(n10669), .Z(n10684) );
  XNOR U11454 ( .A(n10683), .B(n10684), .Z(n10685) );
  XNOR U11455 ( .A(n10686), .B(n10685), .Z(n10689) );
  XNOR U11456 ( .A(n10689), .B(sreg[1430]), .Z(n10691) );
  XNOR U11457 ( .A(n10690), .B(n10691), .Z(c[1430]) );
  NANDN U11458 ( .A(n10672), .B(n10671), .Z(n10676) );
  OR U11459 ( .A(n10674), .B(n10673), .Z(n10675) );
  NAND U11460 ( .A(n10676), .B(n10675), .Z(n10706) );
  AND U11461 ( .A(b[2]), .B(a[409]), .Z(n10697) );
  AND U11462 ( .A(a[410]), .B(b[1]), .Z(n10695) );
  AND U11463 ( .A(a[408]), .B(b[3]), .Z(n10694) );
  XOR U11464 ( .A(n10695), .B(n10694), .Z(n10696) );
  XOR U11465 ( .A(n10697), .B(n10696), .Z(n10700) );
  NAND U11466 ( .A(b[0]), .B(a[411]), .Z(n10701) );
  XNOR U11467 ( .A(n10700), .B(n10701), .Z(n10702) );
  OR U11468 ( .A(n10678), .B(n10677), .Z(n10682) );
  NANDN U11469 ( .A(n10680), .B(n10679), .Z(n10681) );
  AND U11470 ( .A(n10682), .B(n10681), .Z(n10703) );
  XNOR U11471 ( .A(n10702), .B(n10703), .Z(n10707) );
  XNOR U11472 ( .A(n10706), .B(n10707), .Z(n10708) );
  NANDN U11473 ( .A(n10684), .B(n10683), .Z(n10688) );
  NAND U11474 ( .A(n10686), .B(n10685), .Z(n10687) );
  NAND U11475 ( .A(n10688), .B(n10687), .Z(n10709) );
  XNOR U11476 ( .A(n10708), .B(n10709), .Z(n10712) );
  XOR U11477 ( .A(sreg[1431]), .B(n10712), .Z(n10713) );
  NAND U11478 ( .A(n10689), .B(sreg[1430]), .Z(n10693) );
  NANDN U11479 ( .A(n10691), .B(n10690), .Z(n10692) );
  NAND U11480 ( .A(n10693), .B(n10692), .Z(n10714) );
  XOR U11481 ( .A(n10713), .B(n10714), .Z(c[1431]) );
  AND U11482 ( .A(b[2]), .B(a[410]), .Z(n10729) );
  AND U11483 ( .A(a[411]), .B(b[1]), .Z(n10727) );
  AND U11484 ( .A(a[409]), .B(b[3]), .Z(n10726) );
  XOR U11485 ( .A(n10727), .B(n10726), .Z(n10728) );
  XOR U11486 ( .A(n10729), .B(n10728), .Z(n10732) );
  NAND U11487 ( .A(b[0]), .B(a[412]), .Z(n10733) );
  XOR U11488 ( .A(n10732), .B(n10733), .Z(n10735) );
  OR U11489 ( .A(n10695), .B(n10694), .Z(n10699) );
  NANDN U11490 ( .A(n10697), .B(n10696), .Z(n10698) );
  NAND U11491 ( .A(n10699), .B(n10698), .Z(n10734) );
  XNOR U11492 ( .A(n10735), .B(n10734), .Z(n10720) );
  NANDN U11493 ( .A(n10701), .B(n10700), .Z(n10705) );
  NAND U11494 ( .A(n10703), .B(n10702), .Z(n10704) );
  NAND U11495 ( .A(n10705), .B(n10704), .Z(n10721) );
  XNOR U11496 ( .A(n10720), .B(n10721), .Z(n10722) );
  NANDN U11497 ( .A(n10707), .B(n10706), .Z(n10711) );
  NANDN U11498 ( .A(n10709), .B(n10708), .Z(n10710) );
  NAND U11499 ( .A(n10711), .B(n10710), .Z(n10723) );
  XOR U11500 ( .A(n10722), .B(n10723), .Z(n10719) );
  OR U11501 ( .A(n10712), .B(sreg[1431]), .Z(n10716) );
  NANDN U11502 ( .A(n10714), .B(n10713), .Z(n10715) );
  AND U11503 ( .A(n10716), .B(n10715), .Z(n10718) );
  XNOR U11504 ( .A(sreg[1432]), .B(n10718), .Z(n10717) );
  XNOR U11505 ( .A(n10719), .B(n10717), .Z(c[1432]) );
  NANDN U11506 ( .A(n10721), .B(n10720), .Z(n10725) );
  NANDN U11507 ( .A(n10723), .B(n10722), .Z(n10724) );
  NAND U11508 ( .A(n10725), .B(n10724), .Z(n10753) );
  AND U11509 ( .A(b[2]), .B(a[411]), .Z(n10747) );
  AND U11510 ( .A(a[412]), .B(b[1]), .Z(n10745) );
  AND U11511 ( .A(a[410]), .B(b[3]), .Z(n10744) );
  XOR U11512 ( .A(n10745), .B(n10744), .Z(n10746) );
  XOR U11513 ( .A(n10747), .B(n10746), .Z(n10738) );
  NAND U11514 ( .A(b[0]), .B(a[413]), .Z(n10739) );
  XOR U11515 ( .A(n10738), .B(n10739), .Z(n10741) );
  OR U11516 ( .A(n10727), .B(n10726), .Z(n10731) );
  NANDN U11517 ( .A(n10729), .B(n10728), .Z(n10730) );
  NAND U11518 ( .A(n10731), .B(n10730), .Z(n10740) );
  XNOR U11519 ( .A(n10741), .B(n10740), .Z(n10750) );
  NANDN U11520 ( .A(n10733), .B(n10732), .Z(n10737) );
  OR U11521 ( .A(n10735), .B(n10734), .Z(n10736) );
  NAND U11522 ( .A(n10737), .B(n10736), .Z(n10751) );
  XNOR U11523 ( .A(n10750), .B(n10751), .Z(n10752) );
  XNOR U11524 ( .A(n10753), .B(n10752), .Z(n10756) );
  XNOR U11525 ( .A(n10756), .B(sreg[1433]), .Z(n10757) );
  XOR U11526 ( .A(n10758), .B(n10757), .Z(c[1433]) );
  NANDN U11527 ( .A(n10739), .B(n10738), .Z(n10743) );
  OR U11528 ( .A(n10741), .B(n10740), .Z(n10742) );
  NAND U11529 ( .A(n10743), .B(n10742), .Z(n10776) );
  AND U11530 ( .A(b[2]), .B(a[412]), .Z(n10767) );
  AND U11531 ( .A(a[413]), .B(b[1]), .Z(n10765) );
  AND U11532 ( .A(a[411]), .B(b[3]), .Z(n10764) );
  XOR U11533 ( .A(n10765), .B(n10764), .Z(n10766) );
  XOR U11534 ( .A(n10767), .B(n10766), .Z(n10770) );
  NAND U11535 ( .A(b[0]), .B(a[414]), .Z(n10771) );
  XNOR U11536 ( .A(n10770), .B(n10771), .Z(n10772) );
  OR U11537 ( .A(n10745), .B(n10744), .Z(n10749) );
  NANDN U11538 ( .A(n10747), .B(n10746), .Z(n10748) );
  AND U11539 ( .A(n10749), .B(n10748), .Z(n10773) );
  XNOR U11540 ( .A(n10772), .B(n10773), .Z(n10777) );
  XNOR U11541 ( .A(n10776), .B(n10777), .Z(n10778) );
  NANDN U11542 ( .A(n10751), .B(n10750), .Z(n10755) );
  NAND U11543 ( .A(n10753), .B(n10752), .Z(n10754) );
  NAND U11544 ( .A(n10755), .B(n10754), .Z(n10779) );
  XOR U11545 ( .A(n10778), .B(n10779), .Z(n10763) );
  NAND U11546 ( .A(n10756), .B(sreg[1433]), .Z(n10760) );
  OR U11547 ( .A(n10758), .B(n10757), .Z(n10759) );
  AND U11548 ( .A(n10760), .B(n10759), .Z(n10762) );
  XNOR U11549 ( .A(n10762), .B(sreg[1434]), .Z(n10761) );
  XNOR U11550 ( .A(n10763), .B(n10761), .Z(c[1434]) );
  AND U11551 ( .A(b[2]), .B(a[413]), .Z(n10791) );
  AND U11552 ( .A(a[414]), .B(b[1]), .Z(n10789) );
  AND U11553 ( .A(a[412]), .B(b[3]), .Z(n10788) );
  XOR U11554 ( .A(n10789), .B(n10788), .Z(n10790) );
  XOR U11555 ( .A(n10791), .B(n10790), .Z(n10794) );
  NAND U11556 ( .A(b[0]), .B(a[415]), .Z(n10795) );
  XOR U11557 ( .A(n10794), .B(n10795), .Z(n10797) );
  OR U11558 ( .A(n10765), .B(n10764), .Z(n10769) );
  NANDN U11559 ( .A(n10767), .B(n10766), .Z(n10768) );
  NAND U11560 ( .A(n10769), .B(n10768), .Z(n10796) );
  XNOR U11561 ( .A(n10797), .B(n10796), .Z(n10782) );
  NANDN U11562 ( .A(n10771), .B(n10770), .Z(n10775) );
  NAND U11563 ( .A(n10773), .B(n10772), .Z(n10774) );
  NAND U11564 ( .A(n10775), .B(n10774), .Z(n10783) );
  XNOR U11565 ( .A(n10782), .B(n10783), .Z(n10784) );
  NANDN U11566 ( .A(n10777), .B(n10776), .Z(n10781) );
  NANDN U11567 ( .A(n10779), .B(n10778), .Z(n10780) );
  NAND U11568 ( .A(n10781), .B(n10780), .Z(n10785) );
  XOR U11569 ( .A(n10784), .B(n10785), .Z(n10800) );
  XNOR U11570 ( .A(n10800), .B(sreg[1435]), .Z(n10802) );
  XNOR U11571 ( .A(n10801), .B(n10802), .Z(c[1435]) );
  NANDN U11572 ( .A(n10783), .B(n10782), .Z(n10787) );
  NANDN U11573 ( .A(n10785), .B(n10784), .Z(n10786) );
  NAND U11574 ( .A(n10787), .B(n10786), .Z(n10808) );
  AND U11575 ( .A(b[2]), .B(a[414]), .Z(n10814) );
  AND U11576 ( .A(a[415]), .B(b[1]), .Z(n10812) );
  AND U11577 ( .A(a[413]), .B(b[3]), .Z(n10811) );
  XOR U11578 ( .A(n10812), .B(n10811), .Z(n10813) );
  XOR U11579 ( .A(n10814), .B(n10813), .Z(n10817) );
  NAND U11580 ( .A(b[0]), .B(a[416]), .Z(n10818) );
  XOR U11581 ( .A(n10817), .B(n10818), .Z(n10820) );
  OR U11582 ( .A(n10789), .B(n10788), .Z(n10793) );
  NANDN U11583 ( .A(n10791), .B(n10790), .Z(n10792) );
  NAND U11584 ( .A(n10793), .B(n10792), .Z(n10819) );
  XNOR U11585 ( .A(n10820), .B(n10819), .Z(n10805) );
  NANDN U11586 ( .A(n10795), .B(n10794), .Z(n10799) );
  OR U11587 ( .A(n10797), .B(n10796), .Z(n10798) );
  NAND U11588 ( .A(n10799), .B(n10798), .Z(n10806) );
  XNOR U11589 ( .A(n10805), .B(n10806), .Z(n10807) );
  XNOR U11590 ( .A(n10808), .B(n10807), .Z(n10823) );
  XOR U11591 ( .A(sreg[1436]), .B(n10823), .Z(n10824) );
  NAND U11592 ( .A(n10800), .B(sreg[1435]), .Z(n10804) );
  NANDN U11593 ( .A(n10802), .B(n10801), .Z(n10803) );
  NAND U11594 ( .A(n10804), .B(n10803), .Z(n10825) );
  XOR U11595 ( .A(n10824), .B(n10825), .Z(c[1436]) );
  NANDN U11596 ( .A(n10806), .B(n10805), .Z(n10810) );
  NAND U11597 ( .A(n10808), .B(n10807), .Z(n10809) );
  NAND U11598 ( .A(n10810), .B(n10809), .Z(n10834) );
  AND U11599 ( .A(b[2]), .B(a[415]), .Z(n10840) );
  AND U11600 ( .A(a[416]), .B(b[1]), .Z(n10838) );
  AND U11601 ( .A(a[414]), .B(b[3]), .Z(n10837) );
  XOR U11602 ( .A(n10838), .B(n10837), .Z(n10839) );
  XOR U11603 ( .A(n10840), .B(n10839), .Z(n10843) );
  NAND U11604 ( .A(b[0]), .B(a[417]), .Z(n10844) );
  XOR U11605 ( .A(n10843), .B(n10844), .Z(n10846) );
  OR U11606 ( .A(n10812), .B(n10811), .Z(n10816) );
  NANDN U11607 ( .A(n10814), .B(n10813), .Z(n10815) );
  NAND U11608 ( .A(n10816), .B(n10815), .Z(n10845) );
  XNOR U11609 ( .A(n10846), .B(n10845), .Z(n10831) );
  NANDN U11610 ( .A(n10818), .B(n10817), .Z(n10822) );
  OR U11611 ( .A(n10820), .B(n10819), .Z(n10821) );
  NAND U11612 ( .A(n10822), .B(n10821), .Z(n10832) );
  XNOR U11613 ( .A(n10831), .B(n10832), .Z(n10833) );
  XOR U11614 ( .A(n10834), .B(n10833), .Z(n10830) );
  OR U11615 ( .A(n10823), .B(sreg[1436]), .Z(n10827) );
  NANDN U11616 ( .A(n10825), .B(n10824), .Z(n10826) );
  AND U11617 ( .A(n10827), .B(n10826), .Z(n10829) );
  XNOR U11618 ( .A(sreg[1437]), .B(n10829), .Z(n10828) );
  XOR U11619 ( .A(n10830), .B(n10828), .Z(c[1437]) );
  NANDN U11620 ( .A(n10832), .B(n10831), .Z(n10836) );
  NAND U11621 ( .A(n10834), .B(n10833), .Z(n10835) );
  NAND U11622 ( .A(n10836), .B(n10835), .Z(n10852) );
  AND U11623 ( .A(b[2]), .B(a[416]), .Z(n10858) );
  AND U11624 ( .A(a[417]), .B(b[1]), .Z(n10856) );
  AND U11625 ( .A(a[415]), .B(b[3]), .Z(n10855) );
  XOR U11626 ( .A(n10856), .B(n10855), .Z(n10857) );
  XOR U11627 ( .A(n10858), .B(n10857), .Z(n10861) );
  NAND U11628 ( .A(b[0]), .B(a[418]), .Z(n10862) );
  XOR U11629 ( .A(n10861), .B(n10862), .Z(n10864) );
  OR U11630 ( .A(n10838), .B(n10837), .Z(n10842) );
  NANDN U11631 ( .A(n10840), .B(n10839), .Z(n10841) );
  NAND U11632 ( .A(n10842), .B(n10841), .Z(n10863) );
  XNOR U11633 ( .A(n10864), .B(n10863), .Z(n10849) );
  NANDN U11634 ( .A(n10844), .B(n10843), .Z(n10848) );
  OR U11635 ( .A(n10846), .B(n10845), .Z(n10847) );
  NAND U11636 ( .A(n10848), .B(n10847), .Z(n10850) );
  XNOR U11637 ( .A(n10849), .B(n10850), .Z(n10851) );
  XNOR U11638 ( .A(n10852), .B(n10851), .Z(n10867) );
  XNOR U11639 ( .A(n10867), .B(sreg[1438]), .Z(n10868) );
  XOR U11640 ( .A(n10869), .B(n10868), .Z(c[1438]) );
  NANDN U11641 ( .A(n10850), .B(n10849), .Z(n10854) );
  NAND U11642 ( .A(n10852), .B(n10851), .Z(n10853) );
  NAND U11643 ( .A(n10854), .B(n10853), .Z(n10878) );
  AND U11644 ( .A(b[2]), .B(a[417]), .Z(n10884) );
  AND U11645 ( .A(a[418]), .B(b[1]), .Z(n10882) );
  AND U11646 ( .A(a[416]), .B(b[3]), .Z(n10881) );
  XOR U11647 ( .A(n10882), .B(n10881), .Z(n10883) );
  XOR U11648 ( .A(n10884), .B(n10883), .Z(n10887) );
  NAND U11649 ( .A(b[0]), .B(a[419]), .Z(n10888) );
  XOR U11650 ( .A(n10887), .B(n10888), .Z(n10890) );
  OR U11651 ( .A(n10856), .B(n10855), .Z(n10860) );
  NANDN U11652 ( .A(n10858), .B(n10857), .Z(n10859) );
  NAND U11653 ( .A(n10860), .B(n10859), .Z(n10889) );
  XNOR U11654 ( .A(n10890), .B(n10889), .Z(n10875) );
  NANDN U11655 ( .A(n10862), .B(n10861), .Z(n10866) );
  OR U11656 ( .A(n10864), .B(n10863), .Z(n10865) );
  NAND U11657 ( .A(n10866), .B(n10865), .Z(n10876) );
  XNOR U11658 ( .A(n10875), .B(n10876), .Z(n10877) );
  XOR U11659 ( .A(n10878), .B(n10877), .Z(n10874) );
  NAND U11660 ( .A(n10867), .B(sreg[1438]), .Z(n10871) );
  OR U11661 ( .A(n10869), .B(n10868), .Z(n10870) );
  NAND U11662 ( .A(n10871), .B(n10870), .Z(n10873) );
  XNOR U11663 ( .A(sreg[1439]), .B(n10873), .Z(n10872) );
  XOR U11664 ( .A(n10874), .B(n10872), .Z(c[1439]) );
  NANDN U11665 ( .A(n10876), .B(n10875), .Z(n10880) );
  NAND U11666 ( .A(n10878), .B(n10877), .Z(n10879) );
  NAND U11667 ( .A(n10880), .B(n10879), .Z(n10896) );
  AND U11668 ( .A(b[2]), .B(a[418]), .Z(n10902) );
  AND U11669 ( .A(a[419]), .B(b[1]), .Z(n10900) );
  AND U11670 ( .A(a[417]), .B(b[3]), .Z(n10899) );
  XOR U11671 ( .A(n10900), .B(n10899), .Z(n10901) );
  XOR U11672 ( .A(n10902), .B(n10901), .Z(n10905) );
  NAND U11673 ( .A(b[0]), .B(a[420]), .Z(n10906) );
  XOR U11674 ( .A(n10905), .B(n10906), .Z(n10908) );
  OR U11675 ( .A(n10882), .B(n10881), .Z(n10886) );
  NANDN U11676 ( .A(n10884), .B(n10883), .Z(n10885) );
  NAND U11677 ( .A(n10886), .B(n10885), .Z(n10907) );
  XNOR U11678 ( .A(n10908), .B(n10907), .Z(n10893) );
  NANDN U11679 ( .A(n10888), .B(n10887), .Z(n10892) );
  OR U11680 ( .A(n10890), .B(n10889), .Z(n10891) );
  NAND U11681 ( .A(n10892), .B(n10891), .Z(n10894) );
  XNOR U11682 ( .A(n10893), .B(n10894), .Z(n10895) );
  XNOR U11683 ( .A(n10896), .B(n10895), .Z(n10911) );
  XNOR U11684 ( .A(n10911), .B(sreg[1440]), .Z(n10912) );
  XOR U11685 ( .A(n10913), .B(n10912), .Z(c[1440]) );
  NANDN U11686 ( .A(n10894), .B(n10893), .Z(n10898) );
  NAND U11687 ( .A(n10896), .B(n10895), .Z(n10897) );
  NAND U11688 ( .A(n10898), .B(n10897), .Z(n10919) );
  AND U11689 ( .A(b[2]), .B(a[419]), .Z(n10925) );
  AND U11690 ( .A(a[420]), .B(b[1]), .Z(n10923) );
  AND U11691 ( .A(a[418]), .B(b[3]), .Z(n10922) );
  XOR U11692 ( .A(n10923), .B(n10922), .Z(n10924) );
  XOR U11693 ( .A(n10925), .B(n10924), .Z(n10928) );
  NAND U11694 ( .A(b[0]), .B(a[421]), .Z(n10929) );
  XOR U11695 ( .A(n10928), .B(n10929), .Z(n10931) );
  OR U11696 ( .A(n10900), .B(n10899), .Z(n10904) );
  NANDN U11697 ( .A(n10902), .B(n10901), .Z(n10903) );
  NAND U11698 ( .A(n10904), .B(n10903), .Z(n10930) );
  XNOR U11699 ( .A(n10931), .B(n10930), .Z(n10916) );
  NANDN U11700 ( .A(n10906), .B(n10905), .Z(n10910) );
  OR U11701 ( .A(n10908), .B(n10907), .Z(n10909) );
  NAND U11702 ( .A(n10910), .B(n10909), .Z(n10917) );
  XNOR U11703 ( .A(n10916), .B(n10917), .Z(n10918) );
  XNOR U11704 ( .A(n10919), .B(n10918), .Z(n10934) );
  XOR U11705 ( .A(sreg[1441]), .B(n10934), .Z(n10935) );
  NAND U11706 ( .A(n10911), .B(sreg[1440]), .Z(n10915) );
  OR U11707 ( .A(n10913), .B(n10912), .Z(n10914) );
  NAND U11708 ( .A(n10915), .B(n10914), .Z(n10936) );
  XOR U11709 ( .A(n10935), .B(n10936), .Z(c[1441]) );
  NANDN U11710 ( .A(n10917), .B(n10916), .Z(n10921) );
  NAND U11711 ( .A(n10919), .B(n10918), .Z(n10920) );
  NAND U11712 ( .A(n10921), .B(n10920), .Z(n10945) );
  AND U11713 ( .A(b[2]), .B(a[420]), .Z(n10951) );
  AND U11714 ( .A(a[421]), .B(b[1]), .Z(n10949) );
  AND U11715 ( .A(a[419]), .B(b[3]), .Z(n10948) );
  XOR U11716 ( .A(n10949), .B(n10948), .Z(n10950) );
  XOR U11717 ( .A(n10951), .B(n10950), .Z(n10954) );
  NAND U11718 ( .A(b[0]), .B(a[422]), .Z(n10955) );
  XOR U11719 ( .A(n10954), .B(n10955), .Z(n10957) );
  OR U11720 ( .A(n10923), .B(n10922), .Z(n10927) );
  NANDN U11721 ( .A(n10925), .B(n10924), .Z(n10926) );
  NAND U11722 ( .A(n10927), .B(n10926), .Z(n10956) );
  XNOR U11723 ( .A(n10957), .B(n10956), .Z(n10942) );
  NANDN U11724 ( .A(n10929), .B(n10928), .Z(n10933) );
  OR U11725 ( .A(n10931), .B(n10930), .Z(n10932) );
  NAND U11726 ( .A(n10933), .B(n10932), .Z(n10943) );
  XNOR U11727 ( .A(n10942), .B(n10943), .Z(n10944) );
  XOR U11728 ( .A(n10945), .B(n10944), .Z(n10941) );
  OR U11729 ( .A(n10934), .B(sreg[1441]), .Z(n10938) );
  NANDN U11730 ( .A(n10936), .B(n10935), .Z(n10937) );
  AND U11731 ( .A(n10938), .B(n10937), .Z(n10940) );
  XNOR U11732 ( .A(sreg[1442]), .B(n10940), .Z(n10939) );
  XOR U11733 ( .A(n10941), .B(n10939), .Z(c[1442]) );
  NANDN U11734 ( .A(n10943), .B(n10942), .Z(n10947) );
  NAND U11735 ( .A(n10945), .B(n10944), .Z(n10946) );
  NAND U11736 ( .A(n10947), .B(n10946), .Z(n10963) );
  AND U11737 ( .A(b[2]), .B(a[421]), .Z(n10969) );
  AND U11738 ( .A(a[422]), .B(b[1]), .Z(n10967) );
  AND U11739 ( .A(a[420]), .B(b[3]), .Z(n10966) );
  XOR U11740 ( .A(n10967), .B(n10966), .Z(n10968) );
  XOR U11741 ( .A(n10969), .B(n10968), .Z(n10972) );
  NAND U11742 ( .A(b[0]), .B(a[423]), .Z(n10973) );
  XOR U11743 ( .A(n10972), .B(n10973), .Z(n10975) );
  OR U11744 ( .A(n10949), .B(n10948), .Z(n10953) );
  NANDN U11745 ( .A(n10951), .B(n10950), .Z(n10952) );
  NAND U11746 ( .A(n10953), .B(n10952), .Z(n10974) );
  XNOR U11747 ( .A(n10975), .B(n10974), .Z(n10960) );
  NANDN U11748 ( .A(n10955), .B(n10954), .Z(n10959) );
  OR U11749 ( .A(n10957), .B(n10956), .Z(n10958) );
  NAND U11750 ( .A(n10959), .B(n10958), .Z(n10961) );
  XNOR U11751 ( .A(n10960), .B(n10961), .Z(n10962) );
  XNOR U11752 ( .A(n10963), .B(n10962), .Z(n10978) );
  XNOR U11753 ( .A(n10978), .B(sreg[1443]), .Z(n10979) );
  XOR U11754 ( .A(n10980), .B(n10979), .Z(c[1443]) );
  NANDN U11755 ( .A(n10961), .B(n10960), .Z(n10965) );
  NAND U11756 ( .A(n10963), .B(n10962), .Z(n10964) );
  NAND U11757 ( .A(n10965), .B(n10964), .Z(n10986) );
  AND U11758 ( .A(b[2]), .B(a[422]), .Z(n10998) );
  AND U11759 ( .A(a[423]), .B(b[1]), .Z(n10996) );
  AND U11760 ( .A(a[421]), .B(b[3]), .Z(n10995) );
  XOR U11761 ( .A(n10996), .B(n10995), .Z(n10997) );
  XOR U11762 ( .A(n10998), .B(n10997), .Z(n10989) );
  NAND U11763 ( .A(b[0]), .B(a[424]), .Z(n10990) );
  XOR U11764 ( .A(n10989), .B(n10990), .Z(n10992) );
  OR U11765 ( .A(n10967), .B(n10966), .Z(n10971) );
  NANDN U11766 ( .A(n10969), .B(n10968), .Z(n10970) );
  NAND U11767 ( .A(n10971), .B(n10970), .Z(n10991) );
  XNOR U11768 ( .A(n10992), .B(n10991), .Z(n10983) );
  NANDN U11769 ( .A(n10973), .B(n10972), .Z(n10977) );
  OR U11770 ( .A(n10975), .B(n10974), .Z(n10976) );
  NAND U11771 ( .A(n10977), .B(n10976), .Z(n10984) );
  XNOR U11772 ( .A(n10983), .B(n10984), .Z(n10985) );
  XNOR U11773 ( .A(n10986), .B(n10985), .Z(n11001) );
  XOR U11774 ( .A(sreg[1444]), .B(n11001), .Z(n11002) );
  NAND U11775 ( .A(n10978), .B(sreg[1443]), .Z(n10982) );
  OR U11776 ( .A(n10980), .B(n10979), .Z(n10981) );
  NAND U11777 ( .A(n10982), .B(n10981), .Z(n11003) );
  XOR U11778 ( .A(n11002), .B(n11003), .Z(c[1444]) );
  NANDN U11779 ( .A(n10984), .B(n10983), .Z(n10988) );
  NAND U11780 ( .A(n10986), .B(n10985), .Z(n10987) );
  NAND U11781 ( .A(n10988), .B(n10987), .Z(n11012) );
  NANDN U11782 ( .A(n10990), .B(n10989), .Z(n10994) );
  OR U11783 ( .A(n10992), .B(n10991), .Z(n10993) );
  NAND U11784 ( .A(n10994), .B(n10993), .Z(n11009) );
  AND U11785 ( .A(b[2]), .B(a[423]), .Z(n11018) );
  AND U11786 ( .A(a[424]), .B(b[1]), .Z(n11016) );
  AND U11787 ( .A(a[422]), .B(b[3]), .Z(n11015) );
  XOR U11788 ( .A(n11016), .B(n11015), .Z(n11017) );
  XOR U11789 ( .A(n11018), .B(n11017), .Z(n11021) );
  NAND U11790 ( .A(b[0]), .B(a[425]), .Z(n11022) );
  XNOR U11791 ( .A(n11021), .B(n11022), .Z(n11023) );
  OR U11792 ( .A(n10996), .B(n10995), .Z(n11000) );
  NANDN U11793 ( .A(n10998), .B(n10997), .Z(n10999) );
  AND U11794 ( .A(n11000), .B(n10999), .Z(n11024) );
  XNOR U11795 ( .A(n11023), .B(n11024), .Z(n11010) );
  XNOR U11796 ( .A(n11009), .B(n11010), .Z(n11011) );
  XNOR U11797 ( .A(n11012), .B(n11011), .Z(n11008) );
  OR U11798 ( .A(n11001), .B(sreg[1444]), .Z(n11005) );
  NANDN U11799 ( .A(n11003), .B(n11002), .Z(n11004) );
  AND U11800 ( .A(n11005), .B(n11004), .Z(n11007) );
  XNOR U11801 ( .A(sreg[1445]), .B(n11007), .Z(n11006) );
  XNOR U11802 ( .A(n11008), .B(n11006), .Z(c[1445]) );
  NANDN U11803 ( .A(n11010), .B(n11009), .Z(n11014) );
  NANDN U11804 ( .A(n11012), .B(n11011), .Z(n11013) );
  NAND U11805 ( .A(n11014), .B(n11013), .Z(n11042) );
  AND U11806 ( .A(b[2]), .B(a[424]), .Z(n11036) );
  AND U11807 ( .A(a[425]), .B(b[1]), .Z(n11034) );
  AND U11808 ( .A(a[423]), .B(b[3]), .Z(n11033) );
  XOR U11809 ( .A(n11034), .B(n11033), .Z(n11035) );
  XOR U11810 ( .A(n11036), .B(n11035), .Z(n11027) );
  NAND U11811 ( .A(b[0]), .B(a[426]), .Z(n11028) );
  XOR U11812 ( .A(n11027), .B(n11028), .Z(n11030) );
  OR U11813 ( .A(n11016), .B(n11015), .Z(n11020) );
  NANDN U11814 ( .A(n11018), .B(n11017), .Z(n11019) );
  NAND U11815 ( .A(n11020), .B(n11019), .Z(n11029) );
  XNOR U11816 ( .A(n11030), .B(n11029), .Z(n11039) );
  NANDN U11817 ( .A(n11022), .B(n11021), .Z(n11026) );
  NAND U11818 ( .A(n11024), .B(n11023), .Z(n11025) );
  NAND U11819 ( .A(n11026), .B(n11025), .Z(n11040) );
  XNOR U11820 ( .A(n11039), .B(n11040), .Z(n11041) );
  XOR U11821 ( .A(n11042), .B(n11041), .Z(n11045) );
  XNOR U11822 ( .A(n11045), .B(sreg[1446]), .Z(n11046) );
  XOR U11823 ( .A(n11047), .B(n11046), .Z(c[1446]) );
  NANDN U11824 ( .A(n11028), .B(n11027), .Z(n11032) );
  OR U11825 ( .A(n11030), .B(n11029), .Z(n11031) );
  NAND U11826 ( .A(n11032), .B(n11031), .Z(n11050) );
  AND U11827 ( .A(b[2]), .B(a[425]), .Z(n11065) );
  AND U11828 ( .A(a[426]), .B(b[1]), .Z(n11063) );
  AND U11829 ( .A(a[424]), .B(b[3]), .Z(n11062) );
  XOR U11830 ( .A(n11063), .B(n11062), .Z(n11064) );
  XOR U11831 ( .A(n11065), .B(n11064), .Z(n11056) );
  NAND U11832 ( .A(b[0]), .B(a[427]), .Z(n11057) );
  XNOR U11833 ( .A(n11056), .B(n11057), .Z(n11058) );
  OR U11834 ( .A(n11034), .B(n11033), .Z(n11038) );
  NANDN U11835 ( .A(n11036), .B(n11035), .Z(n11037) );
  AND U11836 ( .A(n11038), .B(n11037), .Z(n11059) );
  XNOR U11837 ( .A(n11058), .B(n11059), .Z(n11051) );
  XNOR U11838 ( .A(n11050), .B(n11051), .Z(n11052) );
  NANDN U11839 ( .A(n11040), .B(n11039), .Z(n11044) );
  NANDN U11840 ( .A(n11042), .B(n11041), .Z(n11043) );
  NAND U11841 ( .A(n11044), .B(n11043), .Z(n11053) );
  XNOR U11842 ( .A(n11052), .B(n11053), .Z(n11068) );
  XOR U11843 ( .A(sreg[1447]), .B(n11068), .Z(n11069) );
  NAND U11844 ( .A(n11045), .B(sreg[1446]), .Z(n11049) );
  OR U11845 ( .A(n11047), .B(n11046), .Z(n11048) );
  NAND U11846 ( .A(n11049), .B(n11048), .Z(n11070) );
  XOR U11847 ( .A(n11069), .B(n11070), .Z(c[1447]) );
  NANDN U11848 ( .A(n11051), .B(n11050), .Z(n11055) );
  NANDN U11849 ( .A(n11053), .B(n11052), .Z(n11054) );
  NAND U11850 ( .A(n11055), .B(n11054), .Z(n11079) );
  NANDN U11851 ( .A(n11057), .B(n11056), .Z(n11061) );
  NAND U11852 ( .A(n11059), .B(n11058), .Z(n11060) );
  NAND U11853 ( .A(n11061), .B(n11060), .Z(n11076) );
  AND U11854 ( .A(b[2]), .B(a[426]), .Z(n11085) );
  AND U11855 ( .A(a[427]), .B(b[1]), .Z(n11083) );
  AND U11856 ( .A(a[425]), .B(b[3]), .Z(n11082) );
  XOR U11857 ( .A(n11083), .B(n11082), .Z(n11084) );
  XOR U11858 ( .A(n11085), .B(n11084), .Z(n11088) );
  NAND U11859 ( .A(b[0]), .B(a[428]), .Z(n11089) );
  XNOR U11860 ( .A(n11088), .B(n11089), .Z(n11090) );
  OR U11861 ( .A(n11063), .B(n11062), .Z(n11067) );
  NANDN U11862 ( .A(n11065), .B(n11064), .Z(n11066) );
  AND U11863 ( .A(n11067), .B(n11066), .Z(n11091) );
  XNOR U11864 ( .A(n11090), .B(n11091), .Z(n11077) );
  XNOR U11865 ( .A(n11076), .B(n11077), .Z(n11078) );
  XOR U11866 ( .A(n11079), .B(n11078), .Z(n11075) );
  OR U11867 ( .A(n11068), .B(sreg[1447]), .Z(n11072) );
  NANDN U11868 ( .A(n11070), .B(n11069), .Z(n11071) );
  AND U11869 ( .A(n11072), .B(n11071), .Z(n11074) );
  XOR U11870 ( .A(sreg[1448]), .B(n11074), .Z(n11073) );
  XOR U11871 ( .A(n11075), .B(n11073), .Z(c[1448]) );
  NANDN U11872 ( .A(n11077), .B(n11076), .Z(n11081) );
  NAND U11873 ( .A(n11079), .B(n11078), .Z(n11080) );
  NAND U11874 ( .A(n11081), .B(n11080), .Z(n11097) );
  AND U11875 ( .A(b[2]), .B(a[427]), .Z(n11103) );
  AND U11876 ( .A(a[428]), .B(b[1]), .Z(n11101) );
  AND U11877 ( .A(a[426]), .B(b[3]), .Z(n11100) );
  XOR U11878 ( .A(n11101), .B(n11100), .Z(n11102) );
  XOR U11879 ( .A(n11103), .B(n11102), .Z(n11106) );
  NAND U11880 ( .A(b[0]), .B(a[429]), .Z(n11107) );
  XOR U11881 ( .A(n11106), .B(n11107), .Z(n11109) );
  OR U11882 ( .A(n11083), .B(n11082), .Z(n11087) );
  NANDN U11883 ( .A(n11085), .B(n11084), .Z(n11086) );
  NAND U11884 ( .A(n11087), .B(n11086), .Z(n11108) );
  XNOR U11885 ( .A(n11109), .B(n11108), .Z(n11094) );
  NANDN U11886 ( .A(n11089), .B(n11088), .Z(n11093) );
  NAND U11887 ( .A(n11091), .B(n11090), .Z(n11092) );
  NAND U11888 ( .A(n11093), .B(n11092), .Z(n11095) );
  XNOR U11889 ( .A(n11094), .B(n11095), .Z(n11096) );
  XOR U11890 ( .A(n11097), .B(n11096), .Z(n11112) );
  XNOR U11891 ( .A(n11112), .B(sreg[1449]), .Z(n11114) );
  XNOR U11892 ( .A(n11113), .B(n11114), .Z(c[1449]) );
  NANDN U11893 ( .A(n11095), .B(n11094), .Z(n11099) );
  NANDN U11894 ( .A(n11097), .B(n11096), .Z(n11098) );
  NAND U11895 ( .A(n11099), .B(n11098), .Z(n11123) );
  AND U11896 ( .A(b[2]), .B(a[428]), .Z(n11129) );
  AND U11897 ( .A(a[429]), .B(b[1]), .Z(n11127) );
  AND U11898 ( .A(a[427]), .B(b[3]), .Z(n11126) );
  XOR U11899 ( .A(n11127), .B(n11126), .Z(n11128) );
  XOR U11900 ( .A(n11129), .B(n11128), .Z(n11132) );
  NAND U11901 ( .A(b[0]), .B(a[430]), .Z(n11133) );
  XOR U11902 ( .A(n11132), .B(n11133), .Z(n11135) );
  OR U11903 ( .A(n11101), .B(n11100), .Z(n11105) );
  NANDN U11904 ( .A(n11103), .B(n11102), .Z(n11104) );
  NAND U11905 ( .A(n11105), .B(n11104), .Z(n11134) );
  XNOR U11906 ( .A(n11135), .B(n11134), .Z(n11120) );
  NANDN U11907 ( .A(n11107), .B(n11106), .Z(n11111) );
  OR U11908 ( .A(n11109), .B(n11108), .Z(n11110) );
  NAND U11909 ( .A(n11111), .B(n11110), .Z(n11121) );
  XNOR U11910 ( .A(n11120), .B(n11121), .Z(n11122) );
  XOR U11911 ( .A(n11123), .B(n11122), .Z(n11119) );
  NAND U11912 ( .A(n11112), .B(sreg[1449]), .Z(n11116) );
  NANDN U11913 ( .A(n11114), .B(n11113), .Z(n11115) );
  NAND U11914 ( .A(n11116), .B(n11115), .Z(n11118) );
  XNOR U11915 ( .A(sreg[1450]), .B(n11118), .Z(n11117) );
  XOR U11916 ( .A(n11119), .B(n11117), .Z(c[1450]) );
  NANDN U11917 ( .A(n11121), .B(n11120), .Z(n11125) );
  NAND U11918 ( .A(n11123), .B(n11122), .Z(n11124) );
  NAND U11919 ( .A(n11125), .B(n11124), .Z(n11141) );
  AND U11920 ( .A(b[2]), .B(a[429]), .Z(n11147) );
  AND U11921 ( .A(a[430]), .B(b[1]), .Z(n11145) );
  AND U11922 ( .A(a[428]), .B(b[3]), .Z(n11144) );
  XOR U11923 ( .A(n11145), .B(n11144), .Z(n11146) );
  XOR U11924 ( .A(n11147), .B(n11146), .Z(n11150) );
  NAND U11925 ( .A(b[0]), .B(a[431]), .Z(n11151) );
  XOR U11926 ( .A(n11150), .B(n11151), .Z(n11153) );
  OR U11927 ( .A(n11127), .B(n11126), .Z(n11131) );
  NANDN U11928 ( .A(n11129), .B(n11128), .Z(n11130) );
  NAND U11929 ( .A(n11131), .B(n11130), .Z(n11152) );
  XNOR U11930 ( .A(n11153), .B(n11152), .Z(n11138) );
  NANDN U11931 ( .A(n11133), .B(n11132), .Z(n11137) );
  OR U11932 ( .A(n11135), .B(n11134), .Z(n11136) );
  NAND U11933 ( .A(n11137), .B(n11136), .Z(n11139) );
  XNOR U11934 ( .A(n11138), .B(n11139), .Z(n11140) );
  XNOR U11935 ( .A(n11141), .B(n11140), .Z(n11156) );
  XNOR U11936 ( .A(n11156), .B(sreg[1451]), .Z(n11157) );
  XOR U11937 ( .A(n11158), .B(n11157), .Z(c[1451]) );
  NANDN U11938 ( .A(n11139), .B(n11138), .Z(n11143) );
  NAND U11939 ( .A(n11141), .B(n11140), .Z(n11142) );
  NAND U11940 ( .A(n11143), .B(n11142), .Z(n11164) );
  AND U11941 ( .A(b[2]), .B(a[430]), .Z(n11170) );
  AND U11942 ( .A(a[431]), .B(b[1]), .Z(n11168) );
  AND U11943 ( .A(a[429]), .B(b[3]), .Z(n11167) );
  XOR U11944 ( .A(n11168), .B(n11167), .Z(n11169) );
  XOR U11945 ( .A(n11170), .B(n11169), .Z(n11173) );
  NAND U11946 ( .A(b[0]), .B(a[432]), .Z(n11174) );
  XOR U11947 ( .A(n11173), .B(n11174), .Z(n11176) );
  OR U11948 ( .A(n11145), .B(n11144), .Z(n11149) );
  NANDN U11949 ( .A(n11147), .B(n11146), .Z(n11148) );
  NAND U11950 ( .A(n11149), .B(n11148), .Z(n11175) );
  XNOR U11951 ( .A(n11176), .B(n11175), .Z(n11161) );
  NANDN U11952 ( .A(n11151), .B(n11150), .Z(n11155) );
  OR U11953 ( .A(n11153), .B(n11152), .Z(n11154) );
  NAND U11954 ( .A(n11155), .B(n11154), .Z(n11162) );
  XNOR U11955 ( .A(n11161), .B(n11162), .Z(n11163) );
  XNOR U11956 ( .A(n11164), .B(n11163), .Z(n11179) );
  XOR U11957 ( .A(sreg[1452]), .B(n11179), .Z(n11180) );
  NAND U11958 ( .A(n11156), .B(sreg[1451]), .Z(n11160) );
  OR U11959 ( .A(n11158), .B(n11157), .Z(n11159) );
  NAND U11960 ( .A(n11160), .B(n11159), .Z(n11181) );
  XOR U11961 ( .A(n11180), .B(n11181), .Z(c[1452]) );
  NANDN U11962 ( .A(n11162), .B(n11161), .Z(n11166) );
  NAND U11963 ( .A(n11164), .B(n11163), .Z(n11165) );
  NAND U11964 ( .A(n11166), .B(n11165), .Z(n11190) );
  AND U11965 ( .A(b[2]), .B(a[431]), .Z(n11196) );
  AND U11966 ( .A(a[432]), .B(b[1]), .Z(n11194) );
  AND U11967 ( .A(a[430]), .B(b[3]), .Z(n11193) );
  XOR U11968 ( .A(n11194), .B(n11193), .Z(n11195) );
  XOR U11969 ( .A(n11196), .B(n11195), .Z(n11199) );
  NAND U11970 ( .A(b[0]), .B(a[433]), .Z(n11200) );
  XOR U11971 ( .A(n11199), .B(n11200), .Z(n11202) );
  OR U11972 ( .A(n11168), .B(n11167), .Z(n11172) );
  NANDN U11973 ( .A(n11170), .B(n11169), .Z(n11171) );
  NAND U11974 ( .A(n11172), .B(n11171), .Z(n11201) );
  XNOR U11975 ( .A(n11202), .B(n11201), .Z(n11187) );
  NANDN U11976 ( .A(n11174), .B(n11173), .Z(n11178) );
  OR U11977 ( .A(n11176), .B(n11175), .Z(n11177) );
  NAND U11978 ( .A(n11178), .B(n11177), .Z(n11188) );
  XNOR U11979 ( .A(n11187), .B(n11188), .Z(n11189) );
  XOR U11980 ( .A(n11190), .B(n11189), .Z(n11186) );
  OR U11981 ( .A(n11179), .B(sreg[1452]), .Z(n11183) );
  NANDN U11982 ( .A(n11181), .B(n11180), .Z(n11182) );
  AND U11983 ( .A(n11183), .B(n11182), .Z(n11185) );
  XNOR U11984 ( .A(sreg[1453]), .B(n11185), .Z(n11184) );
  XOR U11985 ( .A(n11186), .B(n11184), .Z(c[1453]) );
  NANDN U11986 ( .A(n11188), .B(n11187), .Z(n11192) );
  NAND U11987 ( .A(n11190), .B(n11189), .Z(n11191) );
  NAND U11988 ( .A(n11192), .B(n11191), .Z(n11208) );
  AND U11989 ( .A(b[2]), .B(a[432]), .Z(n11214) );
  AND U11990 ( .A(a[433]), .B(b[1]), .Z(n11212) );
  AND U11991 ( .A(a[431]), .B(b[3]), .Z(n11211) );
  XOR U11992 ( .A(n11212), .B(n11211), .Z(n11213) );
  XOR U11993 ( .A(n11214), .B(n11213), .Z(n11217) );
  NAND U11994 ( .A(b[0]), .B(a[434]), .Z(n11218) );
  XOR U11995 ( .A(n11217), .B(n11218), .Z(n11220) );
  OR U11996 ( .A(n11194), .B(n11193), .Z(n11198) );
  NANDN U11997 ( .A(n11196), .B(n11195), .Z(n11197) );
  NAND U11998 ( .A(n11198), .B(n11197), .Z(n11219) );
  XNOR U11999 ( .A(n11220), .B(n11219), .Z(n11205) );
  NANDN U12000 ( .A(n11200), .B(n11199), .Z(n11204) );
  OR U12001 ( .A(n11202), .B(n11201), .Z(n11203) );
  NAND U12002 ( .A(n11204), .B(n11203), .Z(n11206) );
  XNOR U12003 ( .A(n11205), .B(n11206), .Z(n11207) );
  XNOR U12004 ( .A(n11208), .B(n11207), .Z(n11223) );
  XNOR U12005 ( .A(n11223), .B(sreg[1454]), .Z(n11224) );
  XOR U12006 ( .A(n11225), .B(n11224), .Z(c[1454]) );
  NANDN U12007 ( .A(n11206), .B(n11205), .Z(n11210) );
  NAND U12008 ( .A(n11208), .B(n11207), .Z(n11209) );
  NAND U12009 ( .A(n11210), .B(n11209), .Z(n11234) );
  AND U12010 ( .A(b[2]), .B(a[433]), .Z(n11240) );
  AND U12011 ( .A(a[434]), .B(b[1]), .Z(n11238) );
  AND U12012 ( .A(a[432]), .B(b[3]), .Z(n11237) );
  XOR U12013 ( .A(n11238), .B(n11237), .Z(n11239) );
  XOR U12014 ( .A(n11240), .B(n11239), .Z(n11243) );
  NAND U12015 ( .A(b[0]), .B(a[435]), .Z(n11244) );
  XOR U12016 ( .A(n11243), .B(n11244), .Z(n11246) );
  OR U12017 ( .A(n11212), .B(n11211), .Z(n11216) );
  NANDN U12018 ( .A(n11214), .B(n11213), .Z(n11215) );
  NAND U12019 ( .A(n11216), .B(n11215), .Z(n11245) );
  XNOR U12020 ( .A(n11246), .B(n11245), .Z(n11231) );
  NANDN U12021 ( .A(n11218), .B(n11217), .Z(n11222) );
  OR U12022 ( .A(n11220), .B(n11219), .Z(n11221) );
  NAND U12023 ( .A(n11222), .B(n11221), .Z(n11232) );
  XNOR U12024 ( .A(n11231), .B(n11232), .Z(n11233) );
  XOR U12025 ( .A(n11234), .B(n11233), .Z(n11230) );
  NAND U12026 ( .A(n11223), .B(sreg[1454]), .Z(n11227) );
  OR U12027 ( .A(n11225), .B(n11224), .Z(n11226) );
  NAND U12028 ( .A(n11227), .B(n11226), .Z(n11229) );
  XNOR U12029 ( .A(sreg[1455]), .B(n11229), .Z(n11228) );
  XOR U12030 ( .A(n11230), .B(n11228), .Z(c[1455]) );
  NANDN U12031 ( .A(n11232), .B(n11231), .Z(n11236) );
  NAND U12032 ( .A(n11234), .B(n11233), .Z(n11235) );
  NAND U12033 ( .A(n11236), .B(n11235), .Z(n11252) );
  AND U12034 ( .A(b[2]), .B(a[434]), .Z(n11258) );
  AND U12035 ( .A(a[435]), .B(b[1]), .Z(n11256) );
  AND U12036 ( .A(a[433]), .B(b[3]), .Z(n11255) );
  XOR U12037 ( .A(n11256), .B(n11255), .Z(n11257) );
  XOR U12038 ( .A(n11258), .B(n11257), .Z(n11261) );
  NAND U12039 ( .A(b[0]), .B(a[436]), .Z(n11262) );
  XOR U12040 ( .A(n11261), .B(n11262), .Z(n11264) );
  OR U12041 ( .A(n11238), .B(n11237), .Z(n11242) );
  NANDN U12042 ( .A(n11240), .B(n11239), .Z(n11241) );
  NAND U12043 ( .A(n11242), .B(n11241), .Z(n11263) );
  XNOR U12044 ( .A(n11264), .B(n11263), .Z(n11249) );
  NANDN U12045 ( .A(n11244), .B(n11243), .Z(n11248) );
  OR U12046 ( .A(n11246), .B(n11245), .Z(n11247) );
  NAND U12047 ( .A(n11248), .B(n11247), .Z(n11250) );
  XNOR U12048 ( .A(n11249), .B(n11250), .Z(n11251) );
  XNOR U12049 ( .A(n11252), .B(n11251), .Z(n11267) );
  XNOR U12050 ( .A(n11267), .B(sreg[1456]), .Z(n11268) );
  XOR U12051 ( .A(n11269), .B(n11268), .Z(c[1456]) );
  NANDN U12052 ( .A(n11250), .B(n11249), .Z(n11254) );
  NAND U12053 ( .A(n11252), .B(n11251), .Z(n11253) );
  NAND U12054 ( .A(n11254), .B(n11253), .Z(n11280) );
  AND U12055 ( .A(b[2]), .B(a[435]), .Z(n11286) );
  AND U12056 ( .A(a[436]), .B(b[1]), .Z(n11284) );
  AND U12057 ( .A(a[434]), .B(b[3]), .Z(n11283) );
  XOR U12058 ( .A(n11284), .B(n11283), .Z(n11285) );
  XOR U12059 ( .A(n11286), .B(n11285), .Z(n11289) );
  NAND U12060 ( .A(b[0]), .B(a[437]), .Z(n11290) );
  XOR U12061 ( .A(n11289), .B(n11290), .Z(n11292) );
  OR U12062 ( .A(n11256), .B(n11255), .Z(n11260) );
  NANDN U12063 ( .A(n11258), .B(n11257), .Z(n11259) );
  NAND U12064 ( .A(n11260), .B(n11259), .Z(n11291) );
  XNOR U12065 ( .A(n11292), .B(n11291), .Z(n11277) );
  NANDN U12066 ( .A(n11262), .B(n11261), .Z(n11266) );
  OR U12067 ( .A(n11264), .B(n11263), .Z(n11265) );
  NAND U12068 ( .A(n11266), .B(n11265), .Z(n11278) );
  XNOR U12069 ( .A(n11277), .B(n11278), .Z(n11279) );
  XNOR U12070 ( .A(n11280), .B(n11279), .Z(n11272) );
  XOR U12071 ( .A(sreg[1457]), .B(n11272), .Z(n11273) );
  NAND U12072 ( .A(n11267), .B(sreg[1456]), .Z(n11271) );
  OR U12073 ( .A(n11269), .B(n11268), .Z(n11270) );
  NAND U12074 ( .A(n11271), .B(n11270), .Z(n11274) );
  XOR U12075 ( .A(n11273), .B(n11274), .Z(c[1457]) );
  OR U12076 ( .A(n11272), .B(sreg[1457]), .Z(n11276) );
  NANDN U12077 ( .A(n11274), .B(n11273), .Z(n11275) );
  AND U12078 ( .A(n11276), .B(n11275), .Z(n11315) );
  NANDN U12079 ( .A(n11278), .B(n11277), .Z(n11282) );
  NAND U12080 ( .A(n11280), .B(n11279), .Z(n11281) );
  NAND U12081 ( .A(n11282), .B(n11281), .Z(n11299) );
  AND U12082 ( .A(b[2]), .B(a[436]), .Z(n11305) );
  AND U12083 ( .A(a[437]), .B(b[1]), .Z(n11303) );
  AND U12084 ( .A(a[435]), .B(b[3]), .Z(n11302) );
  XOR U12085 ( .A(n11303), .B(n11302), .Z(n11304) );
  XOR U12086 ( .A(n11305), .B(n11304), .Z(n11308) );
  NAND U12087 ( .A(b[0]), .B(a[438]), .Z(n11309) );
  XOR U12088 ( .A(n11308), .B(n11309), .Z(n11311) );
  OR U12089 ( .A(n11284), .B(n11283), .Z(n11288) );
  NANDN U12090 ( .A(n11286), .B(n11285), .Z(n11287) );
  NAND U12091 ( .A(n11288), .B(n11287), .Z(n11310) );
  XNOR U12092 ( .A(n11311), .B(n11310), .Z(n11296) );
  NANDN U12093 ( .A(n11290), .B(n11289), .Z(n11294) );
  OR U12094 ( .A(n11292), .B(n11291), .Z(n11293) );
  NAND U12095 ( .A(n11294), .B(n11293), .Z(n11297) );
  XNOR U12096 ( .A(n11296), .B(n11297), .Z(n11298) );
  XNOR U12097 ( .A(n11299), .B(n11298), .Z(n11314) );
  XOR U12098 ( .A(n11314), .B(sreg[1458]), .Z(n11295) );
  XOR U12099 ( .A(n11315), .B(n11295), .Z(c[1458]) );
  NANDN U12100 ( .A(n11297), .B(n11296), .Z(n11301) );
  NAND U12101 ( .A(n11299), .B(n11298), .Z(n11300) );
  NAND U12102 ( .A(n11301), .B(n11300), .Z(n11322) );
  AND U12103 ( .A(b[2]), .B(a[437]), .Z(n11328) );
  AND U12104 ( .A(a[438]), .B(b[1]), .Z(n11326) );
  AND U12105 ( .A(a[436]), .B(b[3]), .Z(n11325) );
  XOR U12106 ( .A(n11326), .B(n11325), .Z(n11327) );
  XOR U12107 ( .A(n11328), .B(n11327), .Z(n11331) );
  NAND U12108 ( .A(b[0]), .B(a[439]), .Z(n11332) );
  XOR U12109 ( .A(n11331), .B(n11332), .Z(n11334) );
  OR U12110 ( .A(n11303), .B(n11302), .Z(n11307) );
  NANDN U12111 ( .A(n11305), .B(n11304), .Z(n11306) );
  NAND U12112 ( .A(n11307), .B(n11306), .Z(n11333) );
  XNOR U12113 ( .A(n11334), .B(n11333), .Z(n11319) );
  NANDN U12114 ( .A(n11309), .B(n11308), .Z(n11313) );
  OR U12115 ( .A(n11311), .B(n11310), .Z(n11312) );
  NAND U12116 ( .A(n11313), .B(n11312), .Z(n11320) );
  XNOR U12117 ( .A(n11319), .B(n11320), .Z(n11321) );
  XOR U12118 ( .A(n11322), .B(n11321), .Z(n11318) );
  XOR U12119 ( .A(sreg[1459]), .B(n11317), .Z(n11316) );
  XOR U12120 ( .A(n11318), .B(n11316), .Z(c[1459]) );
  NANDN U12121 ( .A(n11320), .B(n11319), .Z(n11324) );
  NAND U12122 ( .A(n11322), .B(n11321), .Z(n11323) );
  NAND U12123 ( .A(n11324), .B(n11323), .Z(n11340) );
  AND U12124 ( .A(b[2]), .B(a[438]), .Z(n11346) );
  AND U12125 ( .A(a[439]), .B(b[1]), .Z(n11344) );
  AND U12126 ( .A(a[437]), .B(b[3]), .Z(n11343) );
  XOR U12127 ( .A(n11344), .B(n11343), .Z(n11345) );
  XOR U12128 ( .A(n11346), .B(n11345), .Z(n11349) );
  NAND U12129 ( .A(b[0]), .B(a[440]), .Z(n11350) );
  XOR U12130 ( .A(n11349), .B(n11350), .Z(n11352) );
  OR U12131 ( .A(n11326), .B(n11325), .Z(n11330) );
  NANDN U12132 ( .A(n11328), .B(n11327), .Z(n11329) );
  NAND U12133 ( .A(n11330), .B(n11329), .Z(n11351) );
  XNOR U12134 ( .A(n11352), .B(n11351), .Z(n11337) );
  NANDN U12135 ( .A(n11332), .B(n11331), .Z(n11336) );
  OR U12136 ( .A(n11334), .B(n11333), .Z(n11335) );
  NAND U12137 ( .A(n11336), .B(n11335), .Z(n11338) );
  XNOR U12138 ( .A(n11337), .B(n11338), .Z(n11339) );
  XNOR U12139 ( .A(n11340), .B(n11339), .Z(n11355) );
  XOR U12140 ( .A(sreg[1460]), .B(n11355), .Z(n11357) );
  XNOR U12141 ( .A(n11356), .B(n11357), .Z(c[1460]) );
  NANDN U12142 ( .A(n11338), .B(n11337), .Z(n11342) );
  NAND U12143 ( .A(n11340), .B(n11339), .Z(n11341) );
  NAND U12144 ( .A(n11342), .B(n11341), .Z(n11366) );
  AND U12145 ( .A(b[2]), .B(a[439]), .Z(n11372) );
  AND U12146 ( .A(a[440]), .B(b[1]), .Z(n11370) );
  AND U12147 ( .A(a[438]), .B(b[3]), .Z(n11369) );
  XOR U12148 ( .A(n11370), .B(n11369), .Z(n11371) );
  XOR U12149 ( .A(n11372), .B(n11371), .Z(n11375) );
  NAND U12150 ( .A(b[0]), .B(a[441]), .Z(n11376) );
  XOR U12151 ( .A(n11375), .B(n11376), .Z(n11378) );
  OR U12152 ( .A(n11344), .B(n11343), .Z(n11348) );
  NANDN U12153 ( .A(n11346), .B(n11345), .Z(n11347) );
  NAND U12154 ( .A(n11348), .B(n11347), .Z(n11377) );
  XNOR U12155 ( .A(n11378), .B(n11377), .Z(n11363) );
  NANDN U12156 ( .A(n11350), .B(n11349), .Z(n11354) );
  OR U12157 ( .A(n11352), .B(n11351), .Z(n11353) );
  NAND U12158 ( .A(n11354), .B(n11353), .Z(n11364) );
  XNOR U12159 ( .A(n11363), .B(n11364), .Z(n11365) );
  XOR U12160 ( .A(n11366), .B(n11365), .Z(n11362) );
  OR U12161 ( .A(n11355), .B(sreg[1460]), .Z(n11359) );
  NAND U12162 ( .A(n11357), .B(n11356), .Z(n11358) );
  AND U12163 ( .A(n11359), .B(n11358), .Z(n11361) );
  XNOR U12164 ( .A(sreg[1461]), .B(n11361), .Z(n11360) );
  XOR U12165 ( .A(n11362), .B(n11360), .Z(c[1461]) );
  NANDN U12166 ( .A(n11364), .B(n11363), .Z(n11368) );
  NAND U12167 ( .A(n11366), .B(n11365), .Z(n11367) );
  NAND U12168 ( .A(n11368), .B(n11367), .Z(n11389) );
  AND U12169 ( .A(b[2]), .B(a[440]), .Z(n11401) );
  AND U12170 ( .A(a[441]), .B(b[1]), .Z(n11399) );
  AND U12171 ( .A(a[439]), .B(b[3]), .Z(n11398) );
  XOR U12172 ( .A(n11399), .B(n11398), .Z(n11400) );
  XOR U12173 ( .A(n11401), .B(n11400), .Z(n11392) );
  NAND U12174 ( .A(b[0]), .B(a[442]), .Z(n11393) );
  XOR U12175 ( .A(n11392), .B(n11393), .Z(n11395) );
  OR U12176 ( .A(n11370), .B(n11369), .Z(n11374) );
  NANDN U12177 ( .A(n11372), .B(n11371), .Z(n11373) );
  NAND U12178 ( .A(n11374), .B(n11373), .Z(n11394) );
  XNOR U12179 ( .A(n11395), .B(n11394), .Z(n11386) );
  NANDN U12180 ( .A(n11376), .B(n11375), .Z(n11380) );
  OR U12181 ( .A(n11378), .B(n11377), .Z(n11379) );
  NAND U12182 ( .A(n11380), .B(n11379), .Z(n11387) );
  XNOR U12183 ( .A(n11386), .B(n11387), .Z(n11388) );
  XNOR U12184 ( .A(n11389), .B(n11388), .Z(n11381) );
  XNOR U12185 ( .A(n11381), .B(sreg[1462]), .Z(n11382) );
  XOR U12186 ( .A(n11383), .B(n11382), .Z(c[1462]) );
  NAND U12187 ( .A(n11381), .B(sreg[1462]), .Z(n11385) );
  OR U12188 ( .A(n11383), .B(n11382), .Z(n11384) );
  NAND U12189 ( .A(n11385), .B(n11384), .Z(n11406) );
  NANDN U12190 ( .A(n11387), .B(n11386), .Z(n11391) );
  NAND U12191 ( .A(n11389), .B(n11388), .Z(n11390) );
  AND U12192 ( .A(n11391), .B(n11390), .Z(n11410) );
  NANDN U12193 ( .A(n11393), .B(n11392), .Z(n11397) );
  OR U12194 ( .A(n11395), .B(n11394), .Z(n11396) );
  AND U12195 ( .A(n11397), .B(n11396), .Z(n11409) );
  AND U12196 ( .A(b[2]), .B(a[441]), .Z(n11414) );
  AND U12197 ( .A(a[442]), .B(b[1]), .Z(n11412) );
  AND U12198 ( .A(a[440]), .B(b[3]), .Z(n11411) );
  XOR U12199 ( .A(n11412), .B(n11411), .Z(n11413) );
  XOR U12200 ( .A(n11414), .B(n11413), .Z(n11417) );
  NAND U12201 ( .A(b[0]), .B(a[443]), .Z(n11418) );
  XOR U12202 ( .A(n11417), .B(n11418), .Z(n11420) );
  OR U12203 ( .A(n11399), .B(n11398), .Z(n11403) );
  NANDN U12204 ( .A(n11401), .B(n11400), .Z(n11402) );
  NAND U12205 ( .A(n11403), .B(n11402), .Z(n11419) );
  XOR U12206 ( .A(n11420), .B(n11419), .Z(n11408) );
  XNOR U12207 ( .A(n11409), .B(n11408), .Z(n11404) );
  XOR U12208 ( .A(n11410), .B(n11404), .Z(n11407) );
  XNOR U12209 ( .A(sreg[1463]), .B(n11407), .Z(n11405) );
  XNOR U12210 ( .A(n11406), .B(n11405), .Z(c[1463]) );
  AND U12211 ( .A(b[2]), .B(a[442]), .Z(n11432) );
  AND U12212 ( .A(a[443]), .B(b[1]), .Z(n11430) );
  AND U12213 ( .A(a[441]), .B(b[3]), .Z(n11429) );
  XOR U12214 ( .A(n11430), .B(n11429), .Z(n11431) );
  XOR U12215 ( .A(n11432), .B(n11431), .Z(n11435) );
  NAND U12216 ( .A(b[0]), .B(a[444]), .Z(n11436) );
  XOR U12217 ( .A(n11435), .B(n11436), .Z(n11438) );
  OR U12218 ( .A(n11412), .B(n11411), .Z(n11416) );
  NANDN U12219 ( .A(n11414), .B(n11413), .Z(n11415) );
  NAND U12220 ( .A(n11416), .B(n11415), .Z(n11437) );
  XNOR U12221 ( .A(n11438), .B(n11437), .Z(n11423) );
  NANDN U12222 ( .A(n11418), .B(n11417), .Z(n11422) );
  OR U12223 ( .A(n11420), .B(n11419), .Z(n11421) );
  NAND U12224 ( .A(n11422), .B(n11421), .Z(n11424) );
  XNOR U12225 ( .A(n11423), .B(n11424), .Z(n11425) );
  XOR U12226 ( .A(n11426), .B(n11425), .Z(n11441) );
  XNOR U12227 ( .A(n11441), .B(sreg[1464]), .Z(n11442) );
  XOR U12228 ( .A(n11443), .B(n11442), .Z(c[1464]) );
  NANDN U12229 ( .A(n11424), .B(n11423), .Z(n11428) );
  NANDN U12230 ( .A(n11426), .B(n11425), .Z(n11427) );
  NAND U12231 ( .A(n11428), .B(n11427), .Z(n11454) );
  AND U12232 ( .A(b[2]), .B(a[443]), .Z(n11460) );
  AND U12233 ( .A(a[444]), .B(b[1]), .Z(n11458) );
  AND U12234 ( .A(a[442]), .B(b[3]), .Z(n11457) );
  XOR U12235 ( .A(n11458), .B(n11457), .Z(n11459) );
  XOR U12236 ( .A(n11460), .B(n11459), .Z(n11463) );
  NAND U12237 ( .A(b[0]), .B(a[445]), .Z(n11464) );
  XOR U12238 ( .A(n11463), .B(n11464), .Z(n11466) );
  OR U12239 ( .A(n11430), .B(n11429), .Z(n11434) );
  NANDN U12240 ( .A(n11432), .B(n11431), .Z(n11433) );
  NAND U12241 ( .A(n11434), .B(n11433), .Z(n11465) );
  XNOR U12242 ( .A(n11466), .B(n11465), .Z(n11451) );
  NANDN U12243 ( .A(n11436), .B(n11435), .Z(n11440) );
  OR U12244 ( .A(n11438), .B(n11437), .Z(n11439) );
  NAND U12245 ( .A(n11440), .B(n11439), .Z(n11452) );
  XNOR U12246 ( .A(n11451), .B(n11452), .Z(n11453) );
  XNOR U12247 ( .A(n11454), .B(n11453), .Z(n11446) );
  XNOR U12248 ( .A(n11446), .B(sreg[1465]), .Z(n11448) );
  NAND U12249 ( .A(n11441), .B(sreg[1464]), .Z(n11445) );
  OR U12250 ( .A(n11443), .B(n11442), .Z(n11444) );
  AND U12251 ( .A(n11445), .B(n11444), .Z(n11447) );
  XOR U12252 ( .A(n11448), .B(n11447), .Z(c[1465]) );
  NAND U12253 ( .A(n11446), .B(sreg[1465]), .Z(n11450) );
  OR U12254 ( .A(n11448), .B(n11447), .Z(n11449) );
  NAND U12255 ( .A(n11450), .B(n11449), .Z(n11471) );
  NANDN U12256 ( .A(n11452), .B(n11451), .Z(n11456) );
  NAND U12257 ( .A(n11454), .B(n11453), .Z(n11455) );
  AND U12258 ( .A(n11456), .B(n11455), .Z(n11475) );
  AND U12259 ( .A(b[2]), .B(a[444]), .Z(n11479) );
  AND U12260 ( .A(a[445]), .B(b[1]), .Z(n11477) );
  AND U12261 ( .A(a[443]), .B(b[3]), .Z(n11476) );
  XOR U12262 ( .A(n11477), .B(n11476), .Z(n11478) );
  XOR U12263 ( .A(n11479), .B(n11478), .Z(n11482) );
  NAND U12264 ( .A(b[0]), .B(a[446]), .Z(n11483) );
  XOR U12265 ( .A(n11482), .B(n11483), .Z(n11484) );
  OR U12266 ( .A(n11458), .B(n11457), .Z(n11462) );
  NANDN U12267 ( .A(n11460), .B(n11459), .Z(n11461) );
  AND U12268 ( .A(n11462), .B(n11461), .Z(n11485) );
  XOR U12269 ( .A(n11484), .B(n11485), .Z(n11473) );
  NANDN U12270 ( .A(n11464), .B(n11463), .Z(n11468) );
  OR U12271 ( .A(n11466), .B(n11465), .Z(n11467) );
  AND U12272 ( .A(n11468), .B(n11467), .Z(n11474) );
  XOR U12273 ( .A(n11473), .B(n11474), .Z(n11469) );
  XNOR U12274 ( .A(n11475), .B(n11469), .Z(n11472) );
  XOR U12275 ( .A(sreg[1466]), .B(n11472), .Z(n11470) );
  XNOR U12276 ( .A(n11471), .B(n11470), .Z(c[1466]) );
  AND U12277 ( .A(b[2]), .B(a[445]), .Z(n11495) );
  AND U12278 ( .A(a[446]), .B(b[1]), .Z(n11493) );
  AND U12279 ( .A(a[444]), .B(b[3]), .Z(n11492) );
  XOR U12280 ( .A(n11493), .B(n11492), .Z(n11494) );
  XOR U12281 ( .A(n11495), .B(n11494), .Z(n11498) );
  NAND U12282 ( .A(b[0]), .B(a[447]), .Z(n11499) );
  XOR U12283 ( .A(n11498), .B(n11499), .Z(n11501) );
  OR U12284 ( .A(n11477), .B(n11476), .Z(n11481) );
  NANDN U12285 ( .A(n11479), .B(n11478), .Z(n11480) );
  NAND U12286 ( .A(n11481), .B(n11480), .Z(n11500) );
  XNOR U12287 ( .A(n11501), .B(n11500), .Z(n11486) );
  XNOR U12288 ( .A(n11486), .B(n11487), .Z(n11489) );
  XOR U12289 ( .A(n11488), .B(n11489), .Z(n11504) );
  XOR U12290 ( .A(n11504), .B(sreg[1467]), .Z(n11505) );
  XOR U12291 ( .A(n11506), .B(n11505), .Z(c[1467]) );
  NANDN U12292 ( .A(n11487), .B(n11486), .Z(n11491) );
  NAND U12293 ( .A(n11489), .B(n11488), .Z(n11490) );
  NAND U12294 ( .A(n11491), .B(n11490), .Z(n11512) );
  AND U12295 ( .A(b[2]), .B(a[446]), .Z(n11524) );
  AND U12296 ( .A(a[447]), .B(b[1]), .Z(n11522) );
  AND U12297 ( .A(a[445]), .B(b[3]), .Z(n11521) );
  XOR U12298 ( .A(n11522), .B(n11521), .Z(n11523) );
  XOR U12299 ( .A(n11524), .B(n11523), .Z(n11515) );
  NAND U12300 ( .A(b[0]), .B(a[448]), .Z(n11516) );
  XOR U12301 ( .A(n11515), .B(n11516), .Z(n11518) );
  OR U12302 ( .A(n11493), .B(n11492), .Z(n11497) );
  NANDN U12303 ( .A(n11495), .B(n11494), .Z(n11496) );
  NAND U12304 ( .A(n11497), .B(n11496), .Z(n11517) );
  XNOR U12305 ( .A(n11518), .B(n11517), .Z(n11509) );
  NANDN U12306 ( .A(n11499), .B(n11498), .Z(n11503) );
  OR U12307 ( .A(n11501), .B(n11500), .Z(n11502) );
  NAND U12308 ( .A(n11503), .B(n11502), .Z(n11510) );
  XNOR U12309 ( .A(n11509), .B(n11510), .Z(n11511) );
  XNOR U12310 ( .A(n11512), .B(n11511), .Z(n11528) );
  XOR U12311 ( .A(sreg[1468]), .B(n11528), .Z(n11529) );
  NANDN U12312 ( .A(n11504), .B(sreg[1467]), .Z(n11508) );
  OR U12313 ( .A(n11506), .B(n11505), .Z(n11507) );
  NAND U12314 ( .A(n11508), .B(n11507), .Z(n11530) );
  XOR U12315 ( .A(n11529), .B(n11530), .Z(c[1468]) );
  NANDN U12316 ( .A(n11510), .B(n11509), .Z(n11514) );
  NAND U12317 ( .A(n11512), .B(n11511), .Z(n11513) );
  AND U12318 ( .A(n11514), .B(n11513), .Z(n11536) );
  NANDN U12319 ( .A(n11516), .B(n11515), .Z(n11520) );
  OR U12320 ( .A(n11518), .B(n11517), .Z(n11519) );
  AND U12321 ( .A(n11520), .B(n11519), .Z(n11535) );
  AND U12322 ( .A(b[2]), .B(a[447]), .Z(n11540) );
  AND U12323 ( .A(a[448]), .B(b[1]), .Z(n11538) );
  AND U12324 ( .A(a[446]), .B(b[3]), .Z(n11537) );
  XOR U12325 ( .A(n11538), .B(n11537), .Z(n11539) );
  XOR U12326 ( .A(n11540), .B(n11539), .Z(n11543) );
  NAND U12327 ( .A(b[0]), .B(a[449]), .Z(n11544) );
  XOR U12328 ( .A(n11543), .B(n11544), .Z(n11546) );
  OR U12329 ( .A(n11522), .B(n11521), .Z(n11526) );
  NANDN U12330 ( .A(n11524), .B(n11523), .Z(n11525) );
  NAND U12331 ( .A(n11526), .B(n11525), .Z(n11545) );
  XOR U12332 ( .A(n11546), .B(n11545), .Z(n11534) );
  XNOR U12333 ( .A(n11535), .B(n11534), .Z(n11527) );
  XOR U12334 ( .A(n11536), .B(n11527), .Z(n11550) );
  OR U12335 ( .A(n11528), .B(sreg[1468]), .Z(n11532) );
  NANDN U12336 ( .A(n11530), .B(n11529), .Z(n11531) );
  AND U12337 ( .A(n11532), .B(n11531), .Z(n11549) );
  XNOR U12338 ( .A(sreg[1469]), .B(n11549), .Z(n11533) );
  XNOR U12339 ( .A(n11550), .B(n11533), .Z(c[1469]) );
  AND U12340 ( .A(b[2]), .B(a[448]), .Z(n11561) );
  AND U12341 ( .A(a[449]), .B(b[1]), .Z(n11559) );
  AND U12342 ( .A(a[447]), .B(b[3]), .Z(n11558) );
  XOR U12343 ( .A(n11559), .B(n11558), .Z(n11560) );
  XOR U12344 ( .A(n11561), .B(n11560), .Z(n11564) );
  NAND U12345 ( .A(b[0]), .B(a[450]), .Z(n11565) );
  XOR U12346 ( .A(n11564), .B(n11565), .Z(n11567) );
  OR U12347 ( .A(n11538), .B(n11537), .Z(n11542) );
  NANDN U12348 ( .A(n11540), .B(n11539), .Z(n11541) );
  NAND U12349 ( .A(n11542), .B(n11541), .Z(n11566) );
  XNOR U12350 ( .A(n11567), .B(n11566), .Z(n11552) );
  NANDN U12351 ( .A(n11544), .B(n11543), .Z(n11548) );
  OR U12352 ( .A(n11546), .B(n11545), .Z(n11547) );
  NAND U12353 ( .A(n11548), .B(n11547), .Z(n11553) );
  XNOR U12354 ( .A(n11552), .B(n11553), .Z(n11554) );
  XOR U12355 ( .A(n11555), .B(n11554), .Z(n11571) );
  XNOR U12356 ( .A(sreg[1470]), .B(n11570), .Z(n11551) );
  XNOR U12357 ( .A(n11571), .B(n11551), .Z(c[1470]) );
  NANDN U12358 ( .A(n11553), .B(n11552), .Z(n11557) );
  NANDN U12359 ( .A(n11555), .B(n11554), .Z(n11556) );
  NAND U12360 ( .A(n11557), .B(n11556), .Z(n11576) );
  AND U12361 ( .A(b[2]), .B(a[449]), .Z(n11582) );
  AND U12362 ( .A(a[450]), .B(b[1]), .Z(n11580) );
  AND U12363 ( .A(a[448]), .B(b[3]), .Z(n11579) );
  XOR U12364 ( .A(n11580), .B(n11579), .Z(n11581) );
  XOR U12365 ( .A(n11582), .B(n11581), .Z(n11585) );
  NAND U12366 ( .A(b[0]), .B(a[451]), .Z(n11586) );
  XOR U12367 ( .A(n11585), .B(n11586), .Z(n11588) );
  OR U12368 ( .A(n11559), .B(n11558), .Z(n11563) );
  NANDN U12369 ( .A(n11561), .B(n11560), .Z(n11562) );
  NAND U12370 ( .A(n11563), .B(n11562), .Z(n11587) );
  XNOR U12371 ( .A(n11588), .B(n11587), .Z(n11573) );
  NANDN U12372 ( .A(n11565), .B(n11564), .Z(n11569) );
  OR U12373 ( .A(n11567), .B(n11566), .Z(n11568) );
  NAND U12374 ( .A(n11569), .B(n11568), .Z(n11574) );
  XNOR U12375 ( .A(n11573), .B(n11574), .Z(n11575) );
  XOR U12376 ( .A(n11576), .B(n11575), .Z(n11593) );
  XNOR U12377 ( .A(sreg[1471]), .B(n11592), .Z(n11572) );
  XOR U12378 ( .A(n11593), .B(n11572), .Z(c[1471]) );
  NANDN U12379 ( .A(n11574), .B(n11573), .Z(n11578) );
  NAND U12380 ( .A(n11576), .B(n11575), .Z(n11577) );
  AND U12381 ( .A(n11578), .B(n11577), .Z(n11599) );
  AND U12382 ( .A(b[2]), .B(a[450]), .Z(n11607) );
  AND U12383 ( .A(a[451]), .B(b[1]), .Z(n11605) );
  AND U12384 ( .A(a[449]), .B(b[3]), .Z(n11604) );
  XOR U12385 ( .A(n11605), .B(n11604), .Z(n11606) );
  XOR U12386 ( .A(n11607), .B(n11606), .Z(n11600) );
  NAND U12387 ( .A(b[0]), .B(a[452]), .Z(n11601) );
  XOR U12388 ( .A(n11600), .B(n11601), .Z(n11602) );
  OR U12389 ( .A(n11580), .B(n11579), .Z(n11584) );
  NANDN U12390 ( .A(n11582), .B(n11581), .Z(n11583) );
  AND U12391 ( .A(n11584), .B(n11583), .Z(n11603) );
  XOR U12392 ( .A(n11602), .B(n11603), .Z(n11597) );
  NANDN U12393 ( .A(n11586), .B(n11585), .Z(n11590) );
  OR U12394 ( .A(n11588), .B(n11587), .Z(n11589) );
  AND U12395 ( .A(n11590), .B(n11589), .Z(n11598) );
  XOR U12396 ( .A(n11597), .B(n11598), .Z(n11591) );
  XNOR U12397 ( .A(n11599), .B(n11591), .Z(n11596) );
  XNOR U12398 ( .A(sreg[1472]), .B(n11595), .Z(n11594) );
  XOR U12399 ( .A(n11596), .B(n11594), .Z(c[1472]) );
  AND U12400 ( .A(b[2]), .B(a[451]), .Z(n11613) );
  AND U12401 ( .A(a[452]), .B(b[1]), .Z(n11611) );
  AND U12402 ( .A(a[450]), .B(b[3]), .Z(n11610) );
  XOR U12403 ( .A(n11611), .B(n11610), .Z(n11612) );
  XOR U12404 ( .A(n11613), .B(n11612), .Z(n11616) );
  NAND U12405 ( .A(b[0]), .B(a[453]), .Z(n11617) );
  XNOR U12406 ( .A(n11616), .B(n11617), .Z(n11618) );
  OR U12407 ( .A(n11605), .B(n11604), .Z(n11609) );
  NANDN U12408 ( .A(n11607), .B(n11606), .Z(n11608) );
  AND U12409 ( .A(n11609), .B(n11608), .Z(n11619) );
  XNOR U12410 ( .A(n11618), .B(n11619), .Z(n11623) );
  XNOR U12411 ( .A(n11622), .B(n11623), .Z(n11624) );
  XNOR U12412 ( .A(n11625), .B(n11624), .Z(n11628) );
  XNOR U12413 ( .A(sreg[1473]), .B(n11628), .Z(n11629) );
  XOR U12414 ( .A(n11630), .B(n11629), .Z(c[1473]) );
  AND U12415 ( .A(b[2]), .B(a[452]), .Z(n11642) );
  AND U12416 ( .A(a[453]), .B(b[1]), .Z(n11640) );
  AND U12417 ( .A(a[451]), .B(b[3]), .Z(n11639) );
  XOR U12418 ( .A(n11640), .B(n11639), .Z(n11641) );
  XOR U12419 ( .A(n11642), .B(n11641), .Z(n11645) );
  NAND U12420 ( .A(b[0]), .B(a[454]), .Z(n11646) );
  XOR U12421 ( .A(n11645), .B(n11646), .Z(n11648) );
  OR U12422 ( .A(n11611), .B(n11610), .Z(n11615) );
  NANDN U12423 ( .A(n11613), .B(n11612), .Z(n11614) );
  NAND U12424 ( .A(n11615), .B(n11614), .Z(n11647) );
  XNOR U12425 ( .A(n11648), .B(n11647), .Z(n11633) );
  NANDN U12426 ( .A(n11617), .B(n11616), .Z(n11621) );
  NAND U12427 ( .A(n11619), .B(n11618), .Z(n11620) );
  NAND U12428 ( .A(n11621), .B(n11620), .Z(n11634) );
  XNOR U12429 ( .A(n11633), .B(n11634), .Z(n11635) );
  NANDN U12430 ( .A(n11623), .B(n11622), .Z(n11627) );
  NANDN U12431 ( .A(n11625), .B(n11624), .Z(n11626) );
  NAND U12432 ( .A(n11627), .B(n11626), .Z(n11636) );
  XOR U12433 ( .A(n11635), .B(n11636), .Z(n11651) );
  XNOR U12434 ( .A(n11651), .B(sreg[1474]), .Z(n11653) );
  NAND U12435 ( .A(sreg[1473]), .B(n11628), .Z(n11632) );
  OR U12436 ( .A(n11630), .B(n11629), .Z(n11631) );
  AND U12437 ( .A(n11632), .B(n11631), .Z(n11652) );
  XOR U12438 ( .A(n11653), .B(n11652), .Z(c[1474]) );
  NANDN U12439 ( .A(n11634), .B(n11633), .Z(n11638) );
  NANDN U12440 ( .A(n11636), .B(n11635), .Z(n11637) );
  NAND U12441 ( .A(n11638), .B(n11637), .Z(n11674) );
  AND U12442 ( .A(b[2]), .B(a[453]), .Z(n11668) );
  AND U12443 ( .A(a[454]), .B(b[1]), .Z(n11666) );
  AND U12444 ( .A(a[452]), .B(b[3]), .Z(n11665) );
  XOR U12445 ( .A(n11666), .B(n11665), .Z(n11667) );
  XOR U12446 ( .A(n11668), .B(n11667), .Z(n11659) );
  NAND U12447 ( .A(b[0]), .B(a[455]), .Z(n11660) );
  XOR U12448 ( .A(n11659), .B(n11660), .Z(n11662) );
  OR U12449 ( .A(n11640), .B(n11639), .Z(n11644) );
  NANDN U12450 ( .A(n11642), .B(n11641), .Z(n11643) );
  NAND U12451 ( .A(n11644), .B(n11643), .Z(n11661) );
  XNOR U12452 ( .A(n11662), .B(n11661), .Z(n11671) );
  NANDN U12453 ( .A(n11646), .B(n11645), .Z(n11650) );
  OR U12454 ( .A(n11648), .B(n11647), .Z(n11649) );
  NAND U12455 ( .A(n11650), .B(n11649), .Z(n11672) );
  XNOR U12456 ( .A(n11671), .B(n11672), .Z(n11673) );
  XOR U12457 ( .A(n11674), .B(n11673), .Z(n11658) );
  NAND U12458 ( .A(n11651), .B(sreg[1474]), .Z(n11655) );
  OR U12459 ( .A(n11653), .B(n11652), .Z(n11654) );
  NAND U12460 ( .A(n11655), .B(n11654), .Z(n11657) );
  XNOR U12461 ( .A(sreg[1475]), .B(n11657), .Z(n11656) );
  XOR U12462 ( .A(n11658), .B(n11656), .Z(c[1475]) );
  NANDN U12463 ( .A(n11660), .B(n11659), .Z(n11664) );
  OR U12464 ( .A(n11662), .B(n11661), .Z(n11663) );
  NAND U12465 ( .A(n11664), .B(n11663), .Z(n11689) );
  AND U12466 ( .A(b[2]), .B(a[454]), .Z(n11680) );
  AND U12467 ( .A(a[455]), .B(b[1]), .Z(n11678) );
  AND U12468 ( .A(a[453]), .B(b[3]), .Z(n11677) );
  XOR U12469 ( .A(n11678), .B(n11677), .Z(n11679) );
  XOR U12470 ( .A(n11680), .B(n11679), .Z(n11683) );
  NAND U12471 ( .A(b[0]), .B(a[456]), .Z(n11684) );
  XNOR U12472 ( .A(n11683), .B(n11684), .Z(n11685) );
  OR U12473 ( .A(n11666), .B(n11665), .Z(n11670) );
  NANDN U12474 ( .A(n11668), .B(n11667), .Z(n11669) );
  AND U12475 ( .A(n11670), .B(n11669), .Z(n11686) );
  XNOR U12476 ( .A(n11685), .B(n11686), .Z(n11690) );
  XNOR U12477 ( .A(n11689), .B(n11690), .Z(n11691) );
  NANDN U12478 ( .A(n11672), .B(n11671), .Z(n11676) );
  NAND U12479 ( .A(n11674), .B(n11673), .Z(n11675) );
  AND U12480 ( .A(n11676), .B(n11675), .Z(n11692) );
  XOR U12481 ( .A(n11691), .B(n11692), .Z(n11695) );
  XNOR U12482 ( .A(sreg[1476]), .B(n11695), .Z(n11696) );
  XOR U12483 ( .A(n11697), .B(n11696), .Z(c[1476]) );
  AND U12484 ( .A(b[2]), .B(a[455]), .Z(n11712) );
  AND U12485 ( .A(a[456]), .B(b[1]), .Z(n11710) );
  AND U12486 ( .A(a[454]), .B(b[3]), .Z(n11709) );
  XOR U12487 ( .A(n11710), .B(n11709), .Z(n11711) );
  XOR U12488 ( .A(n11712), .B(n11711), .Z(n11715) );
  NAND U12489 ( .A(b[0]), .B(a[457]), .Z(n11716) );
  XOR U12490 ( .A(n11715), .B(n11716), .Z(n11718) );
  OR U12491 ( .A(n11678), .B(n11677), .Z(n11682) );
  NANDN U12492 ( .A(n11680), .B(n11679), .Z(n11681) );
  NAND U12493 ( .A(n11682), .B(n11681), .Z(n11717) );
  XNOR U12494 ( .A(n11718), .B(n11717), .Z(n11703) );
  NANDN U12495 ( .A(n11684), .B(n11683), .Z(n11688) );
  NAND U12496 ( .A(n11686), .B(n11685), .Z(n11687) );
  NAND U12497 ( .A(n11688), .B(n11687), .Z(n11704) );
  XNOR U12498 ( .A(n11703), .B(n11704), .Z(n11705) );
  NANDN U12499 ( .A(n11690), .B(n11689), .Z(n11694) );
  NAND U12500 ( .A(n11692), .B(n11691), .Z(n11693) );
  AND U12501 ( .A(n11694), .B(n11693), .Z(n11706) );
  XNOR U12502 ( .A(n11705), .B(n11706), .Z(n11702) );
  NAND U12503 ( .A(sreg[1476]), .B(n11695), .Z(n11699) );
  OR U12504 ( .A(n11697), .B(n11696), .Z(n11698) );
  AND U12505 ( .A(n11699), .B(n11698), .Z(n11701) );
  XNOR U12506 ( .A(n11701), .B(sreg[1477]), .Z(n11700) );
  XOR U12507 ( .A(n11702), .B(n11700), .Z(c[1477]) );
  NANDN U12508 ( .A(n11704), .B(n11703), .Z(n11708) );
  NAND U12509 ( .A(n11706), .B(n11705), .Z(n11707) );
  NAND U12510 ( .A(n11708), .B(n11707), .Z(n11729) );
  AND U12511 ( .A(b[2]), .B(a[456]), .Z(n11735) );
  AND U12512 ( .A(a[457]), .B(b[1]), .Z(n11733) );
  AND U12513 ( .A(a[455]), .B(b[3]), .Z(n11732) );
  XOR U12514 ( .A(n11733), .B(n11732), .Z(n11734) );
  XOR U12515 ( .A(n11735), .B(n11734), .Z(n11738) );
  NAND U12516 ( .A(b[0]), .B(a[458]), .Z(n11739) );
  XOR U12517 ( .A(n11738), .B(n11739), .Z(n11741) );
  OR U12518 ( .A(n11710), .B(n11709), .Z(n11714) );
  NANDN U12519 ( .A(n11712), .B(n11711), .Z(n11713) );
  NAND U12520 ( .A(n11714), .B(n11713), .Z(n11740) );
  XNOR U12521 ( .A(n11741), .B(n11740), .Z(n11726) );
  NANDN U12522 ( .A(n11716), .B(n11715), .Z(n11720) );
  OR U12523 ( .A(n11718), .B(n11717), .Z(n11719) );
  NAND U12524 ( .A(n11720), .B(n11719), .Z(n11727) );
  XNOR U12525 ( .A(n11726), .B(n11727), .Z(n11728) );
  XNOR U12526 ( .A(n11729), .B(n11728), .Z(n11721) );
  XOR U12527 ( .A(sreg[1478]), .B(n11721), .Z(n11722) );
  XOR U12528 ( .A(n11723), .B(n11722), .Z(c[1478]) );
  OR U12529 ( .A(n11721), .B(sreg[1478]), .Z(n11725) );
  NANDN U12530 ( .A(n11723), .B(n11722), .Z(n11724) );
  NAND U12531 ( .A(n11725), .B(n11724), .Z(n11764) );
  NANDN U12532 ( .A(n11727), .B(n11726), .Z(n11731) );
  NAND U12533 ( .A(n11729), .B(n11728), .Z(n11730) );
  NAND U12534 ( .A(n11731), .B(n11730), .Z(n11747) );
  AND U12535 ( .A(b[2]), .B(a[457]), .Z(n11753) );
  AND U12536 ( .A(a[458]), .B(b[1]), .Z(n11751) );
  AND U12537 ( .A(a[456]), .B(b[3]), .Z(n11750) );
  XOR U12538 ( .A(n11751), .B(n11750), .Z(n11752) );
  XOR U12539 ( .A(n11753), .B(n11752), .Z(n11756) );
  NAND U12540 ( .A(b[0]), .B(a[459]), .Z(n11757) );
  XOR U12541 ( .A(n11756), .B(n11757), .Z(n11759) );
  OR U12542 ( .A(n11733), .B(n11732), .Z(n11737) );
  NANDN U12543 ( .A(n11735), .B(n11734), .Z(n11736) );
  NAND U12544 ( .A(n11737), .B(n11736), .Z(n11758) );
  XNOR U12545 ( .A(n11759), .B(n11758), .Z(n11744) );
  NANDN U12546 ( .A(n11739), .B(n11738), .Z(n11743) );
  OR U12547 ( .A(n11741), .B(n11740), .Z(n11742) );
  NAND U12548 ( .A(n11743), .B(n11742), .Z(n11745) );
  XNOR U12549 ( .A(n11744), .B(n11745), .Z(n11746) );
  XNOR U12550 ( .A(n11747), .B(n11746), .Z(n11762) );
  XNOR U12551 ( .A(n11762), .B(sreg[1479]), .Z(n11763) );
  XOR U12552 ( .A(n11764), .B(n11763), .Z(c[1479]) );
  NANDN U12553 ( .A(n11745), .B(n11744), .Z(n11749) );
  NAND U12554 ( .A(n11747), .B(n11746), .Z(n11748) );
  NAND U12555 ( .A(n11749), .B(n11748), .Z(n11770) );
  AND U12556 ( .A(b[2]), .B(a[458]), .Z(n11776) );
  AND U12557 ( .A(a[459]), .B(b[1]), .Z(n11774) );
  AND U12558 ( .A(a[457]), .B(b[3]), .Z(n11773) );
  XOR U12559 ( .A(n11774), .B(n11773), .Z(n11775) );
  XOR U12560 ( .A(n11776), .B(n11775), .Z(n11779) );
  NAND U12561 ( .A(b[0]), .B(a[460]), .Z(n11780) );
  XOR U12562 ( .A(n11779), .B(n11780), .Z(n11782) );
  OR U12563 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U12564 ( .A(n11753), .B(n11752), .Z(n11754) );
  NAND U12565 ( .A(n11755), .B(n11754), .Z(n11781) );
  XNOR U12566 ( .A(n11782), .B(n11781), .Z(n11767) );
  NANDN U12567 ( .A(n11757), .B(n11756), .Z(n11761) );
  OR U12568 ( .A(n11759), .B(n11758), .Z(n11760) );
  NAND U12569 ( .A(n11761), .B(n11760), .Z(n11768) );
  XNOR U12570 ( .A(n11767), .B(n11768), .Z(n11769) );
  XNOR U12571 ( .A(n11770), .B(n11769), .Z(n11785) );
  XOR U12572 ( .A(sreg[1480]), .B(n11785), .Z(n11786) );
  NAND U12573 ( .A(n11762), .B(sreg[1479]), .Z(n11766) );
  OR U12574 ( .A(n11764), .B(n11763), .Z(n11765) );
  NAND U12575 ( .A(n11766), .B(n11765), .Z(n11787) );
  XOR U12576 ( .A(n11786), .B(n11787), .Z(c[1480]) );
  NANDN U12577 ( .A(n11768), .B(n11767), .Z(n11772) );
  NAND U12578 ( .A(n11770), .B(n11769), .Z(n11771) );
  NAND U12579 ( .A(n11772), .B(n11771), .Z(n11798) );
  AND U12580 ( .A(b[2]), .B(a[459]), .Z(n11804) );
  AND U12581 ( .A(a[460]), .B(b[1]), .Z(n11802) );
  AND U12582 ( .A(a[458]), .B(b[3]), .Z(n11801) );
  XOR U12583 ( .A(n11802), .B(n11801), .Z(n11803) );
  XOR U12584 ( .A(n11804), .B(n11803), .Z(n11807) );
  NAND U12585 ( .A(b[0]), .B(a[461]), .Z(n11808) );
  XOR U12586 ( .A(n11807), .B(n11808), .Z(n11810) );
  OR U12587 ( .A(n11774), .B(n11773), .Z(n11778) );
  NANDN U12588 ( .A(n11776), .B(n11775), .Z(n11777) );
  NAND U12589 ( .A(n11778), .B(n11777), .Z(n11809) );
  XNOR U12590 ( .A(n11810), .B(n11809), .Z(n11795) );
  NANDN U12591 ( .A(n11780), .B(n11779), .Z(n11784) );
  OR U12592 ( .A(n11782), .B(n11781), .Z(n11783) );
  NAND U12593 ( .A(n11784), .B(n11783), .Z(n11796) );
  XNOR U12594 ( .A(n11795), .B(n11796), .Z(n11797) );
  XNOR U12595 ( .A(n11798), .B(n11797), .Z(n11790) );
  XOR U12596 ( .A(sreg[1481]), .B(n11790), .Z(n11791) );
  OR U12597 ( .A(n11785), .B(sreg[1480]), .Z(n11789) );
  NANDN U12598 ( .A(n11787), .B(n11786), .Z(n11788) );
  AND U12599 ( .A(n11789), .B(n11788), .Z(n11792) );
  XOR U12600 ( .A(n11791), .B(n11792), .Z(c[1481]) );
  OR U12601 ( .A(n11790), .B(sreg[1481]), .Z(n11794) );
  NANDN U12602 ( .A(n11792), .B(n11791), .Z(n11793) );
  NAND U12603 ( .A(n11794), .B(n11793), .Z(n11815) );
  NANDN U12604 ( .A(n11796), .B(n11795), .Z(n11800) );
  NAND U12605 ( .A(n11798), .B(n11797), .Z(n11799) );
  NAND U12606 ( .A(n11800), .B(n11799), .Z(n11821) );
  AND U12607 ( .A(b[2]), .B(a[460]), .Z(n11827) );
  AND U12608 ( .A(a[461]), .B(b[1]), .Z(n11825) );
  AND U12609 ( .A(a[459]), .B(b[3]), .Z(n11824) );
  XOR U12610 ( .A(n11825), .B(n11824), .Z(n11826) );
  XOR U12611 ( .A(n11827), .B(n11826), .Z(n11830) );
  NAND U12612 ( .A(b[0]), .B(a[462]), .Z(n11831) );
  XOR U12613 ( .A(n11830), .B(n11831), .Z(n11833) );
  OR U12614 ( .A(n11802), .B(n11801), .Z(n11806) );
  NANDN U12615 ( .A(n11804), .B(n11803), .Z(n11805) );
  NAND U12616 ( .A(n11806), .B(n11805), .Z(n11832) );
  XNOR U12617 ( .A(n11833), .B(n11832), .Z(n11818) );
  NANDN U12618 ( .A(n11808), .B(n11807), .Z(n11812) );
  OR U12619 ( .A(n11810), .B(n11809), .Z(n11811) );
  NAND U12620 ( .A(n11812), .B(n11811), .Z(n11819) );
  XNOR U12621 ( .A(n11818), .B(n11819), .Z(n11820) );
  XNOR U12622 ( .A(n11821), .B(n11820), .Z(n11813) );
  XNOR U12623 ( .A(n11813), .B(sreg[1482]), .Z(n11814) );
  XOR U12624 ( .A(n11815), .B(n11814), .Z(c[1482]) );
  NAND U12625 ( .A(n11813), .B(sreg[1482]), .Z(n11817) );
  OR U12626 ( .A(n11815), .B(n11814), .Z(n11816) );
  NAND U12627 ( .A(n11817), .B(n11816), .Z(n11856) );
  NANDN U12628 ( .A(n11819), .B(n11818), .Z(n11823) );
  NAND U12629 ( .A(n11821), .B(n11820), .Z(n11822) );
  NAND U12630 ( .A(n11823), .B(n11822), .Z(n11839) );
  AND U12631 ( .A(b[2]), .B(a[461]), .Z(n11845) );
  AND U12632 ( .A(a[462]), .B(b[1]), .Z(n11843) );
  AND U12633 ( .A(a[460]), .B(b[3]), .Z(n11842) );
  XOR U12634 ( .A(n11843), .B(n11842), .Z(n11844) );
  XOR U12635 ( .A(n11845), .B(n11844), .Z(n11848) );
  NAND U12636 ( .A(b[0]), .B(a[463]), .Z(n11849) );
  XOR U12637 ( .A(n11848), .B(n11849), .Z(n11851) );
  OR U12638 ( .A(n11825), .B(n11824), .Z(n11829) );
  NANDN U12639 ( .A(n11827), .B(n11826), .Z(n11828) );
  NAND U12640 ( .A(n11829), .B(n11828), .Z(n11850) );
  XNOR U12641 ( .A(n11851), .B(n11850), .Z(n11836) );
  NANDN U12642 ( .A(n11831), .B(n11830), .Z(n11835) );
  OR U12643 ( .A(n11833), .B(n11832), .Z(n11834) );
  NAND U12644 ( .A(n11835), .B(n11834), .Z(n11837) );
  XNOR U12645 ( .A(n11836), .B(n11837), .Z(n11838) );
  XNOR U12646 ( .A(n11839), .B(n11838), .Z(n11854) );
  XOR U12647 ( .A(sreg[1483]), .B(n11854), .Z(n11855) );
  XOR U12648 ( .A(n11856), .B(n11855), .Z(c[1483]) );
  NANDN U12649 ( .A(n11837), .B(n11836), .Z(n11841) );
  NAND U12650 ( .A(n11839), .B(n11838), .Z(n11840) );
  NAND U12651 ( .A(n11841), .B(n11840), .Z(n11867) );
  AND U12652 ( .A(b[2]), .B(a[462]), .Z(n11873) );
  AND U12653 ( .A(a[463]), .B(b[1]), .Z(n11871) );
  AND U12654 ( .A(a[461]), .B(b[3]), .Z(n11870) );
  XOR U12655 ( .A(n11871), .B(n11870), .Z(n11872) );
  XOR U12656 ( .A(n11873), .B(n11872), .Z(n11876) );
  NAND U12657 ( .A(b[0]), .B(a[464]), .Z(n11877) );
  XOR U12658 ( .A(n11876), .B(n11877), .Z(n11879) );
  OR U12659 ( .A(n11843), .B(n11842), .Z(n11847) );
  NANDN U12660 ( .A(n11845), .B(n11844), .Z(n11846) );
  NAND U12661 ( .A(n11847), .B(n11846), .Z(n11878) );
  XNOR U12662 ( .A(n11879), .B(n11878), .Z(n11864) );
  NANDN U12663 ( .A(n11849), .B(n11848), .Z(n11853) );
  OR U12664 ( .A(n11851), .B(n11850), .Z(n11852) );
  NAND U12665 ( .A(n11853), .B(n11852), .Z(n11865) );
  XNOR U12666 ( .A(n11864), .B(n11865), .Z(n11866) );
  XNOR U12667 ( .A(n11867), .B(n11866), .Z(n11859) );
  XOR U12668 ( .A(sreg[1484]), .B(n11859), .Z(n11860) );
  OR U12669 ( .A(n11854), .B(sreg[1483]), .Z(n11858) );
  NANDN U12670 ( .A(n11856), .B(n11855), .Z(n11857) );
  AND U12671 ( .A(n11858), .B(n11857), .Z(n11861) );
  XOR U12672 ( .A(n11860), .B(n11861), .Z(c[1484]) );
  OR U12673 ( .A(n11859), .B(sreg[1484]), .Z(n11863) );
  NANDN U12674 ( .A(n11861), .B(n11860), .Z(n11862) );
  AND U12675 ( .A(n11863), .B(n11862), .Z(n11883) );
  NANDN U12676 ( .A(n11865), .B(n11864), .Z(n11869) );
  NAND U12677 ( .A(n11867), .B(n11866), .Z(n11868) );
  NAND U12678 ( .A(n11869), .B(n11868), .Z(n11888) );
  AND U12679 ( .A(b[2]), .B(a[463]), .Z(n11894) );
  AND U12680 ( .A(a[464]), .B(b[1]), .Z(n11892) );
  AND U12681 ( .A(a[462]), .B(b[3]), .Z(n11891) );
  XOR U12682 ( .A(n11892), .B(n11891), .Z(n11893) );
  XOR U12683 ( .A(n11894), .B(n11893), .Z(n11897) );
  NAND U12684 ( .A(b[0]), .B(a[465]), .Z(n11898) );
  XOR U12685 ( .A(n11897), .B(n11898), .Z(n11900) );
  OR U12686 ( .A(n11871), .B(n11870), .Z(n11875) );
  NANDN U12687 ( .A(n11873), .B(n11872), .Z(n11874) );
  NAND U12688 ( .A(n11875), .B(n11874), .Z(n11899) );
  XNOR U12689 ( .A(n11900), .B(n11899), .Z(n11885) );
  NANDN U12690 ( .A(n11877), .B(n11876), .Z(n11881) );
  OR U12691 ( .A(n11879), .B(n11878), .Z(n11880) );
  NAND U12692 ( .A(n11881), .B(n11880), .Z(n11886) );
  XNOR U12693 ( .A(n11885), .B(n11886), .Z(n11887) );
  XNOR U12694 ( .A(n11888), .B(n11887), .Z(n11884) );
  XOR U12695 ( .A(sreg[1485]), .B(n11884), .Z(n11882) );
  XOR U12696 ( .A(n11883), .B(n11882), .Z(c[1485]) );
  NANDN U12697 ( .A(n11886), .B(n11885), .Z(n11890) );
  NAND U12698 ( .A(n11888), .B(n11887), .Z(n11889) );
  NAND U12699 ( .A(n11890), .B(n11889), .Z(n11906) );
  AND U12700 ( .A(b[2]), .B(a[464]), .Z(n11912) );
  AND U12701 ( .A(a[465]), .B(b[1]), .Z(n11910) );
  AND U12702 ( .A(a[463]), .B(b[3]), .Z(n11909) );
  XOR U12703 ( .A(n11910), .B(n11909), .Z(n11911) );
  XOR U12704 ( .A(n11912), .B(n11911), .Z(n11915) );
  NAND U12705 ( .A(b[0]), .B(a[466]), .Z(n11916) );
  XOR U12706 ( .A(n11915), .B(n11916), .Z(n11918) );
  OR U12707 ( .A(n11892), .B(n11891), .Z(n11896) );
  NANDN U12708 ( .A(n11894), .B(n11893), .Z(n11895) );
  NAND U12709 ( .A(n11896), .B(n11895), .Z(n11917) );
  XNOR U12710 ( .A(n11918), .B(n11917), .Z(n11903) );
  NANDN U12711 ( .A(n11898), .B(n11897), .Z(n11902) );
  OR U12712 ( .A(n11900), .B(n11899), .Z(n11901) );
  NAND U12713 ( .A(n11902), .B(n11901), .Z(n11904) );
  XNOR U12714 ( .A(n11903), .B(n11904), .Z(n11905) );
  XNOR U12715 ( .A(n11906), .B(n11905), .Z(n11921) );
  XOR U12716 ( .A(sreg[1486]), .B(n11921), .Z(n11922) );
  XOR U12717 ( .A(n11923), .B(n11922), .Z(c[1486]) );
  NANDN U12718 ( .A(n11904), .B(n11903), .Z(n11908) );
  NAND U12719 ( .A(n11906), .B(n11905), .Z(n11907) );
  NAND U12720 ( .A(n11908), .B(n11907), .Z(n11932) );
  AND U12721 ( .A(b[2]), .B(a[465]), .Z(n11938) );
  AND U12722 ( .A(a[466]), .B(b[1]), .Z(n11936) );
  AND U12723 ( .A(a[464]), .B(b[3]), .Z(n11935) );
  XOR U12724 ( .A(n11936), .B(n11935), .Z(n11937) );
  XOR U12725 ( .A(n11938), .B(n11937), .Z(n11941) );
  NAND U12726 ( .A(b[0]), .B(a[467]), .Z(n11942) );
  XOR U12727 ( .A(n11941), .B(n11942), .Z(n11944) );
  OR U12728 ( .A(n11910), .B(n11909), .Z(n11914) );
  NANDN U12729 ( .A(n11912), .B(n11911), .Z(n11913) );
  NAND U12730 ( .A(n11914), .B(n11913), .Z(n11943) );
  XNOR U12731 ( .A(n11944), .B(n11943), .Z(n11929) );
  NANDN U12732 ( .A(n11916), .B(n11915), .Z(n11920) );
  OR U12733 ( .A(n11918), .B(n11917), .Z(n11919) );
  NAND U12734 ( .A(n11920), .B(n11919), .Z(n11930) );
  XNOR U12735 ( .A(n11929), .B(n11930), .Z(n11931) );
  XOR U12736 ( .A(n11932), .B(n11931), .Z(n11928) );
  OR U12737 ( .A(n11921), .B(sreg[1486]), .Z(n11925) );
  NANDN U12738 ( .A(n11923), .B(n11922), .Z(n11924) );
  AND U12739 ( .A(n11925), .B(n11924), .Z(n11927) );
  XNOR U12740 ( .A(sreg[1487]), .B(n11927), .Z(n11926) );
  XOR U12741 ( .A(n11928), .B(n11926), .Z(c[1487]) );
  NANDN U12742 ( .A(n11930), .B(n11929), .Z(n11934) );
  NAND U12743 ( .A(n11932), .B(n11931), .Z(n11933) );
  NAND U12744 ( .A(n11934), .B(n11933), .Z(n11951) );
  AND U12745 ( .A(b[2]), .B(a[466]), .Z(n11957) );
  AND U12746 ( .A(a[467]), .B(b[1]), .Z(n11955) );
  AND U12747 ( .A(a[465]), .B(b[3]), .Z(n11954) );
  XOR U12748 ( .A(n11955), .B(n11954), .Z(n11956) );
  XOR U12749 ( .A(n11957), .B(n11956), .Z(n11960) );
  NAND U12750 ( .A(b[0]), .B(a[468]), .Z(n11961) );
  XOR U12751 ( .A(n11960), .B(n11961), .Z(n11963) );
  OR U12752 ( .A(n11936), .B(n11935), .Z(n11940) );
  NANDN U12753 ( .A(n11938), .B(n11937), .Z(n11939) );
  NAND U12754 ( .A(n11940), .B(n11939), .Z(n11962) );
  XNOR U12755 ( .A(n11963), .B(n11962), .Z(n11948) );
  NANDN U12756 ( .A(n11942), .B(n11941), .Z(n11946) );
  OR U12757 ( .A(n11944), .B(n11943), .Z(n11945) );
  NAND U12758 ( .A(n11946), .B(n11945), .Z(n11949) );
  XNOR U12759 ( .A(n11948), .B(n11949), .Z(n11950) );
  XNOR U12760 ( .A(n11951), .B(n11950), .Z(n11966) );
  XNOR U12761 ( .A(n11966), .B(sreg[1488]), .Z(n11947) );
  XOR U12762 ( .A(n11967), .B(n11947), .Z(c[1488]) );
  NANDN U12763 ( .A(n11949), .B(n11948), .Z(n11953) );
  NAND U12764 ( .A(n11951), .B(n11950), .Z(n11952) );
  NAND U12765 ( .A(n11953), .B(n11952), .Z(n11972) );
  AND U12766 ( .A(b[2]), .B(a[467]), .Z(n11978) );
  AND U12767 ( .A(a[468]), .B(b[1]), .Z(n11976) );
  AND U12768 ( .A(a[466]), .B(b[3]), .Z(n11975) );
  XOR U12769 ( .A(n11976), .B(n11975), .Z(n11977) );
  XOR U12770 ( .A(n11978), .B(n11977), .Z(n11981) );
  NAND U12771 ( .A(b[0]), .B(a[469]), .Z(n11982) );
  XOR U12772 ( .A(n11981), .B(n11982), .Z(n11984) );
  OR U12773 ( .A(n11955), .B(n11954), .Z(n11959) );
  NANDN U12774 ( .A(n11957), .B(n11956), .Z(n11958) );
  NAND U12775 ( .A(n11959), .B(n11958), .Z(n11983) );
  XNOR U12776 ( .A(n11984), .B(n11983), .Z(n11969) );
  NANDN U12777 ( .A(n11961), .B(n11960), .Z(n11965) );
  OR U12778 ( .A(n11963), .B(n11962), .Z(n11964) );
  NAND U12779 ( .A(n11965), .B(n11964), .Z(n11970) );
  XNOR U12780 ( .A(n11969), .B(n11970), .Z(n11971) );
  XNOR U12781 ( .A(n11972), .B(n11971), .Z(n11988) );
  XOR U12782 ( .A(n11987), .B(sreg[1489]), .Z(n11968) );
  XOR U12783 ( .A(n11988), .B(n11968), .Z(c[1489]) );
  NANDN U12784 ( .A(n11970), .B(n11969), .Z(n11974) );
  NAND U12785 ( .A(n11972), .B(n11971), .Z(n11973) );
  NAND U12786 ( .A(n11974), .B(n11973), .Z(n11993) );
  AND U12787 ( .A(b[2]), .B(a[468]), .Z(n11999) );
  AND U12788 ( .A(a[469]), .B(b[1]), .Z(n11997) );
  AND U12789 ( .A(a[467]), .B(b[3]), .Z(n11996) );
  XOR U12790 ( .A(n11997), .B(n11996), .Z(n11998) );
  XOR U12791 ( .A(n11999), .B(n11998), .Z(n12002) );
  NAND U12792 ( .A(b[0]), .B(a[470]), .Z(n12003) );
  XOR U12793 ( .A(n12002), .B(n12003), .Z(n12005) );
  OR U12794 ( .A(n11976), .B(n11975), .Z(n11980) );
  NANDN U12795 ( .A(n11978), .B(n11977), .Z(n11979) );
  NAND U12796 ( .A(n11980), .B(n11979), .Z(n12004) );
  XNOR U12797 ( .A(n12005), .B(n12004), .Z(n11990) );
  NANDN U12798 ( .A(n11982), .B(n11981), .Z(n11986) );
  OR U12799 ( .A(n11984), .B(n11983), .Z(n11985) );
  NAND U12800 ( .A(n11986), .B(n11985), .Z(n11991) );
  XNOR U12801 ( .A(n11990), .B(n11991), .Z(n11992) );
  XNOR U12802 ( .A(n11993), .B(n11992), .Z(n12009) );
  XOR U12803 ( .A(n12008), .B(sreg[1490]), .Z(n11989) );
  XOR U12804 ( .A(n12009), .B(n11989), .Z(c[1490]) );
  NANDN U12805 ( .A(n11991), .B(n11990), .Z(n11995) );
  NAND U12806 ( .A(n11993), .B(n11992), .Z(n11994) );
  NAND U12807 ( .A(n11995), .B(n11994), .Z(n12014) );
  AND U12808 ( .A(b[2]), .B(a[469]), .Z(n12020) );
  AND U12809 ( .A(a[470]), .B(b[1]), .Z(n12018) );
  AND U12810 ( .A(a[468]), .B(b[3]), .Z(n12017) );
  XOR U12811 ( .A(n12018), .B(n12017), .Z(n12019) );
  XOR U12812 ( .A(n12020), .B(n12019), .Z(n12023) );
  NAND U12813 ( .A(b[0]), .B(a[471]), .Z(n12024) );
  XOR U12814 ( .A(n12023), .B(n12024), .Z(n12026) );
  OR U12815 ( .A(n11997), .B(n11996), .Z(n12001) );
  NANDN U12816 ( .A(n11999), .B(n11998), .Z(n12000) );
  NAND U12817 ( .A(n12001), .B(n12000), .Z(n12025) );
  XNOR U12818 ( .A(n12026), .B(n12025), .Z(n12011) );
  NANDN U12819 ( .A(n12003), .B(n12002), .Z(n12007) );
  OR U12820 ( .A(n12005), .B(n12004), .Z(n12006) );
  NAND U12821 ( .A(n12007), .B(n12006), .Z(n12012) );
  XNOR U12822 ( .A(n12011), .B(n12012), .Z(n12013) );
  XOR U12823 ( .A(n12014), .B(n12013), .Z(n12030) );
  XOR U12824 ( .A(sreg[1491]), .B(n12029), .Z(n12010) );
  XOR U12825 ( .A(n12030), .B(n12010), .Z(c[1491]) );
  NANDN U12826 ( .A(n12012), .B(n12011), .Z(n12016) );
  NAND U12827 ( .A(n12014), .B(n12013), .Z(n12015) );
  NAND U12828 ( .A(n12016), .B(n12015), .Z(n12037) );
  AND U12829 ( .A(b[2]), .B(a[470]), .Z(n12043) );
  AND U12830 ( .A(a[471]), .B(b[1]), .Z(n12041) );
  AND U12831 ( .A(a[469]), .B(b[3]), .Z(n12040) );
  XOR U12832 ( .A(n12041), .B(n12040), .Z(n12042) );
  XOR U12833 ( .A(n12043), .B(n12042), .Z(n12046) );
  NAND U12834 ( .A(b[0]), .B(a[472]), .Z(n12047) );
  XOR U12835 ( .A(n12046), .B(n12047), .Z(n12049) );
  OR U12836 ( .A(n12018), .B(n12017), .Z(n12022) );
  NANDN U12837 ( .A(n12020), .B(n12019), .Z(n12021) );
  NAND U12838 ( .A(n12022), .B(n12021), .Z(n12048) );
  XNOR U12839 ( .A(n12049), .B(n12048), .Z(n12034) );
  NANDN U12840 ( .A(n12024), .B(n12023), .Z(n12028) );
  OR U12841 ( .A(n12026), .B(n12025), .Z(n12027) );
  NAND U12842 ( .A(n12028), .B(n12027), .Z(n12035) );
  XNOR U12843 ( .A(n12034), .B(n12035), .Z(n12036) );
  XOR U12844 ( .A(n12037), .B(n12036), .Z(n12033) );
  XNOR U12845 ( .A(sreg[1492]), .B(n12032), .Z(n12031) );
  XOR U12846 ( .A(n12033), .B(n12031), .Z(c[1492]) );
  NANDN U12847 ( .A(n12035), .B(n12034), .Z(n12039) );
  NAND U12848 ( .A(n12037), .B(n12036), .Z(n12038) );
  NAND U12849 ( .A(n12039), .B(n12038), .Z(n12055) );
  AND U12850 ( .A(b[2]), .B(a[471]), .Z(n12061) );
  AND U12851 ( .A(a[472]), .B(b[1]), .Z(n12059) );
  AND U12852 ( .A(a[470]), .B(b[3]), .Z(n12058) );
  XOR U12853 ( .A(n12059), .B(n12058), .Z(n12060) );
  XOR U12854 ( .A(n12061), .B(n12060), .Z(n12064) );
  NAND U12855 ( .A(b[0]), .B(a[473]), .Z(n12065) );
  XOR U12856 ( .A(n12064), .B(n12065), .Z(n12067) );
  OR U12857 ( .A(n12041), .B(n12040), .Z(n12045) );
  NANDN U12858 ( .A(n12043), .B(n12042), .Z(n12044) );
  NAND U12859 ( .A(n12045), .B(n12044), .Z(n12066) );
  XNOR U12860 ( .A(n12067), .B(n12066), .Z(n12052) );
  NANDN U12861 ( .A(n12047), .B(n12046), .Z(n12051) );
  OR U12862 ( .A(n12049), .B(n12048), .Z(n12050) );
  NAND U12863 ( .A(n12051), .B(n12050), .Z(n12053) );
  XNOR U12864 ( .A(n12052), .B(n12053), .Z(n12054) );
  XNOR U12865 ( .A(n12055), .B(n12054), .Z(n12070) );
  XNOR U12866 ( .A(n12070), .B(sreg[1493]), .Z(n12071) );
  XOR U12867 ( .A(n12072), .B(n12071), .Z(c[1493]) );
  NANDN U12868 ( .A(n12053), .B(n12052), .Z(n12057) );
  NAND U12869 ( .A(n12055), .B(n12054), .Z(n12056) );
  NAND U12870 ( .A(n12057), .B(n12056), .Z(n12078) );
  AND U12871 ( .A(b[2]), .B(a[472]), .Z(n12084) );
  AND U12872 ( .A(a[473]), .B(b[1]), .Z(n12082) );
  AND U12873 ( .A(a[471]), .B(b[3]), .Z(n12081) );
  XOR U12874 ( .A(n12082), .B(n12081), .Z(n12083) );
  XOR U12875 ( .A(n12084), .B(n12083), .Z(n12087) );
  NAND U12876 ( .A(b[0]), .B(a[474]), .Z(n12088) );
  XOR U12877 ( .A(n12087), .B(n12088), .Z(n12090) );
  OR U12878 ( .A(n12059), .B(n12058), .Z(n12063) );
  NANDN U12879 ( .A(n12061), .B(n12060), .Z(n12062) );
  NAND U12880 ( .A(n12063), .B(n12062), .Z(n12089) );
  XNOR U12881 ( .A(n12090), .B(n12089), .Z(n12075) );
  NANDN U12882 ( .A(n12065), .B(n12064), .Z(n12069) );
  OR U12883 ( .A(n12067), .B(n12066), .Z(n12068) );
  NAND U12884 ( .A(n12069), .B(n12068), .Z(n12076) );
  XNOR U12885 ( .A(n12075), .B(n12076), .Z(n12077) );
  XNOR U12886 ( .A(n12078), .B(n12077), .Z(n12093) );
  XOR U12887 ( .A(sreg[1494]), .B(n12093), .Z(n12094) );
  NAND U12888 ( .A(n12070), .B(sreg[1493]), .Z(n12074) );
  OR U12889 ( .A(n12072), .B(n12071), .Z(n12073) );
  NAND U12890 ( .A(n12074), .B(n12073), .Z(n12095) );
  XOR U12891 ( .A(n12094), .B(n12095), .Z(c[1494]) );
  NANDN U12892 ( .A(n12076), .B(n12075), .Z(n12080) );
  NAND U12893 ( .A(n12078), .B(n12077), .Z(n12079) );
  NAND U12894 ( .A(n12080), .B(n12079), .Z(n12102) );
  AND U12895 ( .A(b[2]), .B(a[473]), .Z(n12108) );
  AND U12896 ( .A(a[474]), .B(b[1]), .Z(n12106) );
  AND U12897 ( .A(a[472]), .B(b[3]), .Z(n12105) );
  XOR U12898 ( .A(n12106), .B(n12105), .Z(n12107) );
  XOR U12899 ( .A(n12108), .B(n12107), .Z(n12111) );
  NAND U12900 ( .A(b[0]), .B(a[475]), .Z(n12112) );
  XOR U12901 ( .A(n12111), .B(n12112), .Z(n12114) );
  OR U12902 ( .A(n12082), .B(n12081), .Z(n12086) );
  NANDN U12903 ( .A(n12084), .B(n12083), .Z(n12085) );
  NAND U12904 ( .A(n12086), .B(n12085), .Z(n12113) );
  XNOR U12905 ( .A(n12114), .B(n12113), .Z(n12099) );
  NANDN U12906 ( .A(n12088), .B(n12087), .Z(n12092) );
  OR U12907 ( .A(n12090), .B(n12089), .Z(n12091) );
  NAND U12908 ( .A(n12092), .B(n12091), .Z(n12100) );
  XNOR U12909 ( .A(n12099), .B(n12100), .Z(n12101) );
  XOR U12910 ( .A(n12102), .B(n12101), .Z(n12118) );
  OR U12911 ( .A(n12093), .B(sreg[1494]), .Z(n12097) );
  NANDN U12912 ( .A(n12095), .B(n12094), .Z(n12096) );
  AND U12913 ( .A(n12097), .B(n12096), .Z(n12117) );
  XNOR U12914 ( .A(sreg[1495]), .B(n12117), .Z(n12098) );
  XOR U12915 ( .A(n12118), .B(n12098), .Z(c[1495]) );
  NANDN U12916 ( .A(n12100), .B(n12099), .Z(n12104) );
  NAND U12917 ( .A(n12102), .B(n12101), .Z(n12103) );
  NAND U12918 ( .A(n12104), .B(n12103), .Z(n12123) );
  AND U12919 ( .A(b[2]), .B(a[474]), .Z(n12129) );
  AND U12920 ( .A(a[475]), .B(b[1]), .Z(n12127) );
  AND U12921 ( .A(a[473]), .B(b[3]), .Z(n12126) );
  XOR U12922 ( .A(n12127), .B(n12126), .Z(n12128) );
  XOR U12923 ( .A(n12129), .B(n12128), .Z(n12132) );
  NAND U12924 ( .A(b[0]), .B(a[476]), .Z(n12133) );
  XOR U12925 ( .A(n12132), .B(n12133), .Z(n12135) );
  OR U12926 ( .A(n12106), .B(n12105), .Z(n12110) );
  NANDN U12927 ( .A(n12108), .B(n12107), .Z(n12109) );
  NAND U12928 ( .A(n12110), .B(n12109), .Z(n12134) );
  XNOR U12929 ( .A(n12135), .B(n12134), .Z(n12120) );
  NANDN U12930 ( .A(n12112), .B(n12111), .Z(n12116) );
  OR U12931 ( .A(n12114), .B(n12113), .Z(n12115) );
  NAND U12932 ( .A(n12116), .B(n12115), .Z(n12121) );
  XNOR U12933 ( .A(n12120), .B(n12121), .Z(n12122) );
  XOR U12934 ( .A(n12123), .B(n12122), .Z(n12139) );
  XNOR U12935 ( .A(sreg[1496]), .B(n12138), .Z(n12119) );
  XOR U12936 ( .A(n12139), .B(n12119), .Z(c[1496]) );
  NANDN U12937 ( .A(n12121), .B(n12120), .Z(n12125) );
  NAND U12938 ( .A(n12123), .B(n12122), .Z(n12124) );
  NAND U12939 ( .A(n12125), .B(n12124), .Z(n12146) );
  AND U12940 ( .A(b[2]), .B(a[475]), .Z(n12152) );
  AND U12941 ( .A(a[476]), .B(b[1]), .Z(n12150) );
  AND U12942 ( .A(a[474]), .B(b[3]), .Z(n12149) );
  XOR U12943 ( .A(n12150), .B(n12149), .Z(n12151) );
  XOR U12944 ( .A(n12152), .B(n12151), .Z(n12155) );
  NAND U12945 ( .A(b[0]), .B(a[477]), .Z(n12156) );
  XOR U12946 ( .A(n12155), .B(n12156), .Z(n12158) );
  OR U12947 ( .A(n12127), .B(n12126), .Z(n12131) );
  NANDN U12948 ( .A(n12129), .B(n12128), .Z(n12130) );
  NAND U12949 ( .A(n12131), .B(n12130), .Z(n12157) );
  XNOR U12950 ( .A(n12158), .B(n12157), .Z(n12143) );
  NANDN U12951 ( .A(n12133), .B(n12132), .Z(n12137) );
  OR U12952 ( .A(n12135), .B(n12134), .Z(n12136) );
  NAND U12953 ( .A(n12137), .B(n12136), .Z(n12144) );
  XNOR U12954 ( .A(n12143), .B(n12144), .Z(n12145) );
  XNOR U12955 ( .A(n12146), .B(n12145), .Z(n12142) );
  XOR U12956 ( .A(n12141), .B(sreg[1497]), .Z(n12140) );
  XOR U12957 ( .A(n12142), .B(n12140), .Z(c[1497]) );
  NANDN U12958 ( .A(n12144), .B(n12143), .Z(n12148) );
  NAND U12959 ( .A(n12146), .B(n12145), .Z(n12147) );
  NAND U12960 ( .A(n12148), .B(n12147), .Z(n12169) );
  AND U12961 ( .A(b[2]), .B(a[476]), .Z(n12175) );
  AND U12962 ( .A(a[477]), .B(b[1]), .Z(n12173) );
  AND U12963 ( .A(a[475]), .B(b[3]), .Z(n12172) );
  XOR U12964 ( .A(n12173), .B(n12172), .Z(n12174) );
  XOR U12965 ( .A(n12175), .B(n12174), .Z(n12178) );
  NAND U12966 ( .A(b[0]), .B(a[478]), .Z(n12179) );
  XOR U12967 ( .A(n12178), .B(n12179), .Z(n12181) );
  OR U12968 ( .A(n12150), .B(n12149), .Z(n12154) );
  NANDN U12969 ( .A(n12152), .B(n12151), .Z(n12153) );
  NAND U12970 ( .A(n12154), .B(n12153), .Z(n12180) );
  XNOR U12971 ( .A(n12181), .B(n12180), .Z(n12166) );
  NANDN U12972 ( .A(n12156), .B(n12155), .Z(n12160) );
  OR U12973 ( .A(n12158), .B(n12157), .Z(n12159) );
  NAND U12974 ( .A(n12160), .B(n12159), .Z(n12167) );
  XNOR U12975 ( .A(n12166), .B(n12167), .Z(n12168) );
  XNOR U12976 ( .A(n12169), .B(n12168), .Z(n12161) );
  XOR U12977 ( .A(sreg[1498]), .B(n12161), .Z(n12162) );
  XOR U12978 ( .A(n12163), .B(n12162), .Z(c[1498]) );
  OR U12979 ( .A(n12161), .B(sreg[1498]), .Z(n12165) );
  NANDN U12980 ( .A(n12163), .B(n12162), .Z(n12164) );
  NAND U12981 ( .A(n12165), .B(n12164), .Z(n12204) );
  NANDN U12982 ( .A(n12167), .B(n12166), .Z(n12171) );
  NAND U12983 ( .A(n12169), .B(n12168), .Z(n12170) );
  NAND U12984 ( .A(n12171), .B(n12170), .Z(n12187) );
  AND U12985 ( .A(b[2]), .B(a[477]), .Z(n12193) );
  AND U12986 ( .A(a[478]), .B(b[1]), .Z(n12191) );
  AND U12987 ( .A(a[476]), .B(b[3]), .Z(n12190) );
  XOR U12988 ( .A(n12191), .B(n12190), .Z(n12192) );
  XOR U12989 ( .A(n12193), .B(n12192), .Z(n12196) );
  NAND U12990 ( .A(b[0]), .B(a[479]), .Z(n12197) );
  XOR U12991 ( .A(n12196), .B(n12197), .Z(n12199) );
  OR U12992 ( .A(n12173), .B(n12172), .Z(n12177) );
  NANDN U12993 ( .A(n12175), .B(n12174), .Z(n12176) );
  NAND U12994 ( .A(n12177), .B(n12176), .Z(n12198) );
  XNOR U12995 ( .A(n12199), .B(n12198), .Z(n12184) );
  NANDN U12996 ( .A(n12179), .B(n12178), .Z(n12183) );
  OR U12997 ( .A(n12181), .B(n12180), .Z(n12182) );
  NAND U12998 ( .A(n12183), .B(n12182), .Z(n12185) );
  XNOR U12999 ( .A(n12184), .B(n12185), .Z(n12186) );
  XNOR U13000 ( .A(n12187), .B(n12186), .Z(n12202) );
  XNOR U13001 ( .A(n12202), .B(sreg[1499]), .Z(n12203) );
  XOR U13002 ( .A(n12204), .B(n12203), .Z(c[1499]) );
  NANDN U13003 ( .A(n12185), .B(n12184), .Z(n12189) );
  NAND U13004 ( .A(n12187), .B(n12186), .Z(n12188) );
  NAND U13005 ( .A(n12189), .B(n12188), .Z(n12211) );
  AND U13006 ( .A(b[2]), .B(a[478]), .Z(n12223) );
  AND U13007 ( .A(a[479]), .B(b[1]), .Z(n12221) );
  AND U13008 ( .A(a[477]), .B(b[3]), .Z(n12220) );
  XOR U13009 ( .A(n12221), .B(n12220), .Z(n12222) );
  XOR U13010 ( .A(n12223), .B(n12222), .Z(n12214) );
  NAND U13011 ( .A(b[0]), .B(a[480]), .Z(n12215) );
  XOR U13012 ( .A(n12214), .B(n12215), .Z(n12217) );
  OR U13013 ( .A(n12191), .B(n12190), .Z(n12195) );
  NANDN U13014 ( .A(n12193), .B(n12192), .Z(n12194) );
  NAND U13015 ( .A(n12195), .B(n12194), .Z(n12216) );
  XNOR U13016 ( .A(n12217), .B(n12216), .Z(n12208) );
  NANDN U13017 ( .A(n12197), .B(n12196), .Z(n12201) );
  OR U13018 ( .A(n12199), .B(n12198), .Z(n12200) );
  NAND U13019 ( .A(n12201), .B(n12200), .Z(n12209) );
  XNOR U13020 ( .A(n12208), .B(n12209), .Z(n12210) );
  XOR U13021 ( .A(n12211), .B(n12210), .Z(n12228) );
  NAND U13022 ( .A(n12202), .B(sreg[1499]), .Z(n12206) );
  OR U13023 ( .A(n12204), .B(n12203), .Z(n12205) );
  NAND U13024 ( .A(n12206), .B(n12205), .Z(n12227) );
  XNOR U13025 ( .A(sreg[1500]), .B(n12227), .Z(n12207) );
  XOR U13026 ( .A(n12228), .B(n12207), .Z(c[1500]) );
  NANDN U13027 ( .A(n12209), .B(n12208), .Z(n12213) );
  NAND U13028 ( .A(n12211), .B(n12210), .Z(n12212) );
  NAND U13029 ( .A(n12213), .B(n12212), .Z(n12232) );
  NANDN U13030 ( .A(n12215), .B(n12214), .Z(n12219) );
  OR U13031 ( .A(n12217), .B(n12216), .Z(n12218) );
  AND U13032 ( .A(n12219), .B(n12218), .Z(n12231) );
  AND U13033 ( .A(b[2]), .B(a[479]), .Z(n12236) );
  AND U13034 ( .A(a[480]), .B(b[1]), .Z(n12234) );
  AND U13035 ( .A(a[478]), .B(b[3]), .Z(n12233) );
  XOR U13036 ( .A(n12234), .B(n12233), .Z(n12235) );
  XOR U13037 ( .A(n12236), .B(n12235), .Z(n12239) );
  NAND U13038 ( .A(b[0]), .B(a[481]), .Z(n12240) );
  XOR U13039 ( .A(n12239), .B(n12240), .Z(n12242) );
  OR U13040 ( .A(n12221), .B(n12220), .Z(n12225) );
  NANDN U13041 ( .A(n12223), .B(n12222), .Z(n12224) );
  NAND U13042 ( .A(n12225), .B(n12224), .Z(n12241) );
  XOR U13043 ( .A(n12242), .B(n12241), .Z(n12230) );
  XNOR U13044 ( .A(n12231), .B(n12230), .Z(n12226) );
  XNOR U13045 ( .A(n12232), .B(n12226), .Z(n12246) );
  XOR U13046 ( .A(n12245), .B(sreg[1501]), .Z(n12229) );
  XOR U13047 ( .A(n12246), .B(n12229), .Z(c[1501]) );
  AND U13048 ( .A(b[2]), .B(a[480]), .Z(n12259) );
  AND U13049 ( .A(a[481]), .B(b[1]), .Z(n12257) );
  AND U13050 ( .A(a[479]), .B(b[3]), .Z(n12256) );
  XOR U13051 ( .A(n12257), .B(n12256), .Z(n12258) );
  XOR U13052 ( .A(n12259), .B(n12258), .Z(n12262) );
  NAND U13053 ( .A(b[0]), .B(a[482]), .Z(n12263) );
  XOR U13054 ( .A(n12262), .B(n12263), .Z(n12265) );
  OR U13055 ( .A(n12234), .B(n12233), .Z(n12238) );
  NANDN U13056 ( .A(n12236), .B(n12235), .Z(n12237) );
  NAND U13057 ( .A(n12238), .B(n12237), .Z(n12264) );
  XNOR U13058 ( .A(n12265), .B(n12264), .Z(n12250) );
  NANDN U13059 ( .A(n12240), .B(n12239), .Z(n12244) );
  OR U13060 ( .A(n12242), .B(n12241), .Z(n12243) );
  NAND U13061 ( .A(n12244), .B(n12243), .Z(n12251) );
  XNOR U13062 ( .A(n12250), .B(n12251), .Z(n12252) );
  XOR U13063 ( .A(n12253), .B(n12252), .Z(n12249) );
  XOR U13064 ( .A(sreg[1502]), .B(n12248), .Z(n12247) );
  XNOR U13065 ( .A(n12249), .B(n12247), .Z(c[1502]) );
  NANDN U13066 ( .A(n12251), .B(n12250), .Z(n12255) );
  NANDN U13067 ( .A(n12253), .B(n12252), .Z(n12254) );
  NAND U13068 ( .A(n12255), .B(n12254), .Z(n12276) );
  AND U13069 ( .A(b[2]), .B(a[481]), .Z(n12282) );
  AND U13070 ( .A(a[482]), .B(b[1]), .Z(n12280) );
  AND U13071 ( .A(a[480]), .B(b[3]), .Z(n12279) );
  XOR U13072 ( .A(n12280), .B(n12279), .Z(n12281) );
  XOR U13073 ( .A(n12282), .B(n12281), .Z(n12285) );
  NAND U13074 ( .A(b[0]), .B(a[483]), .Z(n12286) );
  XOR U13075 ( .A(n12285), .B(n12286), .Z(n12288) );
  OR U13076 ( .A(n12257), .B(n12256), .Z(n12261) );
  NANDN U13077 ( .A(n12259), .B(n12258), .Z(n12260) );
  NAND U13078 ( .A(n12261), .B(n12260), .Z(n12287) );
  XNOR U13079 ( .A(n12288), .B(n12287), .Z(n12273) );
  NANDN U13080 ( .A(n12263), .B(n12262), .Z(n12267) );
  OR U13081 ( .A(n12265), .B(n12264), .Z(n12266) );
  NAND U13082 ( .A(n12267), .B(n12266), .Z(n12274) );
  XNOR U13083 ( .A(n12273), .B(n12274), .Z(n12275) );
  XNOR U13084 ( .A(n12276), .B(n12275), .Z(n12268) );
  XNOR U13085 ( .A(n12268), .B(sreg[1503]), .Z(n12269) );
  XOR U13086 ( .A(n12270), .B(n12269), .Z(c[1503]) );
  NAND U13087 ( .A(n12268), .B(sreg[1503]), .Z(n12272) );
  OR U13088 ( .A(n12270), .B(n12269), .Z(n12271) );
  AND U13089 ( .A(n12272), .B(n12271), .Z(n12307) );
  NANDN U13090 ( .A(n12274), .B(n12273), .Z(n12278) );
  NAND U13091 ( .A(n12276), .B(n12275), .Z(n12277) );
  AND U13092 ( .A(n12278), .B(n12277), .Z(n12295) );
  AND U13093 ( .A(b[2]), .B(a[482]), .Z(n12299) );
  AND U13094 ( .A(a[483]), .B(b[1]), .Z(n12297) );
  AND U13095 ( .A(a[481]), .B(b[3]), .Z(n12296) );
  XOR U13096 ( .A(n12297), .B(n12296), .Z(n12298) );
  XOR U13097 ( .A(n12299), .B(n12298), .Z(n12302) );
  NAND U13098 ( .A(b[0]), .B(a[484]), .Z(n12303) );
  XOR U13099 ( .A(n12302), .B(n12303), .Z(n12304) );
  OR U13100 ( .A(n12280), .B(n12279), .Z(n12284) );
  NANDN U13101 ( .A(n12282), .B(n12281), .Z(n12283) );
  AND U13102 ( .A(n12284), .B(n12283), .Z(n12305) );
  XOR U13103 ( .A(n12304), .B(n12305), .Z(n12293) );
  NANDN U13104 ( .A(n12286), .B(n12285), .Z(n12290) );
  OR U13105 ( .A(n12288), .B(n12287), .Z(n12289) );
  AND U13106 ( .A(n12290), .B(n12289), .Z(n12294) );
  XOR U13107 ( .A(n12293), .B(n12294), .Z(n12291) );
  XOR U13108 ( .A(n12295), .B(n12291), .Z(n12306) );
  XNOR U13109 ( .A(sreg[1504]), .B(n12306), .Z(n12292) );
  XOR U13110 ( .A(n12307), .B(n12292), .Z(c[1504]) );
  AND U13111 ( .A(b[2]), .B(a[483]), .Z(n12320) );
  AND U13112 ( .A(a[484]), .B(b[1]), .Z(n12318) );
  AND U13113 ( .A(a[482]), .B(b[3]), .Z(n12317) );
  XOR U13114 ( .A(n12318), .B(n12317), .Z(n12319) );
  XOR U13115 ( .A(n12320), .B(n12319), .Z(n12323) );
  NAND U13116 ( .A(b[0]), .B(a[485]), .Z(n12324) );
  XOR U13117 ( .A(n12323), .B(n12324), .Z(n12326) );
  OR U13118 ( .A(n12297), .B(n12296), .Z(n12301) );
  NANDN U13119 ( .A(n12299), .B(n12298), .Z(n12300) );
  NAND U13120 ( .A(n12301), .B(n12300), .Z(n12325) );
  XNOR U13121 ( .A(n12326), .B(n12325), .Z(n12311) );
  XNOR U13122 ( .A(n12311), .B(n12312), .Z(n12314) );
  XOR U13123 ( .A(n12313), .B(n12314), .Z(n12310) );
  XNOR U13124 ( .A(sreg[1505]), .B(n12309), .Z(n12308) );
  XOR U13125 ( .A(n12310), .B(n12308), .Z(c[1505]) );
  NANDN U13126 ( .A(n12312), .B(n12311), .Z(n12316) );
  NAND U13127 ( .A(n12314), .B(n12313), .Z(n12315) );
  NAND U13128 ( .A(n12316), .B(n12315), .Z(n12332) );
  AND U13129 ( .A(b[2]), .B(a[484]), .Z(n12338) );
  AND U13130 ( .A(a[485]), .B(b[1]), .Z(n12336) );
  AND U13131 ( .A(a[483]), .B(b[3]), .Z(n12335) );
  XOR U13132 ( .A(n12336), .B(n12335), .Z(n12337) );
  XOR U13133 ( .A(n12338), .B(n12337), .Z(n12341) );
  NAND U13134 ( .A(b[0]), .B(a[486]), .Z(n12342) );
  XOR U13135 ( .A(n12341), .B(n12342), .Z(n12344) );
  OR U13136 ( .A(n12318), .B(n12317), .Z(n12322) );
  NANDN U13137 ( .A(n12320), .B(n12319), .Z(n12321) );
  NAND U13138 ( .A(n12322), .B(n12321), .Z(n12343) );
  XNOR U13139 ( .A(n12344), .B(n12343), .Z(n12329) );
  NANDN U13140 ( .A(n12324), .B(n12323), .Z(n12328) );
  OR U13141 ( .A(n12326), .B(n12325), .Z(n12327) );
  NAND U13142 ( .A(n12328), .B(n12327), .Z(n12330) );
  XNOR U13143 ( .A(n12329), .B(n12330), .Z(n12331) );
  XNOR U13144 ( .A(n12332), .B(n12331), .Z(n12347) );
  XNOR U13145 ( .A(n12347), .B(sreg[1506]), .Z(n12348) );
  XOR U13146 ( .A(n12349), .B(n12348), .Z(c[1506]) );
  NANDN U13147 ( .A(n12330), .B(n12329), .Z(n12334) );
  NAND U13148 ( .A(n12332), .B(n12331), .Z(n12333) );
  NAND U13149 ( .A(n12334), .B(n12333), .Z(n12360) );
  AND U13150 ( .A(b[2]), .B(a[485]), .Z(n12366) );
  AND U13151 ( .A(a[486]), .B(b[1]), .Z(n12364) );
  AND U13152 ( .A(a[484]), .B(b[3]), .Z(n12363) );
  XOR U13153 ( .A(n12364), .B(n12363), .Z(n12365) );
  XOR U13154 ( .A(n12366), .B(n12365), .Z(n12369) );
  NAND U13155 ( .A(b[0]), .B(a[487]), .Z(n12370) );
  XOR U13156 ( .A(n12369), .B(n12370), .Z(n12372) );
  OR U13157 ( .A(n12336), .B(n12335), .Z(n12340) );
  NANDN U13158 ( .A(n12338), .B(n12337), .Z(n12339) );
  NAND U13159 ( .A(n12340), .B(n12339), .Z(n12371) );
  XNOR U13160 ( .A(n12372), .B(n12371), .Z(n12357) );
  NANDN U13161 ( .A(n12342), .B(n12341), .Z(n12346) );
  OR U13162 ( .A(n12344), .B(n12343), .Z(n12345) );
  NAND U13163 ( .A(n12346), .B(n12345), .Z(n12358) );
  XNOR U13164 ( .A(n12357), .B(n12358), .Z(n12359) );
  XNOR U13165 ( .A(n12360), .B(n12359), .Z(n12352) );
  XOR U13166 ( .A(sreg[1507]), .B(n12352), .Z(n12353) );
  NAND U13167 ( .A(n12347), .B(sreg[1506]), .Z(n12351) );
  OR U13168 ( .A(n12349), .B(n12348), .Z(n12350) );
  NAND U13169 ( .A(n12351), .B(n12350), .Z(n12354) );
  XOR U13170 ( .A(n12353), .B(n12354), .Z(c[1507]) );
  OR U13171 ( .A(n12352), .B(sreg[1507]), .Z(n12356) );
  NANDN U13172 ( .A(n12354), .B(n12353), .Z(n12355) );
  AND U13173 ( .A(n12356), .B(n12355), .Z(n12376) );
  NANDN U13174 ( .A(n12358), .B(n12357), .Z(n12362) );
  NAND U13175 ( .A(n12360), .B(n12359), .Z(n12361) );
  NAND U13176 ( .A(n12362), .B(n12361), .Z(n12381) );
  AND U13177 ( .A(b[2]), .B(a[486]), .Z(n12387) );
  AND U13178 ( .A(a[487]), .B(b[1]), .Z(n12385) );
  AND U13179 ( .A(a[485]), .B(b[3]), .Z(n12384) );
  XOR U13180 ( .A(n12385), .B(n12384), .Z(n12386) );
  XOR U13181 ( .A(n12387), .B(n12386), .Z(n12390) );
  NAND U13182 ( .A(b[0]), .B(a[488]), .Z(n12391) );
  XOR U13183 ( .A(n12390), .B(n12391), .Z(n12393) );
  OR U13184 ( .A(n12364), .B(n12363), .Z(n12368) );
  NANDN U13185 ( .A(n12366), .B(n12365), .Z(n12367) );
  NAND U13186 ( .A(n12368), .B(n12367), .Z(n12392) );
  XNOR U13187 ( .A(n12393), .B(n12392), .Z(n12378) );
  NANDN U13188 ( .A(n12370), .B(n12369), .Z(n12374) );
  OR U13189 ( .A(n12372), .B(n12371), .Z(n12373) );
  NAND U13190 ( .A(n12374), .B(n12373), .Z(n12379) );
  XNOR U13191 ( .A(n12378), .B(n12379), .Z(n12380) );
  XNOR U13192 ( .A(n12381), .B(n12380), .Z(n12377) );
  XOR U13193 ( .A(sreg[1508]), .B(n12377), .Z(n12375) );
  XOR U13194 ( .A(n12376), .B(n12375), .Z(c[1508]) );
  NANDN U13195 ( .A(n12379), .B(n12378), .Z(n12383) );
  NAND U13196 ( .A(n12381), .B(n12380), .Z(n12382) );
  NAND U13197 ( .A(n12383), .B(n12382), .Z(n12399) );
  AND U13198 ( .A(b[2]), .B(a[487]), .Z(n12405) );
  AND U13199 ( .A(a[488]), .B(b[1]), .Z(n12403) );
  AND U13200 ( .A(a[486]), .B(b[3]), .Z(n12402) );
  XOR U13201 ( .A(n12403), .B(n12402), .Z(n12404) );
  XOR U13202 ( .A(n12405), .B(n12404), .Z(n12408) );
  NAND U13203 ( .A(b[0]), .B(a[489]), .Z(n12409) );
  XOR U13204 ( .A(n12408), .B(n12409), .Z(n12411) );
  OR U13205 ( .A(n12385), .B(n12384), .Z(n12389) );
  NANDN U13206 ( .A(n12387), .B(n12386), .Z(n12388) );
  NAND U13207 ( .A(n12389), .B(n12388), .Z(n12410) );
  XNOR U13208 ( .A(n12411), .B(n12410), .Z(n12396) );
  NANDN U13209 ( .A(n12391), .B(n12390), .Z(n12395) );
  OR U13210 ( .A(n12393), .B(n12392), .Z(n12394) );
  NAND U13211 ( .A(n12395), .B(n12394), .Z(n12397) );
  XNOR U13212 ( .A(n12396), .B(n12397), .Z(n12398) );
  XOR U13213 ( .A(n12399), .B(n12398), .Z(n12414) );
  XOR U13214 ( .A(sreg[1509]), .B(n12414), .Z(n12416) );
  XNOR U13215 ( .A(n12415), .B(n12416), .Z(c[1509]) );
  NANDN U13216 ( .A(n12397), .B(n12396), .Z(n12401) );
  NAND U13217 ( .A(n12399), .B(n12398), .Z(n12400) );
  NAND U13218 ( .A(n12401), .B(n12400), .Z(n12422) );
  AND U13219 ( .A(b[2]), .B(a[488]), .Z(n12428) );
  AND U13220 ( .A(a[489]), .B(b[1]), .Z(n12426) );
  AND U13221 ( .A(a[487]), .B(b[3]), .Z(n12425) );
  XOR U13222 ( .A(n12426), .B(n12425), .Z(n12427) );
  XOR U13223 ( .A(n12428), .B(n12427), .Z(n12431) );
  NAND U13224 ( .A(b[0]), .B(a[490]), .Z(n12432) );
  XOR U13225 ( .A(n12431), .B(n12432), .Z(n12434) );
  OR U13226 ( .A(n12403), .B(n12402), .Z(n12407) );
  NANDN U13227 ( .A(n12405), .B(n12404), .Z(n12406) );
  NAND U13228 ( .A(n12407), .B(n12406), .Z(n12433) );
  XNOR U13229 ( .A(n12434), .B(n12433), .Z(n12419) );
  NANDN U13230 ( .A(n12409), .B(n12408), .Z(n12413) );
  OR U13231 ( .A(n12411), .B(n12410), .Z(n12412) );
  NAND U13232 ( .A(n12413), .B(n12412), .Z(n12420) );
  XNOR U13233 ( .A(n12419), .B(n12420), .Z(n12421) );
  XNOR U13234 ( .A(n12422), .B(n12421), .Z(n12437) );
  XOR U13235 ( .A(sreg[1510]), .B(n12437), .Z(n12438) );
  NANDN U13236 ( .A(n12414), .B(sreg[1509]), .Z(n12418) );
  NANDN U13237 ( .A(n12416), .B(n12415), .Z(n12417) );
  NAND U13238 ( .A(n12418), .B(n12417), .Z(n12439) );
  XOR U13239 ( .A(n12438), .B(n12439), .Z(c[1510]) );
  NANDN U13240 ( .A(n12420), .B(n12419), .Z(n12424) );
  NAND U13241 ( .A(n12422), .B(n12421), .Z(n12423) );
  NAND U13242 ( .A(n12424), .B(n12423), .Z(n12446) );
  AND U13243 ( .A(b[2]), .B(a[489]), .Z(n12452) );
  AND U13244 ( .A(a[490]), .B(b[1]), .Z(n12450) );
  AND U13245 ( .A(a[488]), .B(b[3]), .Z(n12449) );
  XOR U13246 ( .A(n12450), .B(n12449), .Z(n12451) );
  XOR U13247 ( .A(n12452), .B(n12451), .Z(n12455) );
  NAND U13248 ( .A(b[0]), .B(a[491]), .Z(n12456) );
  XOR U13249 ( .A(n12455), .B(n12456), .Z(n12458) );
  OR U13250 ( .A(n12426), .B(n12425), .Z(n12430) );
  NANDN U13251 ( .A(n12428), .B(n12427), .Z(n12429) );
  NAND U13252 ( .A(n12430), .B(n12429), .Z(n12457) );
  XNOR U13253 ( .A(n12458), .B(n12457), .Z(n12443) );
  NANDN U13254 ( .A(n12432), .B(n12431), .Z(n12436) );
  OR U13255 ( .A(n12434), .B(n12433), .Z(n12435) );
  NAND U13256 ( .A(n12436), .B(n12435), .Z(n12444) );
  XNOR U13257 ( .A(n12443), .B(n12444), .Z(n12445) );
  XOR U13258 ( .A(n12446), .B(n12445), .Z(n12462) );
  OR U13259 ( .A(n12437), .B(sreg[1510]), .Z(n12441) );
  NANDN U13260 ( .A(n12439), .B(n12438), .Z(n12440) );
  AND U13261 ( .A(n12441), .B(n12440), .Z(n12461) );
  XNOR U13262 ( .A(sreg[1511]), .B(n12461), .Z(n12442) );
  XOR U13263 ( .A(n12462), .B(n12442), .Z(c[1511]) );
  NANDN U13264 ( .A(n12444), .B(n12443), .Z(n12448) );
  NAND U13265 ( .A(n12446), .B(n12445), .Z(n12447) );
  NAND U13266 ( .A(n12448), .B(n12447), .Z(n12469) );
  AND U13267 ( .A(b[2]), .B(a[490]), .Z(n12475) );
  AND U13268 ( .A(a[491]), .B(b[1]), .Z(n12473) );
  AND U13269 ( .A(a[489]), .B(b[3]), .Z(n12472) );
  XOR U13270 ( .A(n12473), .B(n12472), .Z(n12474) );
  XOR U13271 ( .A(n12475), .B(n12474), .Z(n12478) );
  NAND U13272 ( .A(b[0]), .B(a[492]), .Z(n12479) );
  XOR U13273 ( .A(n12478), .B(n12479), .Z(n12481) );
  OR U13274 ( .A(n12450), .B(n12449), .Z(n12454) );
  NANDN U13275 ( .A(n12452), .B(n12451), .Z(n12453) );
  NAND U13276 ( .A(n12454), .B(n12453), .Z(n12480) );
  XNOR U13277 ( .A(n12481), .B(n12480), .Z(n12466) );
  NANDN U13278 ( .A(n12456), .B(n12455), .Z(n12460) );
  OR U13279 ( .A(n12458), .B(n12457), .Z(n12459) );
  NAND U13280 ( .A(n12460), .B(n12459), .Z(n12467) );
  XNOR U13281 ( .A(n12466), .B(n12467), .Z(n12468) );
  XNOR U13282 ( .A(n12469), .B(n12468), .Z(n12465) );
  XOR U13283 ( .A(n12464), .B(sreg[1512]), .Z(n12463) );
  XOR U13284 ( .A(n12465), .B(n12463), .Z(c[1512]) );
  NANDN U13285 ( .A(n12467), .B(n12466), .Z(n12471) );
  NAND U13286 ( .A(n12469), .B(n12468), .Z(n12470) );
  NAND U13287 ( .A(n12471), .B(n12470), .Z(n12487) );
  AND U13288 ( .A(b[2]), .B(a[491]), .Z(n12493) );
  AND U13289 ( .A(a[492]), .B(b[1]), .Z(n12491) );
  AND U13290 ( .A(a[490]), .B(b[3]), .Z(n12490) );
  XOR U13291 ( .A(n12491), .B(n12490), .Z(n12492) );
  XOR U13292 ( .A(n12493), .B(n12492), .Z(n12496) );
  NAND U13293 ( .A(b[0]), .B(a[493]), .Z(n12497) );
  XOR U13294 ( .A(n12496), .B(n12497), .Z(n12499) );
  OR U13295 ( .A(n12473), .B(n12472), .Z(n12477) );
  NANDN U13296 ( .A(n12475), .B(n12474), .Z(n12476) );
  NAND U13297 ( .A(n12477), .B(n12476), .Z(n12498) );
  XNOR U13298 ( .A(n12499), .B(n12498), .Z(n12484) );
  NANDN U13299 ( .A(n12479), .B(n12478), .Z(n12483) );
  OR U13300 ( .A(n12481), .B(n12480), .Z(n12482) );
  NAND U13301 ( .A(n12483), .B(n12482), .Z(n12485) );
  XNOR U13302 ( .A(n12484), .B(n12485), .Z(n12486) );
  XNOR U13303 ( .A(n12487), .B(n12486), .Z(n12502) );
  XNOR U13304 ( .A(n12502), .B(sreg[1513]), .Z(n12504) );
  XNOR U13305 ( .A(n12503), .B(n12504), .Z(c[1513]) );
  NANDN U13306 ( .A(n12485), .B(n12484), .Z(n12489) );
  NAND U13307 ( .A(n12487), .B(n12486), .Z(n12488) );
  NAND U13308 ( .A(n12489), .B(n12488), .Z(n12510) );
  AND U13309 ( .A(b[2]), .B(a[492]), .Z(n12516) );
  AND U13310 ( .A(a[493]), .B(b[1]), .Z(n12514) );
  AND U13311 ( .A(a[491]), .B(b[3]), .Z(n12513) );
  XOR U13312 ( .A(n12514), .B(n12513), .Z(n12515) );
  XOR U13313 ( .A(n12516), .B(n12515), .Z(n12519) );
  NAND U13314 ( .A(b[0]), .B(a[494]), .Z(n12520) );
  XOR U13315 ( .A(n12519), .B(n12520), .Z(n12522) );
  OR U13316 ( .A(n12491), .B(n12490), .Z(n12495) );
  NANDN U13317 ( .A(n12493), .B(n12492), .Z(n12494) );
  NAND U13318 ( .A(n12495), .B(n12494), .Z(n12521) );
  XNOR U13319 ( .A(n12522), .B(n12521), .Z(n12507) );
  NANDN U13320 ( .A(n12497), .B(n12496), .Z(n12501) );
  OR U13321 ( .A(n12499), .B(n12498), .Z(n12500) );
  NAND U13322 ( .A(n12501), .B(n12500), .Z(n12508) );
  XNOR U13323 ( .A(n12507), .B(n12508), .Z(n12509) );
  XNOR U13324 ( .A(n12510), .B(n12509), .Z(n12525) );
  XNOR U13325 ( .A(n12525), .B(sreg[1514]), .Z(n12527) );
  NAND U13326 ( .A(n12502), .B(sreg[1513]), .Z(n12506) );
  NANDN U13327 ( .A(n12504), .B(n12503), .Z(n12505) );
  AND U13328 ( .A(n12506), .B(n12505), .Z(n12526) );
  XOR U13329 ( .A(n12527), .B(n12526), .Z(c[1514]) );
  NANDN U13330 ( .A(n12508), .B(n12507), .Z(n12512) );
  NAND U13331 ( .A(n12510), .B(n12509), .Z(n12511) );
  NAND U13332 ( .A(n12512), .B(n12511), .Z(n12536) );
  AND U13333 ( .A(b[2]), .B(a[493]), .Z(n12542) );
  AND U13334 ( .A(a[494]), .B(b[1]), .Z(n12540) );
  AND U13335 ( .A(a[492]), .B(b[3]), .Z(n12539) );
  XOR U13336 ( .A(n12540), .B(n12539), .Z(n12541) );
  XOR U13337 ( .A(n12542), .B(n12541), .Z(n12545) );
  NAND U13338 ( .A(b[0]), .B(a[495]), .Z(n12546) );
  XOR U13339 ( .A(n12545), .B(n12546), .Z(n12548) );
  OR U13340 ( .A(n12514), .B(n12513), .Z(n12518) );
  NANDN U13341 ( .A(n12516), .B(n12515), .Z(n12517) );
  NAND U13342 ( .A(n12518), .B(n12517), .Z(n12547) );
  XNOR U13343 ( .A(n12548), .B(n12547), .Z(n12533) );
  NANDN U13344 ( .A(n12520), .B(n12519), .Z(n12524) );
  OR U13345 ( .A(n12522), .B(n12521), .Z(n12523) );
  NAND U13346 ( .A(n12524), .B(n12523), .Z(n12534) );
  XNOR U13347 ( .A(n12533), .B(n12534), .Z(n12535) );
  XNOR U13348 ( .A(n12536), .B(n12535), .Z(n12532) );
  NAND U13349 ( .A(n12525), .B(sreg[1514]), .Z(n12529) );
  OR U13350 ( .A(n12527), .B(n12526), .Z(n12528) );
  AND U13351 ( .A(n12529), .B(n12528), .Z(n12531) );
  XNOR U13352 ( .A(n12531), .B(sreg[1515]), .Z(n12530) );
  XOR U13353 ( .A(n12532), .B(n12530), .Z(c[1515]) );
  NANDN U13354 ( .A(n12534), .B(n12533), .Z(n12538) );
  NAND U13355 ( .A(n12536), .B(n12535), .Z(n12537) );
  NAND U13356 ( .A(n12538), .B(n12537), .Z(n12554) );
  AND U13357 ( .A(b[2]), .B(a[494]), .Z(n12560) );
  AND U13358 ( .A(a[495]), .B(b[1]), .Z(n12558) );
  AND U13359 ( .A(a[493]), .B(b[3]), .Z(n12557) );
  XOR U13360 ( .A(n12558), .B(n12557), .Z(n12559) );
  XOR U13361 ( .A(n12560), .B(n12559), .Z(n12563) );
  NAND U13362 ( .A(b[0]), .B(a[496]), .Z(n12564) );
  XOR U13363 ( .A(n12563), .B(n12564), .Z(n12566) );
  OR U13364 ( .A(n12540), .B(n12539), .Z(n12544) );
  NANDN U13365 ( .A(n12542), .B(n12541), .Z(n12543) );
  NAND U13366 ( .A(n12544), .B(n12543), .Z(n12565) );
  XNOR U13367 ( .A(n12566), .B(n12565), .Z(n12551) );
  NANDN U13368 ( .A(n12546), .B(n12545), .Z(n12550) );
  OR U13369 ( .A(n12548), .B(n12547), .Z(n12549) );
  NAND U13370 ( .A(n12550), .B(n12549), .Z(n12552) );
  XNOR U13371 ( .A(n12551), .B(n12552), .Z(n12553) );
  XOR U13372 ( .A(n12554), .B(n12553), .Z(n12569) );
  XOR U13373 ( .A(sreg[1516]), .B(n12569), .Z(n12571) );
  XNOR U13374 ( .A(n12570), .B(n12571), .Z(c[1516]) );
  NANDN U13375 ( .A(n12552), .B(n12551), .Z(n12556) );
  NAND U13376 ( .A(n12554), .B(n12553), .Z(n12555) );
  NAND U13377 ( .A(n12556), .B(n12555), .Z(n12577) );
  AND U13378 ( .A(b[2]), .B(a[495]), .Z(n12583) );
  AND U13379 ( .A(a[496]), .B(b[1]), .Z(n12581) );
  AND U13380 ( .A(a[494]), .B(b[3]), .Z(n12580) );
  XOR U13381 ( .A(n12581), .B(n12580), .Z(n12582) );
  XOR U13382 ( .A(n12583), .B(n12582), .Z(n12586) );
  NAND U13383 ( .A(b[0]), .B(a[497]), .Z(n12587) );
  XOR U13384 ( .A(n12586), .B(n12587), .Z(n12589) );
  OR U13385 ( .A(n12558), .B(n12557), .Z(n12562) );
  NANDN U13386 ( .A(n12560), .B(n12559), .Z(n12561) );
  NAND U13387 ( .A(n12562), .B(n12561), .Z(n12588) );
  XNOR U13388 ( .A(n12589), .B(n12588), .Z(n12574) );
  NANDN U13389 ( .A(n12564), .B(n12563), .Z(n12568) );
  OR U13390 ( .A(n12566), .B(n12565), .Z(n12567) );
  NAND U13391 ( .A(n12568), .B(n12567), .Z(n12575) );
  XNOR U13392 ( .A(n12574), .B(n12575), .Z(n12576) );
  XNOR U13393 ( .A(n12577), .B(n12576), .Z(n12592) );
  XOR U13394 ( .A(sreg[1517]), .B(n12592), .Z(n12593) );
  NANDN U13395 ( .A(n12569), .B(sreg[1516]), .Z(n12573) );
  NANDN U13396 ( .A(n12571), .B(n12570), .Z(n12572) );
  NAND U13397 ( .A(n12573), .B(n12572), .Z(n12594) );
  XOR U13398 ( .A(n12593), .B(n12594), .Z(c[1517]) );
  NANDN U13399 ( .A(n12575), .B(n12574), .Z(n12579) );
  NAND U13400 ( .A(n12577), .B(n12576), .Z(n12578) );
  NAND U13401 ( .A(n12579), .B(n12578), .Z(n12600) );
  AND U13402 ( .A(b[2]), .B(a[496]), .Z(n12606) );
  AND U13403 ( .A(a[497]), .B(b[1]), .Z(n12604) );
  AND U13404 ( .A(a[495]), .B(b[3]), .Z(n12603) );
  XOR U13405 ( .A(n12604), .B(n12603), .Z(n12605) );
  XOR U13406 ( .A(n12606), .B(n12605), .Z(n12609) );
  NAND U13407 ( .A(b[0]), .B(a[498]), .Z(n12610) );
  XOR U13408 ( .A(n12609), .B(n12610), .Z(n12612) );
  OR U13409 ( .A(n12581), .B(n12580), .Z(n12585) );
  NANDN U13410 ( .A(n12583), .B(n12582), .Z(n12584) );
  NAND U13411 ( .A(n12585), .B(n12584), .Z(n12611) );
  XNOR U13412 ( .A(n12612), .B(n12611), .Z(n12597) );
  NANDN U13413 ( .A(n12587), .B(n12586), .Z(n12591) );
  OR U13414 ( .A(n12589), .B(n12588), .Z(n12590) );
  NAND U13415 ( .A(n12591), .B(n12590), .Z(n12598) );
  XNOR U13416 ( .A(n12597), .B(n12598), .Z(n12599) );
  XNOR U13417 ( .A(n12600), .B(n12599), .Z(n12615) );
  XNOR U13418 ( .A(n12615), .B(sreg[1518]), .Z(n12617) );
  OR U13419 ( .A(n12592), .B(sreg[1517]), .Z(n12596) );
  NANDN U13420 ( .A(n12594), .B(n12593), .Z(n12595) );
  NAND U13421 ( .A(n12596), .B(n12595), .Z(n12616) );
  XOR U13422 ( .A(n12617), .B(n12616), .Z(c[1518]) );
  NANDN U13423 ( .A(n12598), .B(n12597), .Z(n12602) );
  NAND U13424 ( .A(n12600), .B(n12599), .Z(n12601) );
  NAND U13425 ( .A(n12602), .B(n12601), .Z(n12623) );
  AND U13426 ( .A(b[2]), .B(a[497]), .Z(n12629) );
  AND U13427 ( .A(a[498]), .B(b[1]), .Z(n12627) );
  AND U13428 ( .A(a[496]), .B(b[3]), .Z(n12626) );
  XOR U13429 ( .A(n12627), .B(n12626), .Z(n12628) );
  XOR U13430 ( .A(n12629), .B(n12628), .Z(n12632) );
  NAND U13431 ( .A(b[0]), .B(a[499]), .Z(n12633) );
  XOR U13432 ( .A(n12632), .B(n12633), .Z(n12635) );
  OR U13433 ( .A(n12604), .B(n12603), .Z(n12608) );
  NANDN U13434 ( .A(n12606), .B(n12605), .Z(n12607) );
  NAND U13435 ( .A(n12608), .B(n12607), .Z(n12634) );
  XNOR U13436 ( .A(n12635), .B(n12634), .Z(n12620) );
  NANDN U13437 ( .A(n12610), .B(n12609), .Z(n12614) );
  OR U13438 ( .A(n12612), .B(n12611), .Z(n12613) );
  NAND U13439 ( .A(n12614), .B(n12613), .Z(n12621) );
  XNOR U13440 ( .A(n12620), .B(n12621), .Z(n12622) );
  XNOR U13441 ( .A(n12623), .B(n12622), .Z(n12638) );
  XNOR U13442 ( .A(n12638), .B(sreg[1519]), .Z(n12640) );
  NAND U13443 ( .A(n12615), .B(sreg[1518]), .Z(n12619) );
  OR U13444 ( .A(n12617), .B(n12616), .Z(n12618) );
  AND U13445 ( .A(n12619), .B(n12618), .Z(n12639) );
  XOR U13446 ( .A(n12640), .B(n12639), .Z(c[1519]) );
  NANDN U13447 ( .A(n12621), .B(n12620), .Z(n12625) );
  NAND U13448 ( .A(n12623), .B(n12622), .Z(n12624) );
  NAND U13449 ( .A(n12625), .B(n12624), .Z(n12649) );
  AND U13450 ( .A(b[2]), .B(a[498]), .Z(n12661) );
  AND U13451 ( .A(a[499]), .B(b[1]), .Z(n12659) );
  AND U13452 ( .A(a[497]), .B(b[3]), .Z(n12658) );
  XOR U13453 ( .A(n12659), .B(n12658), .Z(n12660) );
  XOR U13454 ( .A(n12661), .B(n12660), .Z(n12652) );
  NAND U13455 ( .A(b[0]), .B(a[500]), .Z(n12653) );
  XOR U13456 ( .A(n12652), .B(n12653), .Z(n12655) );
  OR U13457 ( .A(n12627), .B(n12626), .Z(n12631) );
  NANDN U13458 ( .A(n12629), .B(n12628), .Z(n12630) );
  NAND U13459 ( .A(n12631), .B(n12630), .Z(n12654) );
  XNOR U13460 ( .A(n12655), .B(n12654), .Z(n12646) );
  NANDN U13461 ( .A(n12633), .B(n12632), .Z(n12637) );
  OR U13462 ( .A(n12635), .B(n12634), .Z(n12636) );
  NAND U13463 ( .A(n12637), .B(n12636), .Z(n12647) );
  XNOR U13464 ( .A(n12646), .B(n12647), .Z(n12648) );
  XNOR U13465 ( .A(n12649), .B(n12648), .Z(n12645) );
  NAND U13466 ( .A(n12638), .B(sreg[1519]), .Z(n12642) );
  OR U13467 ( .A(n12640), .B(n12639), .Z(n12641) );
  AND U13468 ( .A(n12642), .B(n12641), .Z(n12644) );
  XNOR U13469 ( .A(n12644), .B(sreg[1520]), .Z(n12643) );
  XOR U13470 ( .A(n12645), .B(n12643), .Z(c[1520]) );
  NANDN U13471 ( .A(n12647), .B(n12646), .Z(n12651) );
  NAND U13472 ( .A(n12649), .B(n12648), .Z(n12650) );
  NAND U13473 ( .A(n12651), .B(n12650), .Z(n12679) );
  NANDN U13474 ( .A(n12653), .B(n12652), .Z(n12657) );
  OR U13475 ( .A(n12655), .B(n12654), .Z(n12656) );
  NAND U13476 ( .A(n12657), .B(n12656), .Z(n12676) );
  AND U13477 ( .A(b[2]), .B(a[499]), .Z(n12667) );
  AND U13478 ( .A(a[500]), .B(b[1]), .Z(n12665) );
  AND U13479 ( .A(a[498]), .B(b[3]), .Z(n12664) );
  XOR U13480 ( .A(n12665), .B(n12664), .Z(n12666) );
  XOR U13481 ( .A(n12667), .B(n12666), .Z(n12670) );
  NAND U13482 ( .A(b[0]), .B(a[501]), .Z(n12671) );
  XNOR U13483 ( .A(n12670), .B(n12671), .Z(n12672) );
  OR U13484 ( .A(n12659), .B(n12658), .Z(n12663) );
  NANDN U13485 ( .A(n12661), .B(n12660), .Z(n12662) );
  AND U13486 ( .A(n12663), .B(n12662), .Z(n12673) );
  XNOR U13487 ( .A(n12672), .B(n12673), .Z(n12677) );
  XNOR U13488 ( .A(n12676), .B(n12677), .Z(n12678) );
  XNOR U13489 ( .A(n12679), .B(n12678), .Z(n12682) );
  XNOR U13490 ( .A(sreg[1521]), .B(n12682), .Z(n12684) );
  XNOR U13491 ( .A(n12683), .B(n12684), .Z(c[1521]) );
  AND U13492 ( .A(b[2]), .B(a[500]), .Z(n12697) );
  AND U13493 ( .A(a[501]), .B(b[1]), .Z(n12695) );
  AND U13494 ( .A(a[499]), .B(b[3]), .Z(n12694) );
  XOR U13495 ( .A(n12695), .B(n12694), .Z(n12696) );
  XOR U13496 ( .A(n12697), .B(n12696), .Z(n12700) );
  NAND U13497 ( .A(b[0]), .B(a[502]), .Z(n12701) );
  XOR U13498 ( .A(n12700), .B(n12701), .Z(n12703) );
  OR U13499 ( .A(n12665), .B(n12664), .Z(n12669) );
  NANDN U13500 ( .A(n12667), .B(n12666), .Z(n12668) );
  NAND U13501 ( .A(n12669), .B(n12668), .Z(n12702) );
  XNOR U13502 ( .A(n12703), .B(n12702), .Z(n12688) );
  NANDN U13503 ( .A(n12671), .B(n12670), .Z(n12675) );
  NAND U13504 ( .A(n12673), .B(n12672), .Z(n12674) );
  NAND U13505 ( .A(n12675), .B(n12674), .Z(n12689) );
  XNOR U13506 ( .A(n12688), .B(n12689), .Z(n12690) );
  NANDN U13507 ( .A(n12677), .B(n12676), .Z(n12681) );
  NANDN U13508 ( .A(n12679), .B(n12678), .Z(n12680) );
  AND U13509 ( .A(n12681), .B(n12680), .Z(n12691) );
  XNOR U13510 ( .A(n12690), .B(n12691), .Z(n12707) );
  NAND U13511 ( .A(sreg[1521]), .B(n12682), .Z(n12686) );
  NANDN U13512 ( .A(n12684), .B(n12683), .Z(n12685) );
  AND U13513 ( .A(n12686), .B(n12685), .Z(n12706) );
  XNOR U13514 ( .A(sreg[1522]), .B(n12706), .Z(n12687) );
  XOR U13515 ( .A(n12707), .B(n12687), .Z(c[1522]) );
  NANDN U13516 ( .A(n12689), .B(n12688), .Z(n12693) );
  NAND U13517 ( .A(n12691), .B(n12690), .Z(n12692) );
  NAND U13518 ( .A(n12693), .B(n12692), .Z(n12723) );
  AND U13519 ( .A(b[2]), .B(a[501]), .Z(n12717) );
  AND U13520 ( .A(a[502]), .B(b[1]), .Z(n12715) );
  AND U13521 ( .A(a[500]), .B(b[3]), .Z(n12714) );
  XOR U13522 ( .A(n12715), .B(n12714), .Z(n12716) );
  XOR U13523 ( .A(n12717), .B(n12716), .Z(n12708) );
  NAND U13524 ( .A(b[0]), .B(a[503]), .Z(n12709) );
  XOR U13525 ( .A(n12708), .B(n12709), .Z(n12711) );
  OR U13526 ( .A(n12695), .B(n12694), .Z(n12699) );
  NANDN U13527 ( .A(n12697), .B(n12696), .Z(n12698) );
  NAND U13528 ( .A(n12699), .B(n12698), .Z(n12710) );
  XNOR U13529 ( .A(n12711), .B(n12710), .Z(n12720) );
  NANDN U13530 ( .A(n12701), .B(n12700), .Z(n12705) );
  OR U13531 ( .A(n12703), .B(n12702), .Z(n12704) );
  NAND U13532 ( .A(n12705), .B(n12704), .Z(n12721) );
  XNOR U13533 ( .A(n12720), .B(n12721), .Z(n12722) );
  XNOR U13534 ( .A(n12723), .B(n12722), .Z(n12726) );
  XOR U13535 ( .A(sreg[1523]), .B(n12726), .Z(n12727) );
  XOR U13536 ( .A(n12727), .B(n12728), .Z(c[1523]) );
  NANDN U13537 ( .A(n12709), .B(n12708), .Z(n12713) );
  OR U13538 ( .A(n12711), .B(n12710), .Z(n12712) );
  NAND U13539 ( .A(n12713), .B(n12712), .Z(n12746) );
  AND U13540 ( .A(b[2]), .B(a[502]), .Z(n12737) );
  AND U13541 ( .A(a[503]), .B(b[1]), .Z(n12735) );
  AND U13542 ( .A(a[501]), .B(b[3]), .Z(n12734) );
  XOR U13543 ( .A(n12735), .B(n12734), .Z(n12736) );
  XOR U13544 ( .A(n12737), .B(n12736), .Z(n12740) );
  NAND U13545 ( .A(b[0]), .B(a[504]), .Z(n12741) );
  XNOR U13546 ( .A(n12740), .B(n12741), .Z(n12742) );
  OR U13547 ( .A(n12715), .B(n12714), .Z(n12719) );
  NANDN U13548 ( .A(n12717), .B(n12716), .Z(n12718) );
  AND U13549 ( .A(n12719), .B(n12718), .Z(n12743) );
  XNOR U13550 ( .A(n12742), .B(n12743), .Z(n12747) );
  XNOR U13551 ( .A(n12746), .B(n12747), .Z(n12748) );
  NANDN U13552 ( .A(n12721), .B(n12720), .Z(n12725) );
  NAND U13553 ( .A(n12723), .B(n12722), .Z(n12724) );
  AND U13554 ( .A(n12725), .B(n12724), .Z(n12749) );
  XNOR U13555 ( .A(n12748), .B(n12749), .Z(n12733) );
  OR U13556 ( .A(n12726), .B(sreg[1523]), .Z(n12730) );
  NANDN U13557 ( .A(n12728), .B(n12727), .Z(n12729) );
  AND U13558 ( .A(n12730), .B(n12729), .Z(n12732) );
  XNOR U13559 ( .A(sreg[1524]), .B(n12732), .Z(n12731) );
  XOR U13560 ( .A(n12733), .B(n12731), .Z(c[1524]) );
  AND U13561 ( .A(b[2]), .B(a[503]), .Z(n12761) );
  AND U13562 ( .A(a[504]), .B(b[1]), .Z(n12759) );
  AND U13563 ( .A(a[502]), .B(b[3]), .Z(n12758) );
  XOR U13564 ( .A(n12759), .B(n12758), .Z(n12760) );
  XOR U13565 ( .A(n12761), .B(n12760), .Z(n12764) );
  NAND U13566 ( .A(b[0]), .B(a[505]), .Z(n12765) );
  XOR U13567 ( .A(n12764), .B(n12765), .Z(n12767) );
  OR U13568 ( .A(n12735), .B(n12734), .Z(n12739) );
  NANDN U13569 ( .A(n12737), .B(n12736), .Z(n12738) );
  NAND U13570 ( .A(n12739), .B(n12738), .Z(n12766) );
  XNOR U13571 ( .A(n12767), .B(n12766), .Z(n12752) );
  NANDN U13572 ( .A(n12741), .B(n12740), .Z(n12745) );
  NAND U13573 ( .A(n12743), .B(n12742), .Z(n12744) );
  NAND U13574 ( .A(n12745), .B(n12744), .Z(n12753) );
  XNOR U13575 ( .A(n12752), .B(n12753), .Z(n12754) );
  NANDN U13576 ( .A(n12747), .B(n12746), .Z(n12751) );
  NAND U13577 ( .A(n12749), .B(n12748), .Z(n12750) );
  NAND U13578 ( .A(n12751), .B(n12750), .Z(n12755) );
  XOR U13579 ( .A(n12754), .B(n12755), .Z(n12770) );
  XNOR U13580 ( .A(n12770), .B(sreg[1525]), .Z(n12771) );
  XOR U13581 ( .A(n12772), .B(n12771), .Z(c[1525]) );
  NANDN U13582 ( .A(n12753), .B(n12752), .Z(n12757) );
  NANDN U13583 ( .A(n12755), .B(n12754), .Z(n12756) );
  NAND U13584 ( .A(n12757), .B(n12756), .Z(n12791) );
  AND U13585 ( .A(b[2]), .B(a[504]), .Z(n12785) );
  AND U13586 ( .A(a[505]), .B(b[1]), .Z(n12783) );
  AND U13587 ( .A(a[503]), .B(b[3]), .Z(n12782) );
  XOR U13588 ( .A(n12783), .B(n12782), .Z(n12784) );
  XOR U13589 ( .A(n12785), .B(n12784), .Z(n12776) );
  NAND U13590 ( .A(b[0]), .B(a[506]), .Z(n12777) );
  XOR U13591 ( .A(n12776), .B(n12777), .Z(n12779) );
  OR U13592 ( .A(n12759), .B(n12758), .Z(n12763) );
  NANDN U13593 ( .A(n12761), .B(n12760), .Z(n12762) );
  NAND U13594 ( .A(n12763), .B(n12762), .Z(n12778) );
  XNOR U13595 ( .A(n12779), .B(n12778), .Z(n12788) );
  NANDN U13596 ( .A(n12765), .B(n12764), .Z(n12769) );
  OR U13597 ( .A(n12767), .B(n12766), .Z(n12768) );
  NAND U13598 ( .A(n12769), .B(n12768), .Z(n12789) );
  XNOR U13599 ( .A(n12788), .B(n12789), .Z(n12790) );
  XOR U13600 ( .A(n12791), .B(n12790), .Z(n12795) );
  NAND U13601 ( .A(n12770), .B(sreg[1525]), .Z(n12774) );
  OR U13602 ( .A(n12772), .B(n12771), .Z(n12773) );
  NAND U13603 ( .A(n12774), .B(n12773), .Z(n12794) );
  XNOR U13604 ( .A(sreg[1526]), .B(n12794), .Z(n12775) );
  XOR U13605 ( .A(n12795), .B(n12775), .Z(c[1526]) );
  NANDN U13606 ( .A(n12777), .B(n12776), .Z(n12781) );
  OR U13607 ( .A(n12779), .B(n12778), .Z(n12780) );
  NAND U13608 ( .A(n12781), .B(n12780), .Z(n12797) );
  AND U13609 ( .A(b[2]), .B(a[505]), .Z(n12812) );
  AND U13610 ( .A(a[506]), .B(b[1]), .Z(n12810) );
  AND U13611 ( .A(a[504]), .B(b[3]), .Z(n12809) );
  XOR U13612 ( .A(n12810), .B(n12809), .Z(n12811) );
  XOR U13613 ( .A(n12812), .B(n12811), .Z(n12803) );
  NAND U13614 ( .A(b[0]), .B(a[507]), .Z(n12804) );
  XNOR U13615 ( .A(n12803), .B(n12804), .Z(n12805) );
  OR U13616 ( .A(n12783), .B(n12782), .Z(n12787) );
  NANDN U13617 ( .A(n12785), .B(n12784), .Z(n12786) );
  AND U13618 ( .A(n12787), .B(n12786), .Z(n12806) );
  XNOR U13619 ( .A(n12805), .B(n12806), .Z(n12798) );
  XNOR U13620 ( .A(n12797), .B(n12798), .Z(n12799) );
  NANDN U13621 ( .A(n12789), .B(n12788), .Z(n12793) );
  NAND U13622 ( .A(n12791), .B(n12790), .Z(n12792) );
  AND U13623 ( .A(n12793), .B(n12792), .Z(n12800) );
  XNOR U13624 ( .A(n12799), .B(n12800), .Z(n12818) );
  IV U13625 ( .A(n12816), .Z(n12815) );
  XNOR U13626 ( .A(n12815), .B(sreg[1527]), .Z(n12796) );
  XOR U13627 ( .A(n12818), .B(n12796), .Z(c[1527]) );
  NANDN U13628 ( .A(n12798), .B(n12797), .Z(n12802) );
  NAND U13629 ( .A(n12800), .B(n12799), .Z(n12801) );
  NAND U13630 ( .A(n12802), .B(n12801), .Z(n12827) );
  NANDN U13631 ( .A(n12804), .B(n12803), .Z(n12808) );
  NAND U13632 ( .A(n12806), .B(n12805), .Z(n12807) );
  NAND U13633 ( .A(n12808), .B(n12807), .Z(n12824) );
  AND U13634 ( .A(b[2]), .B(a[506]), .Z(n12833) );
  AND U13635 ( .A(a[507]), .B(b[1]), .Z(n12831) );
  AND U13636 ( .A(a[505]), .B(b[3]), .Z(n12830) );
  XOR U13637 ( .A(n12831), .B(n12830), .Z(n12832) );
  XOR U13638 ( .A(n12833), .B(n12832), .Z(n12836) );
  NAND U13639 ( .A(b[0]), .B(a[508]), .Z(n12837) );
  XNOR U13640 ( .A(n12836), .B(n12837), .Z(n12838) );
  OR U13641 ( .A(n12810), .B(n12809), .Z(n12814) );
  NANDN U13642 ( .A(n12812), .B(n12811), .Z(n12813) );
  AND U13643 ( .A(n12814), .B(n12813), .Z(n12839) );
  XNOR U13644 ( .A(n12838), .B(n12839), .Z(n12825) );
  XNOR U13645 ( .A(n12824), .B(n12825), .Z(n12826) );
  XOR U13646 ( .A(n12827), .B(n12826), .Z(n12823) );
  NAND U13647 ( .A(n12815), .B(sreg[1527]), .Z(n12820) );
  NANDN U13648 ( .A(sreg[1527]), .B(n12816), .Z(n12817) );
  NANDN U13649 ( .A(n12818), .B(n12817), .Z(n12819) );
  AND U13650 ( .A(n12820), .B(n12819), .Z(n12822) );
  XNOR U13651 ( .A(n12822), .B(sreg[1528]), .Z(n12821) );
  XOR U13652 ( .A(n12823), .B(n12821), .Z(c[1528]) );
  NANDN U13653 ( .A(n12825), .B(n12824), .Z(n12829) );
  NAND U13654 ( .A(n12827), .B(n12826), .Z(n12828) );
  NAND U13655 ( .A(n12829), .B(n12828), .Z(n12862) );
  AND U13656 ( .A(b[2]), .B(a[507]), .Z(n12856) );
  AND U13657 ( .A(a[508]), .B(b[1]), .Z(n12854) );
  AND U13658 ( .A(a[506]), .B(b[3]), .Z(n12853) );
  XOR U13659 ( .A(n12854), .B(n12853), .Z(n12855) );
  XOR U13660 ( .A(n12856), .B(n12855), .Z(n12847) );
  NAND U13661 ( .A(b[0]), .B(a[509]), .Z(n12848) );
  XOR U13662 ( .A(n12847), .B(n12848), .Z(n12850) );
  OR U13663 ( .A(n12831), .B(n12830), .Z(n12835) );
  NANDN U13664 ( .A(n12833), .B(n12832), .Z(n12834) );
  NAND U13665 ( .A(n12835), .B(n12834), .Z(n12849) );
  XNOR U13666 ( .A(n12850), .B(n12849), .Z(n12859) );
  NANDN U13667 ( .A(n12837), .B(n12836), .Z(n12841) );
  NAND U13668 ( .A(n12839), .B(n12838), .Z(n12840) );
  NAND U13669 ( .A(n12841), .B(n12840), .Z(n12860) );
  XNOR U13670 ( .A(n12859), .B(n12860), .Z(n12861) );
  XOR U13671 ( .A(n12862), .B(n12861), .Z(n12842) );
  XNOR U13672 ( .A(n12842), .B(sreg[1529]), .Z(n12844) );
  XNOR U13673 ( .A(n12843), .B(n12844), .Z(c[1529]) );
  NAND U13674 ( .A(n12842), .B(sreg[1529]), .Z(n12846) );
  NANDN U13675 ( .A(n12844), .B(n12843), .Z(n12845) );
  NAND U13676 ( .A(n12846), .B(n12845), .Z(n12866) );
  NANDN U13677 ( .A(n12848), .B(n12847), .Z(n12852) );
  OR U13678 ( .A(n12850), .B(n12849), .Z(n12851) );
  NAND U13679 ( .A(n12852), .B(n12851), .Z(n12868) );
  AND U13680 ( .A(b[2]), .B(a[508]), .Z(n12883) );
  AND U13681 ( .A(a[509]), .B(b[1]), .Z(n12881) );
  AND U13682 ( .A(a[507]), .B(b[3]), .Z(n12880) );
  XOR U13683 ( .A(n12881), .B(n12880), .Z(n12882) );
  XOR U13684 ( .A(n12883), .B(n12882), .Z(n12874) );
  NAND U13685 ( .A(b[0]), .B(a[510]), .Z(n12875) );
  XNOR U13686 ( .A(n12874), .B(n12875), .Z(n12876) );
  OR U13687 ( .A(n12854), .B(n12853), .Z(n12858) );
  NANDN U13688 ( .A(n12856), .B(n12855), .Z(n12857) );
  AND U13689 ( .A(n12858), .B(n12857), .Z(n12877) );
  XNOR U13690 ( .A(n12876), .B(n12877), .Z(n12869) );
  XNOR U13691 ( .A(n12868), .B(n12869), .Z(n12870) );
  NANDN U13692 ( .A(n12860), .B(n12859), .Z(n12864) );
  NANDN U13693 ( .A(n12862), .B(n12861), .Z(n12863) );
  AND U13694 ( .A(n12864), .B(n12863), .Z(n12871) );
  XNOR U13695 ( .A(n12870), .B(n12871), .Z(n12867) );
  XOR U13696 ( .A(sreg[1530]), .B(n12867), .Z(n12865) );
  XNOR U13697 ( .A(n12866), .B(n12865), .Z(c[1530]) );
  NANDN U13698 ( .A(n12869), .B(n12868), .Z(n12873) );
  NAND U13699 ( .A(n12871), .B(n12870), .Z(n12872) );
  NAND U13700 ( .A(n12873), .B(n12872), .Z(n12889) );
  NANDN U13701 ( .A(n12875), .B(n12874), .Z(n12879) );
  NAND U13702 ( .A(n12877), .B(n12876), .Z(n12878) );
  NAND U13703 ( .A(n12879), .B(n12878), .Z(n12886) );
  AND U13704 ( .A(b[2]), .B(a[509]), .Z(n12895) );
  AND U13705 ( .A(a[510]), .B(b[1]), .Z(n12893) );
  AND U13706 ( .A(a[508]), .B(b[3]), .Z(n12892) );
  XOR U13707 ( .A(n12893), .B(n12892), .Z(n12894) );
  XOR U13708 ( .A(n12895), .B(n12894), .Z(n12898) );
  NAND U13709 ( .A(b[0]), .B(a[511]), .Z(n12899) );
  XNOR U13710 ( .A(n12898), .B(n12899), .Z(n12900) );
  OR U13711 ( .A(n12881), .B(n12880), .Z(n12885) );
  NANDN U13712 ( .A(n12883), .B(n12882), .Z(n12884) );
  AND U13713 ( .A(n12885), .B(n12884), .Z(n12901) );
  XNOR U13714 ( .A(n12900), .B(n12901), .Z(n12887) );
  XNOR U13715 ( .A(n12886), .B(n12887), .Z(n12888) );
  XOR U13716 ( .A(n12889), .B(n12888), .Z(n12904) );
  XNOR U13717 ( .A(sreg[1531]), .B(n12904), .Z(n12905) );
  XOR U13718 ( .A(n12906), .B(n12905), .Z(c[1531]) );
  NANDN U13719 ( .A(n12887), .B(n12886), .Z(n12891) );
  NAND U13720 ( .A(n12889), .B(n12888), .Z(n12890) );
  NAND U13721 ( .A(n12891), .B(n12890), .Z(n12927) );
  AND U13722 ( .A(b[2]), .B(a[510]), .Z(n12921) );
  AND U13723 ( .A(a[511]), .B(b[1]), .Z(n12919) );
  AND U13724 ( .A(a[509]), .B(b[3]), .Z(n12918) );
  XOR U13725 ( .A(n12919), .B(n12918), .Z(n12920) );
  XOR U13726 ( .A(n12921), .B(n12920), .Z(n12912) );
  NAND U13727 ( .A(b[0]), .B(a[512]), .Z(n12913) );
  XOR U13728 ( .A(n12912), .B(n12913), .Z(n12915) );
  OR U13729 ( .A(n12893), .B(n12892), .Z(n12897) );
  NANDN U13730 ( .A(n12895), .B(n12894), .Z(n12896) );
  NAND U13731 ( .A(n12897), .B(n12896), .Z(n12914) );
  XNOR U13732 ( .A(n12915), .B(n12914), .Z(n12924) );
  NANDN U13733 ( .A(n12899), .B(n12898), .Z(n12903) );
  NAND U13734 ( .A(n12901), .B(n12900), .Z(n12902) );
  NAND U13735 ( .A(n12903), .B(n12902), .Z(n12925) );
  XNOR U13736 ( .A(n12924), .B(n12925), .Z(n12926) );
  XOR U13737 ( .A(n12927), .B(n12926), .Z(n12911) );
  NAND U13738 ( .A(sreg[1531]), .B(n12904), .Z(n12908) );
  OR U13739 ( .A(n12906), .B(n12905), .Z(n12907) );
  NAND U13740 ( .A(n12908), .B(n12907), .Z(n12910) );
  XNOR U13741 ( .A(sreg[1532]), .B(n12910), .Z(n12909) );
  XNOR U13742 ( .A(n12911), .B(n12909), .Z(c[1532]) );
  NANDN U13743 ( .A(n12913), .B(n12912), .Z(n12917) );
  OR U13744 ( .A(n12915), .B(n12914), .Z(n12916) );
  NAND U13745 ( .A(n12917), .B(n12916), .Z(n12930) );
  AND U13746 ( .A(b[2]), .B(a[511]), .Z(n12945) );
  AND U13747 ( .A(a[512]), .B(b[1]), .Z(n12943) );
  AND U13748 ( .A(a[510]), .B(b[3]), .Z(n12942) );
  XOR U13749 ( .A(n12943), .B(n12942), .Z(n12944) );
  XOR U13750 ( .A(n12945), .B(n12944), .Z(n12936) );
  NAND U13751 ( .A(b[0]), .B(a[513]), .Z(n12937) );
  XNOR U13752 ( .A(n12936), .B(n12937), .Z(n12938) );
  OR U13753 ( .A(n12919), .B(n12918), .Z(n12923) );
  NANDN U13754 ( .A(n12921), .B(n12920), .Z(n12922) );
  AND U13755 ( .A(n12923), .B(n12922), .Z(n12939) );
  XNOR U13756 ( .A(n12938), .B(n12939), .Z(n12931) );
  XNOR U13757 ( .A(n12930), .B(n12931), .Z(n12932) );
  NANDN U13758 ( .A(n12925), .B(n12924), .Z(n12929) );
  NANDN U13759 ( .A(n12927), .B(n12926), .Z(n12928) );
  NAND U13760 ( .A(n12929), .B(n12928), .Z(n12933) );
  XOR U13761 ( .A(n12932), .B(n12933), .Z(n12948) );
  XNOR U13762 ( .A(sreg[1533]), .B(n12948), .Z(n12949) );
  XNOR U13763 ( .A(n12950), .B(n12949), .Z(c[1533]) );
  NANDN U13764 ( .A(n12931), .B(n12930), .Z(n12935) );
  NANDN U13765 ( .A(n12933), .B(n12932), .Z(n12934) );
  NAND U13766 ( .A(n12935), .B(n12934), .Z(n12956) );
  NANDN U13767 ( .A(n12937), .B(n12936), .Z(n12941) );
  NAND U13768 ( .A(n12939), .B(n12938), .Z(n12940) );
  NAND U13769 ( .A(n12941), .B(n12940), .Z(n12953) );
  AND U13770 ( .A(b[2]), .B(a[512]), .Z(n12962) );
  AND U13771 ( .A(a[513]), .B(b[1]), .Z(n12960) );
  AND U13772 ( .A(a[511]), .B(b[3]), .Z(n12959) );
  XOR U13773 ( .A(n12960), .B(n12959), .Z(n12961) );
  XOR U13774 ( .A(n12962), .B(n12961), .Z(n12965) );
  NAND U13775 ( .A(b[0]), .B(a[514]), .Z(n12966) );
  XNOR U13776 ( .A(n12965), .B(n12966), .Z(n12967) );
  OR U13777 ( .A(n12943), .B(n12942), .Z(n12947) );
  NANDN U13778 ( .A(n12945), .B(n12944), .Z(n12946) );
  AND U13779 ( .A(n12947), .B(n12946), .Z(n12968) );
  XNOR U13780 ( .A(n12967), .B(n12968), .Z(n12954) );
  XNOR U13781 ( .A(n12953), .B(n12954), .Z(n12955) );
  XOR U13782 ( .A(n12956), .B(n12955), .Z(n12971) );
  XOR U13783 ( .A(sreg[1534]), .B(n12971), .Z(n12972) );
  NANDN U13784 ( .A(sreg[1533]), .B(n12948), .Z(n12952) );
  NAND U13785 ( .A(n12950), .B(n12949), .Z(n12951) );
  AND U13786 ( .A(n12952), .B(n12951), .Z(n12973) );
  XOR U13787 ( .A(n12972), .B(n12973), .Z(c[1534]) );
  NANDN U13788 ( .A(n12954), .B(n12953), .Z(n12958) );
  NAND U13789 ( .A(n12956), .B(n12955), .Z(n12957) );
  NAND U13790 ( .A(n12958), .B(n12957), .Z(n12982) );
  AND U13791 ( .A(b[2]), .B(a[513]), .Z(n12988) );
  AND U13792 ( .A(a[514]), .B(b[1]), .Z(n12986) );
  AND U13793 ( .A(a[512]), .B(b[3]), .Z(n12985) );
  XOR U13794 ( .A(n12986), .B(n12985), .Z(n12987) );
  XOR U13795 ( .A(n12988), .B(n12987), .Z(n12991) );
  NAND U13796 ( .A(b[0]), .B(a[515]), .Z(n12992) );
  XOR U13797 ( .A(n12991), .B(n12992), .Z(n12994) );
  OR U13798 ( .A(n12960), .B(n12959), .Z(n12964) );
  NANDN U13799 ( .A(n12962), .B(n12961), .Z(n12963) );
  NAND U13800 ( .A(n12964), .B(n12963), .Z(n12993) );
  XNOR U13801 ( .A(n12994), .B(n12993), .Z(n12979) );
  NANDN U13802 ( .A(n12966), .B(n12965), .Z(n12970) );
  NAND U13803 ( .A(n12968), .B(n12967), .Z(n12969) );
  NAND U13804 ( .A(n12970), .B(n12969), .Z(n12980) );
  XNOR U13805 ( .A(n12979), .B(n12980), .Z(n12981) );
  XOR U13806 ( .A(n12982), .B(n12981), .Z(n12978) );
  OR U13807 ( .A(n12971), .B(sreg[1534]), .Z(n12975) );
  NANDN U13808 ( .A(n12973), .B(n12972), .Z(n12974) );
  AND U13809 ( .A(n12975), .B(n12974), .Z(n12977) );
  XNOR U13810 ( .A(sreg[1535]), .B(n12977), .Z(n12976) );
  XNOR U13811 ( .A(n12978), .B(n12976), .Z(c[1535]) );
  NANDN U13812 ( .A(n12980), .B(n12979), .Z(n12984) );
  NANDN U13813 ( .A(n12982), .B(n12981), .Z(n12983) );
  AND U13814 ( .A(n12984), .B(n12983), .Z(n13000) );
  AND U13815 ( .A(b[2]), .B(a[514]), .Z(n13008) );
  AND U13816 ( .A(a[515]), .B(b[1]), .Z(n13006) );
  AND U13817 ( .A(a[513]), .B(b[3]), .Z(n13005) );
  XOR U13818 ( .A(n13006), .B(n13005), .Z(n13007) );
  XOR U13819 ( .A(n13008), .B(n13007), .Z(n13001) );
  NAND U13820 ( .A(b[0]), .B(a[516]), .Z(n13002) );
  XOR U13821 ( .A(n13001), .B(n13002), .Z(n13003) );
  OR U13822 ( .A(n12986), .B(n12985), .Z(n12990) );
  NANDN U13823 ( .A(n12988), .B(n12987), .Z(n12989) );
  AND U13824 ( .A(n12990), .B(n12989), .Z(n13004) );
  XOR U13825 ( .A(n13003), .B(n13004), .Z(n12998) );
  NANDN U13826 ( .A(n12992), .B(n12991), .Z(n12996) );
  OR U13827 ( .A(n12994), .B(n12993), .Z(n12995) );
  AND U13828 ( .A(n12996), .B(n12995), .Z(n12999) );
  XOR U13829 ( .A(n12998), .B(n12999), .Z(n12997) );
  XOR U13830 ( .A(n13000), .B(n12997), .Z(n13011) );
  XNOR U13831 ( .A(sreg[1536]), .B(n13011), .Z(n13012) );
  XOR U13832 ( .A(n13013), .B(n13012), .Z(c[1536]) );
  AND U13833 ( .A(b[2]), .B(a[515]), .Z(n13025) );
  AND U13834 ( .A(a[516]), .B(b[1]), .Z(n13023) );
  AND U13835 ( .A(a[514]), .B(b[3]), .Z(n13022) );
  XOR U13836 ( .A(n13023), .B(n13022), .Z(n13024) );
  XOR U13837 ( .A(n13025), .B(n13024), .Z(n13028) );
  NAND U13838 ( .A(b[0]), .B(a[517]), .Z(n13029) );
  XNOR U13839 ( .A(n13028), .B(n13029), .Z(n13030) );
  OR U13840 ( .A(n13006), .B(n13005), .Z(n13010) );
  NANDN U13841 ( .A(n13008), .B(n13007), .Z(n13009) );
  AND U13842 ( .A(n13010), .B(n13009), .Z(n13031) );
  XNOR U13843 ( .A(n13030), .B(n13031), .Z(n13017) );
  XNOR U13844 ( .A(n13016), .B(n13017), .Z(n13018) );
  XNOR U13845 ( .A(n13019), .B(n13018), .Z(n13034) );
  XOR U13846 ( .A(sreg[1537]), .B(n13034), .Z(n13035) );
  NAND U13847 ( .A(sreg[1536]), .B(n13011), .Z(n13015) );
  OR U13848 ( .A(n13013), .B(n13012), .Z(n13014) );
  NAND U13849 ( .A(n13015), .B(n13014), .Z(n13036) );
  XOR U13850 ( .A(n13035), .B(n13036), .Z(c[1537]) );
  NANDN U13851 ( .A(n13017), .B(n13016), .Z(n13021) );
  NANDN U13852 ( .A(n13019), .B(n13018), .Z(n13020) );
  NAND U13853 ( .A(n13021), .B(n13020), .Z(n13045) );
  AND U13854 ( .A(b[2]), .B(a[516]), .Z(n13051) );
  AND U13855 ( .A(a[517]), .B(b[1]), .Z(n13049) );
  AND U13856 ( .A(a[515]), .B(b[3]), .Z(n13048) );
  XOR U13857 ( .A(n13049), .B(n13048), .Z(n13050) );
  XOR U13858 ( .A(n13051), .B(n13050), .Z(n13054) );
  NAND U13859 ( .A(b[0]), .B(a[518]), .Z(n13055) );
  XOR U13860 ( .A(n13054), .B(n13055), .Z(n13057) );
  OR U13861 ( .A(n13023), .B(n13022), .Z(n13027) );
  NANDN U13862 ( .A(n13025), .B(n13024), .Z(n13026) );
  NAND U13863 ( .A(n13027), .B(n13026), .Z(n13056) );
  XNOR U13864 ( .A(n13057), .B(n13056), .Z(n13042) );
  NANDN U13865 ( .A(n13029), .B(n13028), .Z(n13033) );
  NAND U13866 ( .A(n13031), .B(n13030), .Z(n13032) );
  NAND U13867 ( .A(n13033), .B(n13032), .Z(n13043) );
  XNOR U13868 ( .A(n13042), .B(n13043), .Z(n13044) );
  XOR U13869 ( .A(n13045), .B(n13044), .Z(n13041) );
  OR U13870 ( .A(n13034), .B(sreg[1537]), .Z(n13038) );
  NANDN U13871 ( .A(n13036), .B(n13035), .Z(n13037) );
  AND U13872 ( .A(n13038), .B(n13037), .Z(n13040) );
  XNOR U13873 ( .A(sreg[1538]), .B(n13040), .Z(n13039) );
  XNOR U13874 ( .A(n13041), .B(n13039), .Z(c[1538]) );
  NANDN U13875 ( .A(n13043), .B(n13042), .Z(n13047) );
  NANDN U13876 ( .A(n13045), .B(n13044), .Z(n13046) );
  NAND U13877 ( .A(n13047), .B(n13046), .Z(n13063) );
  AND U13878 ( .A(b[2]), .B(a[517]), .Z(n13069) );
  AND U13879 ( .A(a[518]), .B(b[1]), .Z(n13067) );
  AND U13880 ( .A(a[516]), .B(b[3]), .Z(n13066) );
  XOR U13881 ( .A(n13067), .B(n13066), .Z(n13068) );
  XOR U13882 ( .A(n13069), .B(n13068), .Z(n13072) );
  NAND U13883 ( .A(b[0]), .B(a[519]), .Z(n13073) );
  XOR U13884 ( .A(n13072), .B(n13073), .Z(n13075) );
  OR U13885 ( .A(n13049), .B(n13048), .Z(n13053) );
  NANDN U13886 ( .A(n13051), .B(n13050), .Z(n13052) );
  NAND U13887 ( .A(n13053), .B(n13052), .Z(n13074) );
  XNOR U13888 ( .A(n13075), .B(n13074), .Z(n13060) );
  NANDN U13889 ( .A(n13055), .B(n13054), .Z(n13059) );
  OR U13890 ( .A(n13057), .B(n13056), .Z(n13058) );
  NAND U13891 ( .A(n13059), .B(n13058), .Z(n13061) );
  XNOR U13892 ( .A(n13060), .B(n13061), .Z(n13062) );
  XNOR U13893 ( .A(n13063), .B(n13062), .Z(n13078) );
  XNOR U13894 ( .A(n13078), .B(sreg[1539]), .Z(n13079) );
  XOR U13895 ( .A(n13080), .B(n13079), .Z(c[1539]) );
  NANDN U13896 ( .A(n13061), .B(n13060), .Z(n13065) );
  NAND U13897 ( .A(n13063), .B(n13062), .Z(n13064) );
  NAND U13898 ( .A(n13065), .B(n13064), .Z(n13091) );
  AND U13899 ( .A(b[2]), .B(a[518]), .Z(n13097) );
  AND U13900 ( .A(a[519]), .B(b[1]), .Z(n13095) );
  AND U13901 ( .A(a[517]), .B(b[3]), .Z(n13094) );
  XOR U13902 ( .A(n13095), .B(n13094), .Z(n13096) );
  XOR U13903 ( .A(n13097), .B(n13096), .Z(n13100) );
  NAND U13904 ( .A(b[0]), .B(a[520]), .Z(n13101) );
  XOR U13905 ( .A(n13100), .B(n13101), .Z(n13103) );
  OR U13906 ( .A(n13067), .B(n13066), .Z(n13071) );
  NANDN U13907 ( .A(n13069), .B(n13068), .Z(n13070) );
  NAND U13908 ( .A(n13071), .B(n13070), .Z(n13102) );
  XNOR U13909 ( .A(n13103), .B(n13102), .Z(n13088) );
  NANDN U13910 ( .A(n13073), .B(n13072), .Z(n13077) );
  OR U13911 ( .A(n13075), .B(n13074), .Z(n13076) );
  NAND U13912 ( .A(n13077), .B(n13076), .Z(n13089) );
  XNOR U13913 ( .A(n13088), .B(n13089), .Z(n13090) );
  XNOR U13914 ( .A(n13091), .B(n13090), .Z(n13083) );
  XOR U13915 ( .A(sreg[1540]), .B(n13083), .Z(n13084) );
  NAND U13916 ( .A(n13078), .B(sreg[1539]), .Z(n13082) );
  OR U13917 ( .A(n13080), .B(n13079), .Z(n13081) );
  NAND U13918 ( .A(n13082), .B(n13081), .Z(n13085) );
  XOR U13919 ( .A(n13084), .B(n13085), .Z(c[1540]) );
  OR U13920 ( .A(n13083), .B(sreg[1540]), .Z(n13087) );
  NANDN U13921 ( .A(n13085), .B(n13084), .Z(n13086) );
  AND U13922 ( .A(n13087), .B(n13086), .Z(n13125) );
  NANDN U13923 ( .A(n13089), .B(n13088), .Z(n13093) );
  NAND U13924 ( .A(n13091), .B(n13090), .Z(n13092) );
  NAND U13925 ( .A(n13093), .B(n13092), .Z(n13110) );
  AND U13926 ( .A(b[2]), .B(a[519]), .Z(n13116) );
  AND U13927 ( .A(a[520]), .B(b[1]), .Z(n13114) );
  AND U13928 ( .A(a[518]), .B(b[3]), .Z(n13113) );
  XOR U13929 ( .A(n13114), .B(n13113), .Z(n13115) );
  XOR U13930 ( .A(n13116), .B(n13115), .Z(n13119) );
  NAND U13931 ( .A(b[0]), .B(a[521]), .Z(n13120) );
  XOR U13932 ( .A(n13119), .B(n13120), .Z(n13122) );
  OR U13933 ( .A(n13095), .B(n13094), .Z(n13099) );
  NANDN U13934 ( .A(n13097), .B(n13096), .Z(n13098) );
  NAND U13935 ( .A(n13099), .B(n13098), .Z(n13121) );
  XNOR U13936 ( .A(n13122), .B(n13121), .Z(n13107) );
  NANDN U13937 ( .A(n13101), .B(n13100), .Z(n13105) );
  OR U13938 ( .A(n13103), .B(n13102), .Z(n13104) );
  NAND U13939 ( .A(n13105), .B(n13104), .Z(n13108) );
  XNOR U13940 ( .A(n13107), .B(n13108), .Z(n13109) );
  XNOR U13941 ( .A(n13110), .B(n13109), .Z(n13126) );
  XOR U13942 ( .A(sreg[1541]), .B(n13126), .Z(n13106) );
  XOR U13943 ( .A(n13125), .B(n13106), .Z(c[1541]) );
  NANDN U13944 ( .A(n13108), .B(n13107), .Z(n13112) );
  NAND U13945 ( .A(n13110), .B(n13109), .Z(n13111) );
  NAND U13946 ( .A(n13112), .B(n13111), .Z(n13133) );
  AND U13947 ( .A(b[2]), .B(a[520]), .Z(n13139) );
  AND U13948 ( .A(a[521]), .B(b[1]), .Z(n13137) );
  AND U13949 ( .A(a[519]), .B(b[3]), .Z(n13136) );
  XOR U13950 ( .A(n13137), .B(n13136), .Z(n13138) );
  XOR U13951 ( .A(n13139), .B(n13138), .Z(n13142) );
  NAND U13952 ( .A(b[0]), .B(a[522]), .Z(n13143) );
  XOR U13953 ( .A(n13142), .B(n13143), .Z(n13145) );
  OR U13954 ( .A(n13114), .B(n13113), .Z(n13118) );
  NANDN U13955 ( .A(n13116), .B(n13115), .Z(n13117) );
  NAND U13956 ( .A(n13118), .B(n13117), .Z(n13144) );
  XNOR U13957 ( .A(n13145), .B(n13144), .Z(n13130) );
  NANDN U13958 ( .A(n13120), .B(n13119), .Z(n13124) );
  OR U13959 ( .A(n13122), .B(n13121), .Z(n13123) );
  NAND U13960 ( .A(n13124), .B(n13123), .Z(n13131) );
  XNOR U13961 ( .A(n13130), .B(n13131), .Z(n13132) );
  XOR U13962 ( .A(n13133), .B(n13132), .Z(n13128) );
  XNOR U13963 ( .A(sreg[1542]), .B(n13129), .Z(n13127) );
  XOR U13964 ( .A(n13128), .B(n13127), .Z(c[1542]) );
  NANDN U13965 ( .A(n13131), .B(n13130), .Z(n13135) );
  NAND U13966 ( .A(n13133), .B(n13132), .Z(n13134) );
  NAND U13967 ( .A(n13135), .B(n13134), .Z(n13151) );
  AND U13968 ( .A(b[2]), .B(a[521]), .Z(n13157) );
  AND U13969 ( .A(a[522]), .B(b[1]), .Z(n13155) );
  AND U13970 ( .A(a[520]), .B(b[3]), .Z(n13154) );
  XOR U13971 ( .A(n13155), .B(n13154), .Z(n13156) );
  XOR U13972 ( .A(n13157), .B(n13156), .Z(n13160) );
  NAND U13973 ( .A(b[0]), .B(a[523]), .Z(n13161) );
  XOR U13974 ( .A(n13160), .B(n13161), .Z(n13163) );
  OR U13975 ( .A(n13137), .B(n13136), .Z(n13141) );
  NANDN U13976 ( .A(n13139), .B(n13138), .Z(n13140) );
  NAND U13977 ( .A(n13141), .B(n13140), .Z(n13162) );
  XNOR U13978 ( .A(n13163), .B(n13162), .Z(n13148) );
  NANDN U13979 ( .A(n13143), .B(n13142), .Z(n13147) );
  OR U13980 ( .A(n13145), .B(n13144), .Z(n13146) );
  NAND U13981 ( .A(n13147), .B(n13146), .Z(n13149) );
  XNOR U13982 ( .A(n13148), .B(n13149), .Z(n13150) );
  XNOR U13983 ( .A(n13151), .B(n13150), .Z(n13166) );
  XNOR U13984 ( .A(n13166), .B(sreg[1543]), .Z(n13167) );
  XOR U13985 ( .A(n13168), .B(n13167), .Z(c[1543]) );
  NANDN U13986 ( .A(n13149), .B(n13148), .Z(n13153) );
  NAND U13987 ( .A(n13151), .B(n13150), .Z(n13152) );
  NAND U13988 ( .A(n13153), .B(n13152), .Z(n13174) );
  AND U13989 ( .A(b[2]), .B(a[522]), .Z(n13180) );
  AND U13990 ( .A(a[523]), .B(b[1]), .Z(n13178) );
  AND U13991 ( .A(a[521]), .B(b[3]), .Z(n13177) );
  XOR U13992 ( .A(n13178), .B(n13177), .Z(n13179) );
  XOR U13993 ( .A(n13180), .B(n13179), .Z(n13183) );
  NAND U13994 ( .A(b[0]), .B(a[524]), .Z(n13184) );
  XOR U13995 ( .A(n13183), .B(n13184), .Z(n13186) );
  OR U13996 ( .A(n13155), .B(n13154), .Z(n13159) );
  NANDN U13997 ( .A(n13157), .B(n13156), .Z(n13158) );
  NAND U13998 ( .A(n13159), .B(n13158), .Z(n13185) );
  XNOR U13999 ( .A(n13186), .B(n13185), .Z(n13171) );
  NANDN U14000 ( .A(n13161), .B(n13160), .Z(n13165) );
  OR U14001 ( .A(n13163), .B(n13162), .Z(n13164) );
  NAND U14002 ( .A(n13165), .B(n13164), .Z(n13172) );
  XNOR U14003 ( .A(n13171), .B(n13172), .Z(n13173) );
  XNOR U14004 ( .A(n13174), .B(n13173), .Z(n13189) );
  XOR U14005 ( .A(sreg[1544]), .B(n13189), .Z(n13190) );
  NAND U14006 ( .A(n13166), .B(sreg[1543]), .Z(n13170) );
  OR U14007 ( .A(n13168), .B(n13167), .Z(n13169) );
  NAND U14008 ( .A(n13170), .B(n13169), .Z(n13191) );
  XOR U14009 ( .A(n13190), .B(n13191), .Z(c[1544]) );
  NANDN U14010 ( .A(n13172), .B(n13171), .Z(n13176) );
  NAND U14011 ( .A(n13174), .B(n13173), .Z(n13175) );
  NAND U14012 ( .A(n13176), .B(n13175), .Z(n13200) );
  AND U14013 ( .A(b[2]), .B(a[523]), .Z(n13206) );
  AND U14014 ( .A(a[524]), .B(b[1]), .Z(n13204) );
  AND U14015 ( .A(a[522]), .B(b[3]), .Z(n13203) );
  XOR U14016 ( .A(n13204), .B(n13203), .Z(n13205) );
  XOR U14017 ( .A(n13206), .B(n13205), .Z(n13209) );
  NAND U14018 ( .A(b[0]), .B(a[525]), .Z(n13210) );
  XOR U14019 ( .A(n13209), .B(n13210), .Z(n13212) );
  OR U14020 ( .A(n13178), .B(n13177), .Z(n13182) );
  NANDN U14021 ( .A(n13180), .B(n13179), .Z(n13181) );
  NAND U14022 ( .A(n13182), .B(n13181), .Z(n13211) );
  XNOR U14023 ( .A(n13212), .B(n13211), .Z(n13197) );
  NANDN U14024 ( .A(n13184), .B(n13183), .Z(n13188) );
  OR U14025 ( .A(n13186), .B(n13185), .Z(n13187) );
  NAND U14026 ( .A(n13188), .B(n13187), .Z(n13198) );
  XNOR U14027 ( .A(n13197), .B(n13198), .Z(n13199) );
  XOR U14028 ( .A(n13200), .B(n13199), .Z(n13196) );
  OR U14029 ( .A(n13189), .B(sreg[1544]), .Z(n13193) );
  NANDN U14030 ( .A(n13191), .B(n13190), .Z(n13192) );
  AND U14031 ( .A(n13193), .B(n13192), .Z(n13195) );
  XNOR U14032 ( .A(sreg[1545]), .B(n13195), .Z(n13194) );
  XOR U14033 ( .A(n13196), .B(n13194), .Z(c[1545]) );
  NANDN U14034 ( .A(n13198), .B(n13197), .Z(n13202) );
  NAND U14035 ( .A(n13200), .B(n13199), .Z(n13201) );
  NAND U14036 ( .A(n13202), .B(n13201), .Z(n13218) );
  AND U14037 ( .A(b[2]), .B(a[524]), .Z(n13224) );
  AND U14038 ( .A(a[525]), .B(b[1]), .Z(n13222) );
  AND U14039 ( .A(a[523]), .B(b[3]), .Z(n13221) );
  XOR U14040 ( .A(n13222), .B(n13221), .Z(n13223) );
  XOR U14041 ( .A(n13224), .B(n13223), .Z(n13227) );
  NAND U14042 ( .A(b[0]), .B(a[526]), .Z(n13228) );
  XOR U14043 ( .A(n13227), .B(n13228), .Z(n13230) );
  OR U14044 ( .A(n13204), .B(n13203), .Z(n13208) );
  NANDN U14045 ( .A(n13206), .B(n13205), .Z(n13207) );
  NAND U14046 ( .A(n13208), .B(n13207), .Z(n13229) );
  XNOR U14047 ( .A(n13230), .B(n13229), .Z(n13215) );
  NANDN U14048 ( .A(n13210), .B(n13209), .Z(n13214) );
  OR U14049 ( .A(n13212), .B(n13211), .Z(n13213) );
  NAND U14050 ( .A(n13214), .B(n13213), .Z(n13216) );
  XNOR U14051 ( .A(n13215), .B(n13216), .Z(n13217) );
  XNOR U14052 ( .A(n13218), .B(n13217), .Z(n13233) );
  XNOR U14053 ( .A(n13233), .B(sreg[1546]), .Z(n13234) );
  XOR U14054 ( .A(n13235), .B(n13234), .Z(c[1546]) );
  NANDN U14055 ( .A(n13216), .B(n13215), .Z(n13220) );
  NAND U14056 ( .A(n13218), .B(n13217), .Z(n13219) );
  NAND U14057 ( .A(n13220), .B(n13219), .Z(n13244) );
  AND U14058 ( .A(b[2]), .B(a[525]), .Z(n13250) );
  AND U14059 ( .A(a[526]), .B(b[1]), .Z(n13248) );
  AND U14060 ( .A(a[524]), .B(b[3]), .Z(n13247) );
  XOR U14061 ( .A(n13248), .B(n13247), .Z(n13249) );
  XOR U14062 ( .A(n13250), .B(n13249), .Z(n13253) );
  NAND U14063 ( .A(b[0]), .B(a[527]), .Z(n13254) );
  XOR U14064 ( .A(n13253), .B(n13254), .Z(n13256) );
  OR U14065 ( .A(n13222), .B(n13221), .Z(n13226) );
  NANDN U14066 ( .A(n13224), .B(n13223), .Z(n13225) );
  NAND U14067 ( .A(n13226), .B(n13225), .Z(n13255) );
  XNOR U14068 ( .A(n13256), .B(n13255), .Z(n13241) );
  NANDN U14069 ( .A(n13228), .B(n13227), .Z(n13232) );
  OR U14070 ( .A(n13230), .B(n13229), .Z(n13231) );
  NAND U14071 ( .A(n13232), .B(n13231), .Z(n13242) );
  XNOR U14072 ( .A(n13241), .B(n13242), .Z(n13243) );
  XOR U14073 ( .A(n13244), .B(n13243), .Z(n13240) );
  NAND U14074 ( .A(n13233), .B(sreg[1546]), .Z(n13237) );
  OR U14075 ( .A(n13235), .B(n13234), .Z(n13236) );
  NAND U14076 ( .A(n13237), .B(n13236), .Z(n13239) );
  XNOR U14077 ( .A(sreg[1547]), .B(n13239), .Z(n13238) );
  XOR U14078 ( .A(n13240), .B(n13238), .Z(c[1547]) );
  NANDN U14079 ( .A(n13242), .B(n13241), .Z(n13246) );
  NAND U14080 ( .A(n13244), .B(n13243), .Z(n13245) );
  NAND U14081 ( .A(n13246), .B(n13245), .Z(n13262) );
  AND U14082 ( .A(b[2]), .B(a[526]), .Z(n13268) );
  AND U14083 ( .A(a[527]), .B(b[1]), .Z(n13266) );
  AND U14084 ( .A(a[525]), .B(b[3]), .Z(n13265) );
  XOR U14085 ( .A(n13266), .B(n13265), .Z(n13267) );
  XOR U14086 ( .A(n13268), .B(n13267), .Z(n13271) );
  NAND U14087 ( .A(b[0]), .B(a[528]), .Z(n13272) );
  XOR U14088 ( .A(n13271), .B(n13272), .Z(n13274) );
  OR U14089 ( .A(n13248), .B(n13247), .Z(n13252) );
  NANDN U14090 ( .A(n13250), .B(n13249), .Z(n13251) );
  NAND U14091 ( .A(n13252), .B(n13251), .Z(n13273) );
  XNOR U14092 ( .A(n13274), .B(n13273), .Z(n13259) );
  NANDN U14093 ( .A(n13254), .B(n13253), .Z(n13258) );
  OR U14094 ( .A(n13256), .B(n13255), .Z(n13257) );
  NAND U14095 ( .A(n13258), .B(n13257), .Z(n13260) );
  XNOR U14096 ( .A(n13259), .B(n13260), .Z(n13261) );
  XNOR U14097 ( .A(n13262), .B(n13261), .Z(n13277) );
  XNOR U14098 ( .A(n13277), .B(sreg[1548]), .Z(n13278) );
  XOR U14099 ( .A(n13279), .B(n13278), .Z(c[1548]) );
  NANDN U14100 ( .A(n13260), .B(n13259), .Z(n13264) );
  NAND U14101 ( .A(n13262), .B(n13261), .Z(n13263) );
  NAND U14102 ( .A(n13264), .B(n13263), .Z(n13285) );
  AND U14103 ( .A(b[2]), .B(a[527]), .Z(n13291) );
  AND U14104 ( .A(a[528]), .B(b[1]), .Z(n13289) );
  AND U14105 ( .A(a[526]), .B(b[3]), .Z(n13288) );
  XOR U14106 ( .A(n13289), .B(n13288), .Z(n13290) );
  XOR U14107 ( .A(n13291), .B(n13290), .Z(n13294) );
  NAND U14108 ( .A(b[0]), .B(a[529]), .Z(n13295) );
  XOR U14109 ( .A(n13294), .B(n13295), .Z(n13297) );
  OR U14110 ( .A(n13266), .B(n13265), .Z(n13270) );
  NANDN U14111 ( .A(n13268), .B(n13267), .Z(n13269) );
  NAND U14112 ( .A(n13270), .B(n13269), .Z(n13296) );
  XNOR U14113 ( .A(n13297), .B(n13296), .Z(n13282) );
  NANDN U14114 ( .A(n13272), .B(n13271), .Z(n13276) );
  OR U14115 ( .A(n13274), .B(n13273), .Z(n13275) );
  NAND U14116 ( .A(n13276), .B(n13275), .Z(n13283) );
  XNOR U14117 ( .A(n13282), .B(n13283), .Z(n13284) );
  XNOR U14118 ( .A(n13285), .B(n13284), .Z(n13300) );
  XNOR U14119 ( .A(n13300), .B(sreg[1549]), .Z(n13302) );
  NAND U14120 ( .A(n13277), .B(sreg[1548]), .Z(n13281) );
  OR U14121 ( .A(n13279), .B(n13278), .Z(n13280) );
  AND U14122 ( .A(n13281), .B(n13280), .Z(n13301) );
  XOR U14123 ( .A(n13302), .B(n13301), .Z(c[1549]) );
  NANDN U14124 ( .A(n13283), .B(n13282), .Z(n13287) );
  NAND U14125 ( .A(n13285), .B(n13284), .Z(n13286) );
  NAND U14126 ( .A(n13287), .B(n13286), .Z(n13309) );
  AND U14127 ( .A(b[2]), .B(a[528]), .Z(n13315) );
  AND U14128 ( .A(a[529]), .B(b[1]), .Z(n13313) );
  AND U14129 ( .A(a[527]), .B(b[3]), .Z(n13312) );
  XOR U14130 ( .A(n13313), .B(n13312), .Z(n13314) );
  XOR U14131 ( .A(n13315), .B(n13314), .Z(n13318) );
  NAND U14132 ( .A(b[0]), .B(a[530]), .Z(n13319) );
  XOR U14133 ( .A(n13318), .B(n13319), .Z(n13321) );
  OR U14134 ( .A(n13289), .B(n13288), .Z(n13293) );
  NANDN U14135 ( .A(n13291), .B(n13290), .Z(n13292) );
  NAND U14136 ( .A(n13293), .B(n13292), .Z(n13320) );
  XNOR U14137 ( .A(n13321), .B(n13320), .Z(n13306) );
  NANDN U14138 ( .A(n13295), .B(n13294), .Z(n13299) );
  OR U14139 ( .A(n13297), .B(n13296), .Z(n13298) );
  NAND U14140 ( .A(n13299), .B(n13298), .Z(n13307) );
  XNOR U14141 ( .A(n13306), .B(n13307), .Z(n13308) );
  XOR U14142 ( .A(n13309), .B(n13308), .Z(n13325) );
  NAND U14143 ( .A(n13300), .B(sreg[1549]), .Z(n13304) );
  OR U14144 ( .A(n13302), .B(n13301), .Z(n13303) );
  NAND U14145 ( .A(n13304), .B(n13303), .Z(n13324) );
  XNOR U14146 ( .A(sreg[1550]), .B(n13324), .Z(n13305) );
  XOR U14147 ( .A(n13325), .B(n13305), .Z(c[1550]) );
  NANDN U14148 ( .A(n13307), .B(n13306), .Z(n13311) );
  NAND U14149 ( .A(n13309), .B(n13308), .Z(n13310) );
  NAND U14150 ( .A(n13311), .B(n13310), .Z(n13330) );
  AND U14151 ( .A(b[2]), .B(a[529]), .Z(n13336) );
  AND U14152 ( .A(a[530]), .B(b[1]), .Z(n13334) );
  AND U14153 ( .A(a[528]), .B(b[3]), .Z(n13333) );
  XOR U14154 ( .A(n13334), .B(n13333), .Z(n13335) );
  XOR U14155 ( .A(n13336), .B(n13335), .Z(n13339) );
  NAND U14156 ( .A(b[0]), .B(a[531]), .Z(n13340) );
  XOR U14157 ( .A(n13339), .B(n13340), .Z(n13342) );
  OR U14158 ( .A(n13313), .B(n13312), .Z(n13317) );
  NANDN U14159 ( .A(n13315), .B(n13314), .Z(n13316) );
  NAND U14160 ( .A(n13317), .B(n13316), .Z(n13341) );
  XNOR U14161 ( .A(n13342), .B(n13341), .Z(n13327) );
  NANDN U14162 ( .A(n13319), .B(n13318), .Z(n13323) );
  OR U14163 ( .A(n13321), .B(n13320), .Z(n13322) );
  NAND U14164 ( .A(n13323), .B(n13322), .Z(n13328) );
  XNOR U14165 ( .A(n13327), .B(n13328), .Z(n13329) );
  XOR U14166 ( .A(n13330), .B(n13329), .Z(n13346) );
  XNOR U14167 ( .A(sreg[1551]), .B(n13345), .Z(n13326) );
  XOR U14168 ( .A(n13346), .B(n13326), .Z(c[1551]) );
  NANDN U14169 ( .A(n13328), .B(n13327), .Z(n13332) );
  NAND U14170 ( .A(n13330), .B(n13329), .Z(n13331) );
  NAND U14171 ( .A(n13332), .B(n13331), .Z(n13353) );
  AND U14172 ( .A(b[2]), .B(a[530]), .Z(n13365) );
  AND U14173 ( .A(a[531]), .B(b[1]), .Z(n13363) );
  AND U14174 ( .A(a[529]), .B(b[3]), .Z(n13362) );
  XOR U14175 ( .A(n13363), .B(n13362), .Z(n13364) );
  XOR U14176 ( .A(n13365), .B(n13364), .Z(n13356) );
  NAND U14177 ( .A(b[0]), .B(a[532]), .Z(n13357) );
  XOR U14178 ( .A(n13356), .B(n13357), .Z(n13359) );
  OR U14179 ( .A(n13334), .B(n13333), .Z(n13338) );
  NANDN U14180 ( .A(n13336), .B(n13335), .Z(n13337) );
  NAND U14181 ( .A(n13338), .B(n13337), .Z(n13358) );
  XNOR U14182 ( .A(n13359), .B(n13358), .Z(n13350) );
  NANDN U14183 ( .A(n13340), .B(n13339), .Z(n13344) );
  OR U14184 ( .A(n13342), .B(n13341), .Z(n13343) );
  NAND U14185 ( .A(n13344), .B(n13343), .Z(n13351) );
  XNOR U14186 ( .A(n13350), .B(n13351), .Z(n13352) );
  XNOR U14187 ( .A(n13353), .B(n13352), .Z(n13349) );
  XOR U14188 ( .A(n13348), .B(sreg[1552]), .Z(n13347) );
  XOR U14189 ( .A(n13349), .B(n13347), .Z(c[1552]) );
  NANDN U14190 ( .A(n13351), .B(n13350), .Z(n13355) );
  NAND U14191 ( .A(n13353), .B(n13352), .Z(n13354) );
  NAND U14192 ( .A(n13355), .B(n13354), .Z(n13383) );
  NANDN U14193 ( .A(n13357), .B(n13356), .Z(n13361) );
  OR U14194 ( .A(n13359), .B(n13358), .Z(n13360) );
  NAND U14195 ( .A(n13361), .B(n13360), .Z(n13380) );
  AND U14196 ( .A(b[2]), .B(a[531]), .Z(n13371) );
  AND U14197 ( .A(a[532]), .B(b[1]), .Z(n13369) );
  AND U14198 ( .A(a[530]), .B(b[3]), .Z(n13368) );
  XOR U14199 ( .A(n13369), .B(n13368), .Z(n13370) );
  XOR U14200 ( .A(n13371), .B(n13370), .Z(n13374) );
  NAND U14201 ( .A(b[0]), .B(a[533]), .Z(n13375) );
  XNOR U14202 ( .A(n13374), .B(n13375), .Z(n13376) );
  OR U14203 ( .A(n13363), .B(n13362), .Z(n13367) );
  NANDN U14204 ( .A(n13365), .B(n13364), .Z(n13366) );
  AND U14205 ( .A(n13367), .B(n13366), .Z(n13377) );
  XNOR U14206 ( .A(n13376), .B(n13377), .Z(n13381) );
  XNOR U14207 ( .A(n13380), .B(n13381), .Z(n13382) );
  XNOR U14208 ( .A(n13383), .B(n13382), .Z(n13386) );
  XNOR U14209 ( .A(sreg[1553]), .B(n13386), .Z(n13388) );
  XNOR U14210 ( .A(n13387), .B(n13388), .Z(c[1553]) );
  AND U14211 ( .A(b[2]), .B(a[532]), .Z(n13403) );
  AND U14212 ( .A(a[533]), .B(b[1]), .Z(n13401) );
  AND U14213 ( .A(a[531]), .B(b[3]), .Z(n13400) );
  XOR U14214 ( .A(n13401), .B(n13400), .Z(n13402) );
  XOR U14215 ( .A(n13403), .B(n13402), .Z(n13406) );
  NAND U14216 ( .A(b[0]), .B(a[534]), .Z(n13407) );
  XOR U14217 ( .A(n13406), .B(n13407), .Z(n13409) );
  OR U14218 ( .A(n13369), .B(n13368), .Z(n13373) );
  NANDN U14219 ( .A(n13371), .B(n13370), .Z(n13372) );
  NAND U14220 ( .A(n13373), .B(n13372), .Z(n13408) );
  XNOR U14221 ( .A(n13409), .B(n13408), .Z(n13394) );
  NANDN U14222 ( .A(n13375), .B(n13374), .Z(n13379) );
  NAND U14223 ( .A(n13377), .B(n13376), .Z(n13378) );
  NAND U14224 ( .A(n13379), .B(n13378), .Z(n13395) );
  XNOR U14225 ( .A(n13394), .B(n13395), .Z(n13396) );
  NANDN U14226 ( .A(n13381), .B(n13380), .Z(n13385) );
  NANDN U14227 ( .A(n13383), .B(n13382), .Z(n13384) );
  AND U14228 ( .A(n13385), .B(n13384), .Z(n13397) );
  XNOR U14229 ( .A(n13396), .B(n13397), .Z(n13393) );
  NAND U14230 ( .A(sreg[1553]), .B(n13386), .Z(n13390) );
  NANDN U14231 ( .A(n13388), .B(n13387), .Z(n13389) );
  AND U14232 ( .A(n13390), .B(n13389), .Z(n13392) );
  XNOR U14233 ( .A(n13392), .B(sreg[1554]), .Z(n13391) );
  XOR U14234 ( .A(n13393), .B(n13391), .Z(c[1554]) );
  NANDN U14235 ( .A(n13395), .B(n13394), .Z(n13399) );
  NAND U14236 ( .A(n13397), .B(n13396), .Z(n13398) );
  NAND U14237 ( .A(n13399), .B(n13398), .Z(n13427) );
  AND U14238 ( .A(b[2]), .B(a[533]), .Z(n13421) );
  AND U14239 ( .A(a[534]), .B(b[1]), .Z(n13419) );
  AND U14240 ( .A(a[532]), .B(b[3]), .Z(n13418) );
  XOR U14241 ( .A(n13419), .B(n13418), .Z(n13420) );
  XOR U14242 ( .A(n13421), .B(n13420), .Z(n13412) );
  NAND U14243 ( .A(b[0]), .B(a[535]), .Z(n13413) );
  XOR U14244 ( .A(n13412), .B(n13413), .Z(n13415) );
  OR U14245 ( .A(n13401), .B(n13400), .Z(n13405) );
  NANDN U14246 ( .A(n13403), .B(n13402), .Z(n13404) );
  NAND U14247 ( .A(n13405), .B(n13404), .Z(n13414) );
  XNOR U14248 ( .A(n13415), .B(n13414), .Z(n13424) );
  NANDN U14249 ( .A(n13407), .B(n13406), .Z(n13411) );
  OR U14250 ( .A(n13409), .B(n13408), .Z(n13410) );
  NAND U14251 ( .A(n13411), .B(n13410), .Z(n13425) );
  XNOR U14252 ( .A(n13424), .B(n13425), .Z(n13426) );
  XNOR U14253 ( .A(n13427), .B(n13426), .Z(n13430) );
  XNOR U14254 ( .A(n13430), .B(sreg[1555]), .Z(n13432) );
  XNOR U14255 ( .A(n13431), .B(n13432), .Z(c[1555]) );
  NANDN U14256 ( .A(n13413), .B(n13412), .Z(n13417) );
  OR U14257 ( .A(n13415), .B(n13414), .Z(n13416) );
  NAND U14258 ( .A(n13417), .B(n13416), .Z(n13450) );
  AND U14259 ( .A(b[2]), .B(a[534]), .Z(n13441) );
  AND U14260 ( .A(a[535]), .B(b[1]), .Z(n13439) );
  AND U14261 ( .A(a[533]), .B(b[3]), .Z(n13438) );
  XOR U14262 ( .A(n13439), .B(n13438), .Z(n13440) );
  XOR U14263 ( .A(n13441), .B(n13440), .Z(n13444) );
  NAND U14264 ( .A(b[0]), .B(a[536]), .Z(n13445) );
  XNOR U14265 ( .A(n13444), .B(n13445), .Z(n13446) );
  OR U14266 ( .A(n13419), .B(n13418), .Z(n13423) );
  NANDN U14267 ( .A(n13421), .B(n13420), .Z(n13422) );
  AND U14268 ( .A(n13423), .B(n13422), .Z(n13447) );
  XNOR U14269 ( .A(n13446), .B(n13447), .Z(n13451) );
  XNOR U14270 ( .A(n13450), .B(n13451), .Z(n13452) );
  NANDN U14271 ( .A(n13425), .B(n13424), .Z(n13429) );
  NAND U14272 ( .A(n13427), .B(n13426), .Z(n13428) );
  NAND U14273 ( .A(n13429), .B(n13428), .Z(n13453) );
  XOR U14274 ( .A(n13452), .B(n13453), .Z(n13437) );
  NAND U14275 ( .A(n13430), .B(sreg[1555]), .Z(n13434) );
  NANDN U14276 ( .A(n13432), .B(n13431), .Z(n13433) );
  AND U14277 ( .A(n13434), .B(n13433), .Z(n13436) );
  XNOR U14278 ( .A(n13436), .B(sreg[1556]), .Z(n13435) );
  XNOR U14279 ( .A(n13437), .B(n13435), .Z(c[1556]) );
  AND U14280 ( .A(b[2]), .B(a[535]), .Z(n13465) );
  AND U14281 ( .A(a[536]), .B(b[1]), .Z(n13463) );
  AND U14282 ( .A(a[534]), .B(b[3]), .Z(n13462) );
  XOR U14283 ( .A(n13463), .B(n13462), .Z(n13464) );
  XOR U14284 ( .A(n13465), .B(n13464), .Z(n13468) );
  NAND U14285 ( .A(b[0]), .B(a[537]), .Z(n13469) );
  XOR U14286 ( .A(n13468), .B(n13469), .Z(n13471) );
  OR U14287 ( .A(n13439), .B(n13438), .Z(n13443) );
  NANDN U14288 ( .A(n13441), .B(n13440), .Z(n13442) );
  NAND U14289 ( .A(n13443), .B(n13442), .Z(n13470) );
  XNOR U14290 ( .A(n13471), .B(n13470), .Z(n13456) );
  NANDN U14291 ( .A(n13445), .B(n13444), .Z(n13449) );
  NAND U14292 ( .A(n13447), .B(n13446), .Z(n13448) );
  NAND U14293 ( .A(n13449), .B(n13448), .Z(n13457) );
  XNOR U14294 ( .A(n13456), .B(n13457), .Z(n13458) );
  NANDN U14295 ( .A(n13451), .B(n13450), .Z(n13455) );
  NANDN U14296 ( .A(n13453), .B(n13452), .Z(n13454) );
  NAND U14297 ( .A(n13455), .B(n13454), .Z(n13459) );
  XOR U14298 ( .A(n13458), .B(n13459), .Z(n13474) );
  XNOR U14299 ( .A(n13474), .B(sreg[1557]), .Z(n13476) );
  XNOR U14300 ( .A(n13475), .B(n13476), .Z(c[1557]) );
  NANDN U14301 ( .A(n13457), .B(n13456), .Z(n13461) );
  NANDN U14302 ( .A(n13459), .B(n13458), .Z(n13460) );
  NAND U14303 ( .A(n13461), .B(n13460), .Z(n13482) );
  AND U14304 ( .A(b[2]), .B(a[536]), .Z(n13488) );
  AND U14305 ( .A(a[537]), .B(b[1]), .Z(n13486) );
  AND U14306 ( .A(a[535]), .B(b[3]), .Z(n13485) );
  XOR U14307 ( .A(n13486), .B(n13485), .Z(n13487) );
  XOR U14308 ( .A(n13488), .B(n13487), .Z(n13491) );
  NAND U14309 ( .A(b[0]), .B(a[538]), .Z(n13492) );
  XOR U14310 ( .A(n13491), .B(n13492), .Z(n13494) );
  OR U14311 ( .A(n13463), .B(n13462), .Z(n13467) );
  NANDN U14312 ( .A(n13465), .B(n13464), .Z(n13466) );
  NAND U14313 ( .A(n13467), .B(n13466), .Z(n13493) );
  XNOR U14314 ( .A(n13494), .B(n13493), .Z(n13479) );
  NANDN U14315 ( .A(n13469), .B(n13468), .Z(n13473) );
  OR U14316 ( .A(n13471), .B(n13470), .Z(n13472) );
  NAND U14317 ( .A(n13473), .B(n13472), .Z(n13480) );
  XNOR U14318 ( .A(n13479), .B(n13480), .Z(n13481) );
  XNOR U14319 ( .A(n13482), .B(n13481), .Z(n13497) );
  XOR U14320 ( .A(sreg[1558]), .B(n13497), .Z(n13498) );
  NAND U14321 ( .A(n13474), .B(sreg[1557]), .Z(n13478) );
  NANDN U14322 ( .A(n13476), .B(n13475), .Z(n13477) );
  NAND U14323 ( .A(n13478), .B(n13477), .Z(n13499) );
  XOR U14324 ( .A(n13498), .B(n13499), .Z(c[1558]) );
  NANDN U14325 ( .A(n13480), .B(n13479), .Z(n13484) );
  NAND U14326 ( .A(n13482), .B(n13481), .Z(n13483) );
  NAND U14327 ( .A(n13484), .B(n13483), .Z(n13506) );
  AND U14328 ( .A(b[2]), .B(a[537]), .Z(n13512) );
  AND U14329 ( .A(a[538]), .B(b[1]), .Z(n13510) );
  AND U14330 ( .A(a[536]), .B(b[3]), .Z(n13509) );
  XOR U14331 ( .A(n13510), .B(n13509), .Z(n13511) );
  XOR U14332 ( .A(n13512), .B(n13511), .Z(n13515) );
  NAND U14333 ( .A(b[0]), .B(a[539]), .Z(n13516) );
  XOR U14334 ( .A(n13515), .B(n13516), .Z(n13518) );
  OR U14335 ( .A(n13486), .B(n13485), .Z(n13490) );
  NANDN U14336 ( .A(n13488), .B(n13487), .Z(n13489) );
  NAND U14337 ( .A(n13490), .B(n13489), .Z(n13517) );
  XNOR U14338 ( .A(n13518), .B(n13517), .Z(n13503) );
  NANDN U14339 ( .A(n13492), .B(n13491), .Z(n13496) );
  OR U14340 ( .A(n13494), .B(n13493), .Z(n13495) );
  NAND U14341 ( .A(n13496), .B(n13495), .Z(n13504) );
  XNOR U14342 ( .A(n13503), .B(n13504), .Z(n13505) );
  XOR U14343 ( .A(n13506), .B(n13505), .Z(n13522) );
  OR U14344 ( .A(n13497), .B(sreg[1558]), .Z(n13501) );
  NANDN U14345 ( .A(n13499), .B(n13498), .Z(n13500) );
  AND U14346 ( .A(n13501), .B(n13500), .Z(n13521) );
  XNOR U14347 ( .A(sreg[1559]), .B(n13521), .Z(n13502) );
  XOR U14348 ( .A(n13522), .B(n13502), .Z(c[1559]) );
  NANDN U14349 ( .A(n13504), .B(n13503), .Z(n13508) );
  NAND U14350 ( .A(n13506), .B(n13505), .Z(n13507) );
  NAND U14351 ( .A(n13508), .B(n13507), .Z(n13527) );
  AND U14352 ( .A(b[2]), .B(a[538]), .Z(n13533) );
  AND U14353 ( .A(a[539]), .B(b[1]), .Z(n13531) );
  AND U14354 ( .A(a[537]), .B(b[3]), .Z(n13530) );
  XOR U14355 ( .A(n13531), .B(n13530), .Z(n13532) );
  XOR U14356 ( .A(n13533), .B(n13532), .Z(n13536) );
  NAND U14357 ( .A(b[0]), .B(a[540]), .Z(n13537) );
  XOR U14358 ( .A(n13536), .B(n13537), .Z(n13539) );
  OR U14359 ( .A(n13510), .B(n13509), .Z(n13514) );
  NANDN U14360 ( .A(n13512), .B(n13511), .Z(n13513) );
  NAND U14361 ( .A(n13514), .B(n13513), .Z(n13538) );
  XNOR U14362 ( .A(n13539), .B(n13538), .Z(n13524) );
  NANDN U14363 ( .A(n13516), .B(n13515), .Z(n13520) );
  OR U14364 ( .A(n13518), .B(n13517), .Z(n13519) );
  NAND U14365 ( .A(n13520), .B(n13519), .Z(n13525) );
  XNOR U14366 ( .A(n13524), .B(n13525), .Z(n13526) );
  XOR U14367 ( .A(n13527), .B(n13526), .Z(n13543) );
  XNOR U14368 ( .A(sreg[1560]), .B(n13542), .Z(n13523) );
  XOR U14369 ( .A(n13543), .B(n13523), .Z(c[1560]) );
  NANDN U14370 ( .A(n13525), .B(n13524), .Z(n13529) );
  NAND U14371 ( .A(n13527), .B(n13526), .Z(n13528) );
  NAND U14372 ( .A(n13529), .B(n13528), .Z(n13550) );
  AND U14373 ( .A(b[2]), .B(a[539]), .Z(n13556) );
  AND U14374 ( .A(a[540]), .B(b[1]), .Z(n13554) );
  AND U14375 ( .A(a[538]), .B(b[3]), .Z(n13553) );
  XOR U14376 ( .A(n13554), .B(n13553), .Z(n13555) );
  XOR U14377 ( .A(n13556), .B(n13555), .Z(n13559) );
  NAND U14378 ( .A(b[0]), .B(a[541]), .Z(n13560) );
  XOR U14379 ( .A(n13559), .B(n13560), .Z(n13562) );
  OR U14380 ( .A(n13531), .B(n13530), .Z(n13535) );
  NANDN U14381 ( .A(n13533), .B(n13532), .Z(n13534) );
  NAND U14382 ( .A(n13535), .B(n13534), .Z(n13561) );
  XNOR U14383 ( .A(n13562), .B(n13561), .Z(n13547) );
  NANDN U14384 ( .A(n13537), .B(n13536), .Z(n13541) );
  OR U14385 ( .A(n13539), .B(n13538), .Z(n13540) );
  NAND U14386 ( .A(n13541), .B(n13540), .Z(n13548) );
  XNOR U14387 ( .A(n13547), .B(n13548), .Z(n13549) );
  XOR U14388 ( .A(n13550), .B(n13549), .Z(n13546) );
  XNOR U14389 ( .A(sreg[1561]), .B(n13545), .Z(n13544) );
  XOR U14390 ( .A(n13546), .B(n13544), .Z(c[1561]) );
  NANDN U14391 ( .A(n13548), .B(n13547), .Z(n13552) );
  NAND U14392 ( .A(n13550), .B(n13549), .Z(n13551) );
  NAND U14393 ( .A(n13552), .B(n13551), .Z(n13568) );
  AND U14394 ( .A(b[2]), .B(a[540]), .Z(n13574) );
  AND U14395 ( .A(a[541]), .B(b[1]), .Z(n13572) );
  AND U14396 ( .A(a[539]), .B(b[3]), .Z(n13571) );
  XOR U14397 ( .A(n13572), .B(n13571), .Z(n13573) );
  XOR U14398 ( .A(n13574), .B(n13573), .Z(n13577) );
  NAND U14399 ( .A(b[0]), .B(a[542]), .Z(n13578) );
  XOR U14400 ( .A(n13577), .B(n13578), .Z(n13580) );
  OR U14401 ( .A(n13554), .B(n13553), .Z(n13558) );
  NANDN U14402 ( .A(n13556), .B(n13555), .Z(n13557) );
  NAND U14403 ( .A(n13558), .B(n13557), .Z(n13579) );
  XNOR U14404 ( .A(n13580), .B(n13579), .Z(n13565) );
  NANDN U14405 ( .A(n13560), .B(n13559), .Z(n13564) );
  OR U14406 ( .A(n13562), .B(n13561), .Z(n13563) );
  NAND U14407 ( .A(n13564), .B(n13563), .Z(n13566) );
  XNOR U14408 ( .A(n13565), .B(n13566), .Z(n13567) );
  XNOR U14409 ( .A(n13568), .B(n13567), .Z(n13583) );
  XNOR U14410 ( .A(n13583), .B(sreg[1562]), .Z(n13584) );
  XOR U14411 ( .A(n13585), .B(n13584), .Z(c[1562]) );
  NANDN U14412 ( .A(n13566), .B(n13565), .Z(n13570) );
  NAND U14413 ( .A(n13568), .B(n13567), .Z(n13569) );
  NAND U14414 ( .A(n13570), .B(n13569), .Z(n13596) );
  AND U14415 ( .A(b[2]), .B(a[541]), .Z(n13602) );
  AND U14416 ( .A(a[542]), .B(b[1]), .Z(n13600) );
  AND U14417 ( .A(a[540]), .B(b[3]), .Z(n13599) );
  XOR U14418 ( .A(n13600), .B(n13599), .Z(n13601) );
  XOR U14419 ( .A(n13602), .B(n13601), .Z(n13605) );
  NAND U14420 ( .A(b[0]), .B(a[543]), .Z(n13606) );
  XOR U14421 ( .A(n13605), .B(n13606), .Z(n13608) );
  OR U14422 ( .A(n13572), .B(n13571), .Z(n13576) );
  NANDN U14423 ( .A(n13574), .B(n13573), .Z(n13575) );
  NAND U14424 ( .A(n13576), .B(n13575), .Z(n13607) );
  XNOR U14425 ( .A(n13608), .B(n13607), .Z(n13593) );
  NANDN U14426 ( .A(n13578), .B(n13577), .Z(n13582) );
  OR U14427 ( .A(n13580), .B(n13579), .Z(n13581) );
  NAND U14428 ( .A(n13582), .B(n13581), .Z(n13594) );
  XNOR U14429 ( .A(n13593), .B(n13594), .Z(n13595) );
  XNOR U14430 ( .A(n13596), .B(n13595), .Z(n13588) );
  XOR U14431 ( .A(sreg[1563]), .B(n13588), .Z(n13589) );
  NAND U14432 ( .A(n13583), .B(sreg[1562]), .Z(n13587) );
  OR U14433 ( .A(n13585), .B(n13584), .Z(n13586) );
  NAND U14434 ( .A(n13587), .B(n13586), .Z(n13590) );
  XOR U14435 ( .A(n13589), .B(n13590), .Z(c[1563]) );
  OR U14436 ( .A(n13588), .B(sreg[1563]), .Z(n13592) );
  NANDN U14437 ( .A(n13590), .B(n13589), .Z(n13591) );
  NAND U14438 ( .A(n13592), .B(n13591), .Z(n13631) );
  NANDN U14439 ( .A(n13594), .B(n13593), .Z(n13598) );
  NAND U14440 ( .A(n13596), .B(n13595), .Z(n13597) );
  NAND U14441 ( .A(n13598), .B(n13597), .Z(n13614) );
  AND U14442 ( .A(b[2]), .B(a[542]), .Z(n13620) );
  AND U14443 ( .A(a[543]), .B(b[1]), .Z(n13618) );
  AND U14444 ( .A(a[541]), .B(b[3]), .Z(n13617) );
  XOR U14445 ( .A(n13618), .B(n13617), .Z(n13619) );
  XOR U14446 ( .A(n13620), .B(n13619), .Z(n13623) );
  NAND U14447 ( .A(b[0]), .B(a[544]), .Z(n13624) );
  XOR U14448 ( .A(n13623), .B(n13624), .Z(n13626) );
  OR U14449 ( .A(n13600), .B(n13599), .Z(n13604) );
  NANDN U14450 ( .A(n13602), .B(n13601), .Z(n13603) );
  NAND U14451 ( .A(n13604), .B(n13603), .Z(n13625) );
  XNOR U14452 ( .A(n13626), .B(n13625), .Z(n13611) );
  NANDN U14453 ( .A(n13606), .B(n13605), .Z(n13610) );
  OR U14454 ( .A(n13608), .B(n13607), .Z(n13609) );
  NAND U14455 ( .A(n13610), .B(n13609), .Z(n13612) );
  XNOR U14456 ( .A(n13611), .B(n13612), .Z(n13613) );
  XNOR U14457 ( .A(n13614), .B(n13613), .Z(n13629) );
  XNOR U14458 ( .A(n13629), .B(sreg[1564]), .Z(n13630) );
  XOR U14459 ( .A(n13631), .B(n13630), .Z(c[1564]) );
  NANDN U14460 ( .A(n13612), .B(n13611), .Z(n13616) );
  NAND U14461 ( .A(n13614), .B(n13613), .Z(n13615) );
  NAND U14462 ( .A(n13616), .B(n13615), .Z(n13642) );
  AND U14463 ( .A(b[2]), .B(a[543]), .Z(n13648) );
  AND U14464 ( .A(a[544]), .B(b[1]), .Z(n13646) );
  AND U14465 ( .A(a[542]), .B(b[3]), .Z(n13645) );
  XOR U14466 ( .A(n13646), .B(n13645), .Z(n13647) );
  XOR U14467 ( .A(n13648), .B(n13647), .Z(n13651) );
  NAND U14468 ( .A(b[0]), .B(a[545]), .Z(n13652) );
  XOR U14469 ( .A(n13651), .B(n13652), .Z(n13654) );
  OR U14470 ( .A(n13618), .B(n13617), .Z(n13622) );
  NANDN U14471 ( .A(n13620), .B(n13619), .Z(n13621) );
  NAND U14472 ( .A(n13622), .B(n13621), .Z(n13653) );
  XNOR U14473 ( .A(n13654), .B(n13653), .Z(n13639) );
  NANDN U14474 ( .A(n13624), .B(n13623), .Z(n13628) );
  OR U14475 ( .A(n13626), .B(n13625), .Z(n13627) );
  NAND U14476 ( .A(n13628), .B(n13627), .Z(n13640) );
  XNOR U14477 ( .A(n13639), .B(n13640), .Z(n13641) );
  XNOR U14478 ( .A(n13642), .B(n13641), .Z(n13634) );
  XNOR U14479 ( .A(n13634), .B(sreg[1565]), .Z(n13636) );
  NAND U14480 ( .A(n13629), .B(sreg[1564]), .Z(n13633) );
  OR U14481 ( .A(n13631), .B(n13630), .Z(n13632) );
  AND U14482 ( .A(n13633), .B(n13632), .Z(n13635) );
  XOR U14483 ( .A(n13636), .B(n13635), .Z(c[1565]) );
  NAND U14484 ( .A(n13634), .B(sreg[1565]), .Z(n13638) );
  OR U14485 ( .A(n13636), .B(n13635), .Z(n13637) );
  NAND U14486 ( .A(n13638), .B(n13637), .Z(n13659) );
  NANDN U14487 ( .A(n13640), .B(n13639), .Z(n13644) );
  NAND U14488 ( .A(n13642), .B(n13641), .Z(n13643) );
  NAND U14489 ( .A(n13644), .B(n13643), .Z(n13665) );
  AND U14490 ( .A(b[2]), .B(a[544]), .Z(n13671) );
  AND U14491 ( .A(a[545]), .B(b[1]), .Z(n13669) );
  AND U14492 ( .A(a[543]), .B(b[3]), .Z(n13668) );
  XOR U14493 ( .A(n13669), .B(n13668), .Z(n13670) );
  XOR U14494 ( .A(n13671), .B(n13670), .Z(n13674) );
  NAND U14495 ( .A(b[0]), .B(a[546]), .Z(n13675) );
  XOR U14496 ( .A(n13674), .B(n13675), .Z(n13677) );
  OR U14497 ( .A(n13646), .B(n13645), .Z(n13650) );
  NANDN U14498 ( .A(n13648), .B(n13647), .Z(n13649) );
  NAND U14499 ( .A(n13650), .B(n13649), .Z(n13676) );
  XNOR U14500 ( .A(n13677), .B(n13676), .Z(n13662) );
  NANDN U14501 ( .A(n13652), .B(n13651), .Z(n13656) );
  OR U14502 ( .A(n13654), .B(n13653), .Z(n13655) );
  NAND U14503 ( .A(n13656), .B(n13655), .Z(n13663) );
  XNOR U14504 ( .A(n13662), .B(n13663), .Z(n13664) );
  XNOR U14505 ( .A(n13665), .B(n13664), .Z(n13657) );
  XOR U14506 ( .A(sreg[1566]), .B(n13657), .Z(n13658) );
  XOR U14507 ( .A(n13659), .B(n13658), .Z(c[1566]) );
  OR U14508 ( .A(n13657), .B(sreg[1566]), .Z(n13661) );
  NANDN U14509 ( .A(n13659), .B(n13658), .Z(n13660) );
  AND U14510 ( .A(n13661), .B(n13660), .Z(n13681) );
  NANDN U14511 ( .A(n13663), .B(n13662), .Z(n13667) );
  NAND U14512 ( .A(n13665), .B(n13664), .Z(n13666) );
  NAND U14513 ( .A(n13667), .B(n13666), .Z(n13686) );
  AND U14514 ( .A(b[2]), .B(a[545]), .Z(n13692) );
  AND U14515 ( .A(a[546]), .B(b[1]), .Z(n13690) );
  AND U14516 ( .A(a[544]), .B(b[3]), .Z(n13689) );
  XOR U14517 ( .A(n13690), .B(n13689), .Z(n13691) );
  XOR U14518 ( .A(n13692), .B(n13691), .Z(n13695) );
  NAND U14519 ( .A(b[0]), .B(a[547]), .Z(n13696) );
  XOR U14520 ( .A(n13695), .B(n13696), .Z(n13698) );
  OR U14521 ( .A(n13669), .B(n13668), .Z(n13673) );
  NANDN U14522 ( .A(n13671), .B(n13670), .Z(n13672) );
  NAND U14523 ( .A(n13673), .B(n13672), .Z(n13697) );
  XNOR U14524 ( .A(n13698), .B(n13697), .Z(n13683) );
  NANDN U14525 ( .A(n13675), .B(n13674), .Z(n13679) );
  OR U14526 ( .A(n13677), .B(n13676), .Z(n13678) );
  NAND U14527 ( .A(n13679), .B(n13678), .Z(n13684) );
  XNOR U14528 ( .A(n13683), .B(n13684), .Z(n13685) );
  XNOR U14529 ( .A(n13686), .B(n13685), .Z(n13682) );
  XOR U14530 ( .A(sreg[1567]), .B(n13682), .Z(n13680) );
  XOR U14531 ( .A(n13681), .B(n13680), .Z(c[1567]) );
  NANDN U14532 ( .A(n13684), .B(n13683), .Z(n13688) );
  NAND U14533 ( .A(n13686), .B(n13685), .Z(n13687) );
  NAND U14534 ( .A(n13688), .B(n13687), .Z(n13704) );
  AND U14535 ( .A(b[2]), .B(a[546]), .Z(n13716) );
  AND U14536 ( .A(a[547]), .B(b[1]), .Z(n13714) );
  AND U14537 ( .A(a[545]), .B(b[3]), .Z(n13713) );
  XOR U14538 ( .A(n13714), .B(n13713), .Z(n13715) );
  XOR U14539 ( .A(n13716), .B(n13715), .Z(n13707) );
  NAND U14540 ( .A(b[0]), .B(a[548]), .Z(n13708) );
  XOR U14541 ( .A(n13707), .B(n13708), .Z(n13710) );
  OR U14542 ( .A(n13690), .B(n13689), .Z(n13694) );
  NANDN U14543 ( .A(n13692), .B(n13691), .Z(n13693) );
  NAND U14544 ( .A(n13694), .B(n13693), .Z(n13709) );
  XNOR U14545 ( .A(n13710), .B(n13709), .Z(n13701) );
  NANDN U14546 ( .A(n13696), .B(n13695), .Z(n13700) );
  OR U14547 ( .A(n13698), .B(n13697), .Z(n13699) );
  NAND U14548 ( .A(n13700), .B(n13699), .Z(n13702) );
  XNOR U14549 ( .A(n13701), .B(n13702), .Z(n13703) );
  XNOR U14550 ( .A(n13704), .B(n13703), .Z(n13719) );
  XNOR U14551 ( .A(n13719), .B(sreg[1568]), .Z(n13721) );
  XNOR U14552 ( .A(n13720), .B(n13721), .Z(c[1568]) );
  NANDN U14553 ( .A(n13702), .B(n13701), .Z(n13706) );
  NAND U14554 ( .A(n13704), .B(n13703), .Z(n13705) );
  NAND U14555 ( .A(n13706), .B(n13705), .Z(n13744) );
  NANDN U14556 ( .A(n13708), .B(n13707), .Z(n13712) );
  OR U14557 ( .A(n13710), .B(n13709), .Z(n13711) );
  NAND U14558 ( .A(n13712), .B(n13711), .Z(n13741) );
  AND U14559 ( .A(b[2]), .B(a[547]), .Z(n13732) );
  AND U14560 ( .A(a[548]), .B(b[1]), .Z(n13730) );
  AND U14561 ( .A(a[546]), .B(b[3]), .Z(n13729) );
  XOR U14562 ( .A(n13730), .B(n13729), .Z(n13731) );
  XOR U14563 ( .A(n13732), .B(n13731), .Z(n13735) );
  NAND U14564 ( .A(b[0]), .B(a[549]), .Z(n13736) );
  XNOR U14565 ( .A(n13735), .B(n13736), .Z(n13737) );
  OR U14566 ( .A(n13714), .B(n13713), .Z(n13718) );
  NANDN U14567 ( .A(n13716), .B(n13715), .Z(n13717) );
  AND U14568 ( .A(n13718), .B(n13717), .Z(n13738) );
  XNOR U14569 ( .A(n13737), .B(n13738), .Z(n13742) );
  XNOR U14570 ( .A(n13741), .B(n13742), .Z(n13743) );
  XNOR U14571 ( .A(n13744), .B(n13743), .Z(n13724) );
  XOR U14572 ( .A(sreg[1569]), .B(n13724), .Z(n13725) );
  NAND U14573 ( .A(n13719), .B(sreg[1568]), .Z(n13723) );
  NANDN U14574 ( .A(n13721), .B(n13720), .Z(n13722) );
  NAND U14575 ( .A(n13723), .B(n13722), .Z(n13726) );
  XOR U14576 ( .A(n13725), .B(n13726), .Z(c[1569]) );
  OR U14577 ( .A(n13724), .B(sreg[1569]), .Z(n13728) );
  NANDN U14578 ( .A(n13726), .B(n13725), .Z(n13727) );
  NAND U14579 ( .A(n13728), .B(n13727), .Z(n13767) );
  AND U14580 ( .A(b[2]), .B(a[548]), .Z(n13756) );
  AND U14581 ( .A(a[549]), .B(b[1]), .Z(n13754) );
  AND U14582 ( .A(a[547]), .B(b[3]), .Z(n13753) );
  XOR U14583 ( .A(n13754), .B(n13753), .Z(n13755) );
  XOR U14584 ( .A(n13756), .B(n13755), .Z(n13759) );
  NAND U14585 ( .A(b[0]), .B(a[550]), .Z(n13760) );
  XOR U14586 ( .A(n13759), .B(n13760), .Z(n13762) );
  OR U14587 ( .A(n13730), .B(n13729), .Z(n13734) );
  NANDN U14588 ( .A(n13732), .B(n13731), .Z(n13733) );
  NAND U14589 ( .A(n13734), .B(n13733), .Z(n13761) );
  XNOR U14590 ( .A(n13762), .B(n13761), .Z(n13747) );
  NANDN U14591 ( .A(n13736), .B(n13735), .Z(n13740) );
  NAND U14592 ( .A(n13738), .B(n13737), .Z(n13739) );
  NAND U14593 ( .A(n13740), .B(n13739), .Z(n13748) );
  XNOR U14594 ( .A(n13747), .B(n13748), .Z(n13749) );
  NANDN U14595 ( .A(n13742), .B(n13741), .Z(n13746) );
  NANDN U14596 ( .A(n13744), .B(n13743), .Z(n13745) );
  NAND U14597 ( .A(n13746), .B(n13745), .Z(n13750) );
  XOR U14598 ( .A(n13749), .B(n13750), .Z(n13765) );
  XNOR U14599 ( .A(n13765), .B(sreg[1570]), .Z(n13766) );
  XOR U14600 ( .A(n13767), .B(n13766), .Z(c[1570]) );
  NANDN U14601 ( .A(n13748), .B(n13747), .Z(n13752) );
  NANDN U14602 ( .A(n13750), .B(n13749), .Z(n13751) );
  NAND U14603 ( .A(n13752), .B(n13751), .Z(n13790) );
  AND U14604 ( .A(b[2]), .B(a[549]), .Z(n13784) );
  AND U14605 ( .A(a[550]), .B(b[1]), .Z(n13782) );
  AND U14606 ( .A(a[548]), .B(b[3]), .Z(n13781) );
  XOR U14607 ( .A(n13782), .B(n13781), .Z(n13783) );
  XOR U14608 ( .A(n13784), .B(n13783), .Z(n13775) );
  NAND U14609 ( .A(b[0]), .B(a[551]), .Z(n13776) );
  XOR U14610 ( .A(n13775), .B(n13776), .Z(n13778) );
  OR U14611 ( .A(n13754), .B(n13753), .Z(n13758) );
  NANDN U14612 ( .A(n13756), .B(n13755), .Z(n13757) );
  NAND U14613 ( .A(n13758), .B(n13757), .Z(n13777) );
  XNOR U14614 ( .A(n13778), .B(n13777), .Z(n13787) );
  NANDN U14615 ( .A(n13760), .B(n13759), .Z(n13764) );
  OR U14616 ( .A(n13762), .B(n13761), .Z(n13763) );
  NAND U14617 ( .A(n13764), .B(n13763), .Z(n13788) );
  XNOR U14618 ( .A(n13787), .B(n13788), .Z(n13789) );
  XNOR U14619 ( .A(n13790), .B(n13789), .Z(n13770) );
  XNOR U14620 ( .A(n13770), .B(sreg[1571]), .Z(n13772) );
  NAND U14621 ( .A(n13765), .B(sreg[1570]), .Z(n13769) );
  OR U14622 ( .A(n13767), .B(n13766), .Z(n13768) );
  AND U14623 ( .A(n13769), .B(n13768), .Z(n13771) );
  XOR U14624 ( .A(n13772), .B(n13771), .Z(c[1571]) );
  NAND U14625 ( .A(n13770), .B(sreg[1571]), .Z(n13774) );
  OR U14626 ( .A(n13772), .B(n13771), .Z(n13773) );
  NAND U14627 ( .A(n13774), .B(n13773), .Z(n13794) );
  NANDN U14628 ( .A(n13776), .B(n13775), .Z(n13780) );
  OR U14629 ( .A(n13778), .B(n13777), .Z(n13779) );
  NAND U14630 ( .A(n13780), .B(n13779), .Z(n13808) );
  AND U14631 ( .A(b[2]), .B(a[550]), .Z(n13799) );
  AND U14632 ( .A(a[551]), .B(b[1]), .Z(n13797) );
  AND U14633 ( .A(a[549]), .B(b[3]), .Z(n13796) );
  XOR U14634 ( .A(n13797), .B(n13796), .Z(n13798) );
  XOR U14635 ( .A(n13799), .B(n13798), .Z(n13802) );
  NAND U14636 ( .A(b[0]), .B(a[552]), .Z(n13803) );
  XNOR U14637 ( .A(n13802), .B(n13803), .Z(n13804) );
  OR U14638 ( .A(n13782), .B(n13781), .Z(n13786) );
  NANDN U14639 ( .A(n13784), .B(n13783), .Z(n13785) );
  AND U14640 ( .A(n13786), .B(n13785), .Z(n13805) );
  XNOR U14641 ( .A(n13804), .B(n13805), .Z(n13809) );
  XNOR U14642 ( .A(n13808), .B(n13809), .Z(n13810) );
  NANDN U14643 ( .A(n13788), .B(n13787), .Z(n13792) );
  NAND U14644 ( .A(n13790), .B(n13789), .Z(n13791) );
  AND U14645 ( .A(n13792), .B(n13791), .Z(n13811) );
  XNOR U14646 ( .A(n13810), .B(n13811), .Z(n13795) );
  XOR U14647 ( .A(sreg[1572]), .B(n13795), .Z(n13793) );
  XNOR U14648 ( .A(n13794), .B(n13793), .Z(c[1572]) );
  AND U14649 ( .A(b[2]), .B(a[551]), .Z(n13823) );
  AND U14650 ( .A(a[552]), .B(b[1]), .Z(n13821) );
  AND U14651 ( .A(a[550]), .B(b[3]), .Z(n13820) );
  XOR U14652 ( .A(n13821), .B(n13820), .Z(n13822) );
  XOR U14653 ( .A(n13823), .B(n13822), .Z(n13826) );
  NAND U14654 ( .A(b[0]), .B(a[553]), .Z(n13827) );
  XOR U14655 ( .A(n13826), .B(n13827), .Z(n13829) );
  OR U14656 ( .A(n13797), .B(n13796), .Z(n13801) );
  NANDN U14657 ( .A(n13799), .B(n13798), .Z(n13800) );
  NAND U14658 ( .A(n13801), .B(n13800), .Z(n13828) );
  XNOR U14659 ( .A(n13829), .B(n13828), .Z(n13814) );
  NANDN U14660 ( .A(n13803), .B(n13802), .Z(n13807) );
  NAND U14661 ( .A(n13805), .B(n13804), .Z(n13806) );
  NAND U14662 ( .A(n13807), .B(n13806), .Z(n13815) );
  XNOR U14663 ( .A(n13814), .B(n13815), .Z(n13816) );
  NANDN U14664 ( .A(n13809), .B(n13808), .Z(n13813) );
  NAND U14665 ( .A(n13811), .B(n13810), .Z(n13812) );
  NAND U14666 ( .A(n13813), .B(n13812), .Z(n13817) );
  XOR U14667 ( .A(n13816), .B(n13817), .Z(n13832) );
  XNOR U14668 ( .A(n13832), .B(sreg[1573]), .Z(n13833) );
  XOR U14669 ( .A(n13834), .B(n13833), .Z(c[1573]) );
  NANDN U14670 ( .A(n13815), .B(n13814), .Z(n13819) );
  NANDN U14671 ( .A(n13817), .B(n13816), .Z(n13818) );
  NAND U14672 ( .A(n13819), .B(n13818), .Z(n13853) );
  AND U14673 ( .A(b[2]), .B(a[552]), .Z(n13847) );
  AND U14674 ( .A(a[553]), .B(b[1]), .Z(n13845) );
  AND U14675 ( .A(a[551]), .B(b[3]), .Z(n13844) );
  XOR U14676 ( .A(n13845), .B(n13844), .Z(n13846) );
  XOR U14677 ( .A(n13847), .B(n13846), .Z(n13838) );
  NAND U14678 ( .A(b[0]), .B(a[554]), .Z(n13839) );
  XOR U14679 ( .A(n13838), .B(n13839), .Z(n13841) );
  OR U14680 ( .A(n13821), .B(n13820), .Z(n13825) );
  NANDN U14681 ( .A(n13823), .B(n13822), .Z(n13824) );
  NAND U14682 ( .A(n13825), .B(n13824), .Z(n13840) );
  XNOR U14683 ( .A(n13841), .B(n13840), .Z(n13850) );
  NANDN U14684 ( .A(n13827), .B(n13826), .Z(n13831) );
  OR U14685 ( .A(n13829), .B(n13828), .Z(n13830) );
  NAND U14686 ( .A(n13831), .B(n13830), .Z(n13851) );
  XNOR U14687 ( .A(n13850), .B(n13851), .Z(n13852) );
  XOR U14688 ( .A(n13853), .B(n13852), .Z(n13857) );
  NAND U14689 ( .A(n13832), .B(sreg[1573]), .Z(n13836) );
  OR U14690 ( .A(n13834), .B(n13833), .Z(n13835) );
  NAND U14691 ( .A(n13836), .B(n13835), .Z(n13856) );
  XNOR U14692 ( .A(sreg[1574]), .B(n13856), .Z(n13837) );
  XOR U14693 ( .A(n13857), .B(n13837), .Z(c[1574]) );
  NANDN U14694 ( .A(n13839), .B(n13838), .Z(n13843) );
  OR U14695 ( .A(n13841), .B(n13840), .Z(n13842) );
  NAND U14696 ( .A(n13843), .B(n13842), .Z(n13861) );
  AND U14697 ( .A(b[2]), .B(a[553]), .Z(n13870) );
  AND U14698 ( .A(a[554]), .B(b[1]), .Z(n13868) );
  AND U14699 ( .A(a[552]), .B(b[3]), .Z(n13867) );
  XOR U14700 ( .A(n13868), .B(n13867), .Z(n13869) );
  XOR U14701 ( .A(n13870), .B(n13869), .Z(n13873) );
  NAND U14702 ( .A(b[0]), .B(a[555]), .Z(n13874) );
  XNOR U14703 ( .A(n13873), .B(n13874), .Z(n13875) );
  OR U14704 ( .A(n13845), .B(n13844), .Z(n13849) );
  NANDN U14705 ( .A(n13847), .B(n13846), .Z(n13848) );
  AND U14706 ( .A(n13849), .B(n13848), .Z(n13876) );
  XNOR U14707 ( .A(n13875), .B(n13876), .Z(n13862) );
  XNOR U14708 ( .A(n13861), .B(n13862), .Z(n13863) );
  NANDN U14709 ( .A(n13851), .B(n13850), .Z(n13855) );
  NAND U14710 ( .A(n13853), .B(n13852), .Z(n13854) );
  AND U14711 ( .A(n13855), .B(n13854), .Z(n13864) );
  XNOR U14712 ( .A(n13863), .B(n13864), .Z(n13860) );
  XNOR U14713 ( .A(sreg[1575]), .B(n13859), .Z(n13858) );
  XOR U14714 ( .A(n13860), .B(n13858), .Z(c[1575]) );
  NANDN U14715 ( .A(n13862), .B(n13861), .Z(n13866) );
  NAND U14716 ( .A(n13864), .B(n13863), .Z(n13865) );
  NAND U14717 ( .A(n13866), .B(n13865), .Z(n13882) );
  AND U14718 ( .A(b[2]), .B(a[554]), .Z(n13888) );
  AND U14719 ( .A(a[555]), .B(b[1]), .Z(n13886) );
  AND U14720 ( .A(a[553]), .B(b[3]), .Z(n13885) );
  XOR U14721 ( .A(n13886), .B(n13885), .Z(n13887) );
  XOR U14722 ( .A(n13888), .B(n13887), .Z(n13891) );
  NAND U14723 ( .A(b[0]), .B(a[556]), .Z(n13892) );
  XOR U14724 ( .A(n13891), .B(n13892), .Z(n13894) );
  OR U14725 ( .A(n13868), .B(n13867), .Z(n13872) );
  NANDN U14726 ( .A(n13870), .B(n13869), .Z(n13871) );
  NAND U14727 ( .A(n13872), .B(n13871), .Z(n13893) );
  XNOR U14728 ( .A(n13894), .B(n13893), .Z(n13879) );
  NANDN U14729 ( .A(n13874), .B(n13873), .Z(n13878) );
  NAND U14730 ( .A(n13876), .B(n13875), .Z(n13877) );
  NAND U14731 ( .A(n13878), .B(n13877), .Z(n13880) );
  XNOR U14732 ( .A(n13879), .B(n13880), .Z(n13881) );
  XOR U14733 ( .A(n13882), .B(n13881), .Z(n13897) );
  XNOR U14734 ( .A(n13897), .B(sreg[1576]), .Z(n13898) );
  XOR U14735 ( .A(n13899), .B(n13898), .Z(c[1576]) );
  NANDN U14736 ( .A(n13880), .B(n13879), .Z(n13884) );
  NANDN U14737 ( .A(n13882), .B(n13881), .Z(n13883) );
  NAND U14738 ( .A(n13884), .B(n13883), .Z(n13917) );
  AND U14739 ( .A(b[2]), .B(a[555]), .Z(n13911) );
  AND U14740 ( .A(a[556]), .B(b[1]), .Z(n13909) );
  AND U14741 ( .A(a[554]), .B(b[3]), .Z(n13908) );
  XOR U14742 ( .A(n13909), .B(n13908), .Z(n13910) );
  XOR U14743 ( .A(n13911), .B(n13910), .Z(n13902) );
  NAND U14744 ( .A(b[0]), .B(a[557]), .Z(n13903) );
  XOR U14745 ( .A(n13902), .B(n13903), .Z(n13905) );
  OR U14746 ( .A(n13886), .B(n13885), .Z(n13890) );
  NANDN U14747 ( .A(n13888), .B(n13887), .Z(n13889) );
  NAND U14748 ( .A(n13890), .B(n13889), .Z(n13904) );
  XNOR U14749 ( .A(n13905), .B(n13904), .Z(n13914) );
  NANDN U14750 ( .A(n13892), .B(n13891), .Z(n13896) );
  OR U14751 ( .A(n13894), .B(n13893), .Z(n13895) );
  NAND U14752 ( .A(n13896), .B(n13895), .Z(n13915) );
  XNOR U14753 ( .A(n13914), .B(n13915), .Z(n13916) );
  XNOR U14754 ( .A(n13917), .B(n13916), .Z(n13920) );
  XNOR U14755 ( .A(n13920), .B(sreg[1577]), .Z(n13922) );
  NAND U14756 ( .A(n13897), .B(sreg[1576]), .Z(n13901) );
  OR U14757 ( .A(n13899), .B(n13898), .Z(n13900) );
  AND U14758 ( .A(n13901), .B(n13900), .Z(n13921) );
  XOR U14759 ( .A(n13922), .B(n13921), .Z(c[1577]) );
  NANDN U14760 ( .A(n13903), .B(n13902), .Z(n13907) );
  OR U14761 ( .A(n13905), .B(n13904), .Z(n13906) );
  NAND U14762 ( .A(n13907), .B(n13906), .Z(n13925) );
  AND U14763 ( .A(b[2]), .B(a[556]), .Z(n13934) );
  AND U14764 ( .A(a[557]), .B(b[1]), .Z(n13932) );
  AND U14765 ( .A(a[555]), .B(b[3]), .Z(n13931) );
  XOR U14766 ( .A(n13932), .B(n13931), .Z(n13933) );
  XOR U14767 ( .A(n13934), .B(n13933), .Z(n13937) );
  NAND U14768 ( .A(b[0]), .B(a[558]), .Z(n13938) );
  XNOR U14769 ( .A(n13937), .B(n13938), .Z(n13939) );
  OR U14770 ( .A(n13909), .B(n13908), .Z(n13913) );
  NANDN U14771 ( .A(n13911), .B(n13910), .Z(n13912) );
  AND U14772 ( .A(n13913), .B(n13912), .Z(n13940) );
  XNOR U14773 ( .A(n13939), .B(n13940), .Z(n13926) );
  XNOR U14774 ( .A(n13925), .B(n13926), .Z(n13927) );
  NANDN U14775 ( .A(n13915), .B(n13914), .Z(n13919) );
  NAND U14776 ( .A(n13917), .B(n13916), .Z(n13918) );
  AND U14777 ( .A(n13919), .B(n13918), .Z(n13928) );
  XOR U14778 ( .A(n13927), .B(n13928), .Z(n13943) );
  XNOR U14779 ( .A(sreg[1578]), .B(n13943), .Z(n13945) );
  NAND U14780 ( .A(n13920), .B(sreg[1577]), .Z(n13924) );
  OR U14781 ( .A(n13922), .B(n13921), .Z(n13923) );
  AND U14782 ( .A(n13924), .B(n13923), .Z(n13944) );
  XOR U14783 ( .A(n13945), .B(n13944), .Z(c[1578]) );
  NANDN U14784 ( .A(n13926), .B(n13925), .Z(n13930) );
  NAND U14785 ( .A(n13928), .B(n13927), .Z(n13929) );
  NAND U14786 ( .A(n13930), .B(n13929), .Z(n13951) );
  AND U14787 ( .A(b[2]), .B(a[557]), .Z(n13957) );
  AND U14788 ( .A(a[558]), .B(b[1]), .Z(n13955) );
  AND U14789 ( .A(a[556]), .B(b[3]), .Z(n13954) );
  XOR U14790 ( .A(n13955), .B(n13954), .Z(n13956) );
  XOR U14791 ( .A(n13957), .B(n13956), .Z(n13960) );
  NAND U14792 ( .A(b[0]), .B(a[559]), .Z(n13961) );
  XOR U14793 ( .A(n13960), .B(n13961), .Z(n13963) );
  OR U14794 ( .A(n13932), .B(n13931), .Z(n13936) );
  NANDN U14795 ( .A(n13934), .B(n13933), .Z(n13935) );
  NAND U14796 ( .A(n13936), .B(n13935), .Z(n13962) );
  XNOR U14797 ( .A(n13963), .B(n13962), .Z(n13948) );
  NANDN U14798 ( .A(n13938), .B(n13937), .Z(n13942) );
  NAND U14799 ( .A(n13940), .B(n13939), .Z(n13941) );
  NAND U14800 ( .A(n13942), .B(n13941), .Z(n13949) );
  XNOR U14801 ( .A(n13948), .B(n13949), .Z(n13950) );
  XOR U14802 ( .A(n13951), .B(n13950), .Z(n13966) );
  XNOR U14803 ( .A(n13966), .B(sreg[1579]), .Z(n13968) );
  NAND U14804 ( .A(sreg[1578]), .B(n13943), .Z(n13947) );
  OR U14805 ( .A(n13945), .B(n13944), .Z(n13946) );
  AND U14806 ( .A(n13947), .B(n13946), .Z(n13967) );
  XOR U14807 ( .A(n13968), .B(n13967), .Z(c[1579]) );
  NANDN U14808 ( .A(n13949), .B(n13948), .Z(n13953) );
  NANDN U14809 ( .A(n13951), .B(n13950), .Z(n13952) );
  NAND U14810 ( .A(n13953), .B(n13952), .Z(n13991) );
  AND U14811 ( .A(b[2]), .B(a[558]), .Z(n13985) );
  AND U14812 ( .A(a[559]), .B(b[1]), .Z(n13983) );
  AND U14813 ( .A(a[557]), .B(b[3]), .Z(n13982) );
  XOR U14814 ( .A(n13983), .B(n13982), .Z(n13984) );
  XOR U14815 ( .A(n13985), .B(n13984), .Z(n13976) );
  NAND U14816 ( .A(b[0]), .B(a[560]), .Z(n13977) );
  XOR U14817 ( .A(n13976), .B(n13977), .Z(n13979) );
  OR U14818 ( .A(n13955), .B(n13954), .Z(n13959) );
  NANDN U14819 ( .A(n13957), .B(n13956), .Z(n13958) );
  NAND U14820 ( .A(n13959), .B(n13958), .Z(n13978) );
  XNOR U14821 ( .A(n13979), .B(n13978), .Z(n13988) );
  NANDN U14822 ( .A(n13961), .B(n13960), .Z(n13965) );
  OR U14823 ( .A(n13963), .B(n13962), .Z(n13964) );
  NAND U14824 ( .A(n13965), .B(n13964), .Z(n13989) );
  XNOR U14825 ( .A(n13988), .B(n13989), .Z(n13990) );
  XNOR U14826 ( .A(n13991), .B(n13990), .Z(n13971) );
  XNOR U14827 ( .A(n13971), .B(sreg[1580]), .Z(n13973) );
  NAND U14828 ( .A(n13966), .B(sreg[1579]), .Z(n13970) );
  OR U14829 ( .A(n13968), .B(n13967), .Z(n13969) );
  AND U14830 ( .A(n13970), .B(n13969), .Z(n13972) );
  XOR U14831 ( .A(n13973), .B(n13972), .Z(c[1580]) );
  NAND U14832 ( .A(n13971), .B(sreg[1580]), .Z(n13975) );
  OR U14833 ( .A(n13973), .B(n13972), .Z(n13974) );
  NAND U14834 ( .A(n13975), .B(n13974), .Z(n14013) );
  NANDN U14835 ( .A(n13977), .B(n13976), .Z(n13981) );
  OR U14836 ( .A(n13979), .B(n13978), .Z(n13980) );
  NAND U14837 ( .A(n13981), .B(n13980), .Z(n13995) );
  AND U14838 ( .A(b[2]), .B(a[559]), .Z(n14004) );
  AND U14839 ( .A(a[560]), .B(b[1]), .Z(n14002) );
  AND U14840 ( .A(a[558]), .B(b[3]), .Z(n14001) );
  XOR U14841 ( .A(n14002), .B(n14001), .Z(n14003) );
  XOR U14842 ( .A(n14004), .B(n14003), .Z(n14007) );
  NAND U14843 ( .A(b[0]), .B(a[561]), .Z(n14008) );
  XNOR U14844 ( .A(n14007), .B(n14008), .Z(n14009) );
  OR U14845 ( .A(n13983), .B(n13982), .Z(n13987) );
  NANDN U14846 ( .A(n13985), .B(n13984), .Z(n13986) );
  AND U14847 ( .A(n13987), .B(n13986), .Z(n14010) );
  XNOR U14848 ( .A(n14009), .B(n14010), .Z(n13996) );
  XNOR U14849 ( .A(n13995), .B(n13996), .Z(n13997) );
  NANDN U14850 ( .A(n13989), .B(n13988), .Z(n13993) );
  NAND U14851 ( .A(n13991), .B(n13990), .Z(n13992) );
  AND U14852 ( .A(n13993), .B(n13992), .Z(n13998) );
  XNOR U14853 ( .A(n13997), .B(n13998), .Z(n14014) );
  XOR U14854 ( .A(sreg[1581]), .B(n14014), .Z(n13994) );
  XNOR U14855 ( .A(n14013), .B(n13994), .Z(c[1581]) );
  NANDN U14856 ( .A(n13996), .B(n13995), .Z(n14000) );
  NAND U14857 ( .A(n13998), .B(n13997), .Z(n13999) );
  NAND U14858 ( .A(n14000), .B(n13999), .Z(n14021) );
  AND U14859 ( .A(b[2]), .B(a[560]), .Z(n14027) );
  AND U14860 ( .A(a[561]), .B(b[1]), .Z(n14025) );
  AND U14861 ( .A(a[559]), .B(b[3]), .Z(n14024) );
  XOR U14862 ( .A(n14025), .B(n14024), .Z(n14026) );
  XOR U14863 ( .A(n14027), .B(n14026), .Z(n14030) );
  NAND U14864 ( .A(b[0]), .B(a[562]), .Z(n14031) );
  XOR U14865 ( .A(n14030), .B(n14031), .Z(n14033) );
  OR U14866 ( .A(n14002), .B(n14001), .Z(n14006) );
  NANDN U14867 ( .A(n14004), .B(n14003), .Z(n14005) );
  NAND U14868 ( .A(n14006), .B(n14005), .Z(n14032) );
  XNOR U14869 ( .A(n14033), .B(n14032), .Z(n14018) );
  NANDN U14870 ( .A(n14008), .B(n14007), .Z(n14012) );
  NAND U14871 ( .A(n14010), .B(n14009), .Z(n14011) );
  NAND U14872 ( .A(n14012), .B(n14011), .Z(n14019) );
  XNOR U14873 ( .A(n14018), .B(n14019), .Z(n14020) );
  XOR U14874 ( .A(n14021), .B(n14020), .Z(n14017) );
  XNOR U14875 ( .A(sreg[1582]), .B(n14016), .Z(n14015) );
  XNOR U14876 ( .A(n14017), .B(n14015), .Z(c[1582]) );
  NANDN U14877 ( .A(n14019), .B(n14018), .Z(n14023) );
  NANDN U14878 ( .A(n14021), .B(n14020), .Z(n14022) );
  NAND U14879 ( .A(n14023), .B(n14022), .Z(n14039) );
  AND U14880 ( .A(b[2]), .B(a[561]), .Z(n14045) );
  AND U14881 ( .A(a[562]), .B(b[1]), .Z(n14043) );
  AND U14882 ( .A(a[560]), .B(b[3]), .Z(n14042) );
  XOR U14883 ( .A(n14043), .B(n14042), .Z(n14044) );
  XOR U14884 ( .A(n14045), .B(n14044), .Z(n14048) );
  NAND U14885 ( .A(b[0]), .B(a[563]), .Z(n14049) );
  XOR U14886 ( .A(n14048), .B(n14049), .Z(n14051) );
  OR U14887 ( .A(n14025), .B(n14024), .Z(n14029) );
  NANDN U14888 ( .A(n14027), .B(n14026), .Z(n14028) );
  NAND U14889 ( .A(n14029), .B(n14028), .Z(n14050) );
  XNOR U14890 ( .A(n14051), .B(n14050), .Z(n14036) );
  NANDN U14891 ( .A(n14031), .B(n14030), .Z(n14035) );
  OR U14892 ( .A(n14033), .B(n14032), .Z(n14034) );
  NAND U14893 ( .A(n14035), .B(n14034), .Z(n14037) );
  XNOR U14894 ( .A(n14036), .B(n14037), .Z(n14038) );
  XNOR U14895 ( .A(n14039), .B(n14038), .Z(n14055) );
  XNOR U14896 ( .A(n14055), .B(sreg[1583]), .Z(n14056) );
  XOR U14897 ( .A(n14057), .B(n14056), .Z(c[1583]) );
  NANDN U14898 ( .A(n14037), .B(n14036), .Z(n14041) );
  NAND U14899 ( .A(n14039), .B(n14038), .Z(n14040) );
  NAND U14900 ( .A(n14041), .B(n14040), .Z(n14062) );
  AND U14901 ( .A(b[2]), .B(a[562]), .Z(n14070) );
  AND U14902 ( .A(a[563]), .B(b[1]), .Z(n14068) );
  AND U14903 ( .A(a[561]), .B(b[3]), .Z(n14067) );
  XOR U14904 ( .A(n14068), .B(n14067), .Z(n14069) );
  XOR U14905 ( .A(n14070), .B(n14069), .Z(n14063) );
  NAND U14906 ( .A(b[0]), .B(a[564]), .Z(n14064) );
  XOR U14907 ( .A(n14063), .B(n14064), .Z(n14065) );
  OR U14908 ( .A(n14043), .B(n14042), .Z(n14047) );
  NANDN U14909 ( .A(n14045), .B(n14044), .Z(n14046) );
  AND U14910 ( .A(n14047), .B(n14046), .Z(n14066) );
  XOR U14911 ( .A(n14065), .B(n14066), .Z(n14060) );
  NANDN U14912 ( .A(n14049), .B(n14048), .Z(n14053) );
  OR U14913 ( .A(n14051), .B(n14050), .Z(n14052) );
  AND U14914 ( .A(n14053), .B(n14052), .Z(n14061) );
  XOR U14915 ( .A(n14060), .B(n14061), .Z(n14054) );
  XOR U14916 ( .A(n14062), .B(n14054), .Z(n14073) );
  XOR U14917 ( .A(sreg[1584]), .B(n14073), .Z(n14075) );
  NAND U14918 ( .A(n14055), .B(sreg[1583]), .Z(n14059) );
  OR U14919 ( .A(n14057), .B(n14056), .Z(n14058) );
  NAND U14920 ( .A(n14059), .B(n14058), .Z(n14074) );
  XNOR U14921 ( .A(n14075), .B(n14074), .Z(c[1584]) );
  AND U14922 ( .A(b[2]), .B(a[563]), .Z(n14082) );
  AND U14923 ( .A(a[564]), .B(b[1]), .Z(n14080) );
  AND U14924 ( .A(a[562]), .B(b[3]), .Z(n14079) );
  XOR U14925 ( .A(n14080), .B(n14079), .Z(n14081) );
  XOR U14926 ( .A(n14082), .B(n14081), .Z(n14085) );
  NAND U14927 ( .A(b[0]), .B(a[565]), .Z(n14086) );
  XNOR U14928 ( .A(n14085), .B(n14086), .Z(n14087) );
  OR U14929 ( .A(n14068), .B(n14067), .Z(n14072) );
  NANDN U14930 ( .A(n14070), .B(n14069), .Z(n14071) );
  AND U14931 ( .A(n14072), .B(n14071), .Z(n14088) );
  XNOR U14932 ( .A(n14087), .B(n14088), .Z(n14092) );
  XNOR U14933 ( .A(n14091), .B(n14092), .Z(n14093) );
  XOR U14934 ( .A(n14094), .B(n14093), .Z(n14097) );
  NANDN U14935 ( .A(sreg[1584]), .B(n14073), .Z(n14077) );
  OR U14936 ( .A(n14075), .B(n14074), .Z(n14076) );
  NAND U14937 ( .A(n14077), .B(n14076), .Z(n14098) );
  XNOR U14938 ( .A(n14098), .B(sreg[1585]), .Z(n14078) );
  XNOR U14939 ( .A(n14097), .B(n14078), .Z(c[1585]) );
  AND U14940 ( .A(b[2]), .B(a[564]), .Z(n14111) );
  AND U14941 ( .A(a[565]), .B(b[1]), .Z(n14109) );
  AND U14942 ( .A(a[563]), .B(b[3]), .Z(n14108) );
  XOR U14943 ( .A(n14109), .B(n14108), .Z(n14110) );
  XOR U14944 ( .A(n14111), .B(n14110), .Z(n14114) );
  NAND U14945 ( .A(b[0]), .B(a[566]), .Z(n14115) );
  XOR U14946 ( .A(n14114), .B(n14115), .Z(n14117) );
  OR U14947 ( .A(n14080), .B(n14079), .Z(n14084) );
  NANDN U14948 ( .A(n14082), .B(n14081), .Z(n14083) );
  NAND U14949 ( .A(n14084), .B(n14083), .Z(n14116) );
  XNOR U14950 ( .A(n14117), .B(n14116), .Z(n14102) );
  NANDN U14951 ( .A(n14086), .B(n14085), .Z(n14090) );
  NAND U14952 ( .A(n14088), .B(n14087), .Z(n14089) );
  NAND U14953 ( .A(n14090), .B(n14089), .Z(n14103) );
  XNOR U14954 ( .A(n14102), .B(n14103), .Z(n14104) );
  NANDN U14955 ( .A(n14092), .B(n14091), .Z(n14096) );
  NANDN U14956 ( .A(n14094), .B(n14093), .Z(n14095) );
  NAND U14957 ( .A(n14096), .B(n14095), .Z(n14105) );
  XOR U14958 ( .A(n14104), .B(n14105), .Z(n14101) );
  XOR U14959 ( .A(sreg[1586]), .B(n14100), .Z(n14099) );
  XNOR U14960 ( .A(n14101), .B(n14099), .Z(c[1586]) );
  NANDN U14961 ( .A(n14103), .B(n14102), .Z(n14107) );
  NANDN U14962 ( .A(n14105), .B(n14104), .Z(n14106) );
  NAND U14963 ( .A(n14107), .B(n14106), .Z(n14140) );
  AND U14964 ( .A(b[2]), .B(a[565]), .Z(n14134) );
  AND U14965 ( .A(a[566]), .B(b[1]), .Z(n14132) );
  AND U14966 ( .A(a[564]), .B(b[3]), .Z(n14131) );
  XOR U14967 ( .A(n14132), .B(n14131), .Z(n14133) );
  XOR U14968 ( .A(n14134), .B(n14133), .Z(n14125) );
  NAND U14969 ( .A(b[0]), .B(a[567]), .Z(n14126) );
  XOR U14970 ( .A(n14125), .B(n14126), .Z(n14128) );
  OR U14971 ( .A(n14109), .B(n14108), .Z(n14113) );
  NANDN U14972 ( .A(n14111), .B(n14110), .Z(n14112) );
  NAND U14973 ( .A(n14113), .B(n14112), .Z(n14127) );
  XNOR U14974 ( .A(n14128), .B(n14127), .Z(n14137) );
  NANDN U14975 ( .A(n14115), .B(n14114), .Z(n14119) );
  OR U14976 ( .A(n14117), .B(n14116), .Z(n14118) );
  NAND U14977 ( .A(n14119), .B(n14118), .Z(n14138) );
  XNOR U14978 ( .A(n14137), .B(n14138), .Z(n14139) );
  XNOR U14979 ( .A(n14140), .B(n14139), .Z(n14120) );
  XNOR U14980 ( .A(n14120), .B(sreg[1587]), .Z(n14121) );
  XOR U14981 ( .A(n14122), .B(n14121), .Z(c[1587]) );
  NAND U14982 ( .A(n14120), .B(sreg[1587]), .Z(n14124) );
  OR U14983 ( .A(n14122), .B(n14121), .Z(n14123) );
  AND U14984 ( .A(n14124), .B(n14123), .Z(n14163) );
  NANDN U14985 ( .A(n14126), .B(n14125), .Z(n14130) );
  OR U14986 ( .A(n14128), .B(n14127), .Z(n14129) );
  NAND U14987 ( .A(n14130), .B(n14129), .Z(n14156) );
  AND U14988 ( .A(b[2]), .B(a[566]), .Z(n14147) );
  AND U14989 ( .A(a[567]), .B(b[1]), .Z(n14145) );
  AND U14990 ( .A(a[565]), .B(b[3]), .Z(n14144) );
  XOR U14991 ( .A(n14145), .B(n14144), .Z(n14146) );
  XOR U14992 ( .A(n14147), .B(n14146), .Z(n14150) );
  NAND U14993 ( .A(b[0]), .B(a[568]), .Z(n14151) );
  XNOR U14994 ( .A(n14150), .B(n14151), .Z(n14152) );
  OR U14995 ( .A(n14132), .B(n14131), .Z(n14136) );
  NANDN U14996 ( .A(n14134), .B(n14133), .Z(n14135) );
  AND U14997 ( .A(n14136), .B(n14135), .Z(n14153) );
  XNOR U14998 ( .A(n14152), .B(n14153), .Z(n14157) );
  XNOR U14999 ( .A(n14156), .B(n14157), .Z(n14158) );
  NANDN U15000 ( .A(n14138), .B(n14137), .Z(n14142) );
  NAND U15001 ( .A(n14140), .B(n14139), .Z(n14141) );
  AND U15002 ( .A(n14142), .B(n14141), .Z(n14159) );
  XOR U15003 ( .A(n14158), .B(n14159), .Z(n14162) );
  XNOR U15004 ( .A(sreg[1588]), .B(n14162), .Z(n14143) );
  XOR U15005 ( .A(n14163), .B(n14143), .Z(c[1588]) );
  AND U15006 ( .A(b[2]), .B(a[567]), .Z(n14176) );
  AND U15007 ( .A(a[568]), .B(b[1]), .Z(n14174) );
  AND U15008 ( .A(a[566]), .B(b[3]), .Z(n14173) );
  XOR U15009 ( .A(n14174), .B(n14173), .Z(n14175) );
  XOR U15010 ( .A(n14176), .B(n14175), .Z(n14179) );
  NAND U15011 ( .A(b[0]), .B(a[569]), .Z(n14180) );
  XOR U15012 ( .A(n14179), .B(n14180), .Z(n14182) );
  OR U15013 ( .A(n14145), .B(n14144), .Z(n14149) );
  NANDN U15014 ( .A(n14147), .B(n14146), .Z(n14148) );
  NAND U15015 ( .A(n14149), .B(n14148), .Z(n14181) );
  XNOR U15016 ( .A(n14182), .B(n14181), .Z(n14167) );
  NANDN U15017 ( .A(n14151), .B(n14150), .Z(n14155) );
  NAND U15018 ( .A(n14153), .B(n14152), .Z(n14154) );
  NAND U15019 ( .A(n14155), .B(n14154), .Z(n14168) );
  XNOR U15020 ( .A(n14167), .B(n14168), .Z(n14169) );
  NANDN U15021 ( .A(n14157), .B(n14156), .Z(n14161) );
  NAND U15022 ( .A(n14159), .B(n14158), .Z(n14160) );
  NAND U15023 ( .A(n14161), .B(n14160), .Z(n14170) );
  XOR U15024 ( .A(n14169), .B(n14170), .Z(n14166) );
  XNOR U15025 ( .A(sreg[1589]), .B(n14165), .Z(n14164) );
  XNOR U15026 ( .A(n14166), .B(n14164), .Z(c[1589]) );
  NANDN U15027 ( .A(n14168), .B(n14167), .Z(n14172) );
  NANDN U15028 ( .A(n14170), .B(n14169), .Z(n14171) );
  NAND U15029 ( .A(n14172), .B(n14171), .Z(n14188) );
  AND U15030 ( .A(b[2]), .B(a[568]), .Z(n14194) );
  AND U15031 ( .A(a[569]), .B(b[1]), .Z(n14192) );
  AND U15032 ( .A(a[567]), .B(b[3]), .Z(n14191) );
  XOR U15033 ( .A(n14192), .B(n14191), .Z(n14193) );
  XOR U15034 ( .A(n14194), .B(n14193), .Z(n14197) );
  NAND U15035 ( .A(b[0]), .B(a[570]), .Z(n14198) );
  XOR U15036 ( .A(n14197), .B(n14198), .Z(n14200) );
  OR U15037 ( .A(n14174), .B(n14173), .Z(n14178) );
  NANDN U15038 ( .A(n14176), .B(n14175), .Z(n14177) );
  NAND U15039 ( .A(n14178), .B(n14177), .Z(n14199) );
  XNOR U15040 ( .A(n14200), .B(n14199), .Z(n14185) );
  NANDN U15041 ( .A(n14180), .B(n14179), .Z(n14184) );
  OR U15042 ( .A(n14182), .B(n14181), .Z(n14183) );
  NAND U15043 ( .A(n14184), .B(n14183), .Z(n14186) );
  XNOR U15044 ( .A(n14185), .B(n14186), .Z(n14187) );
  XNOR U15045 ( .A(n14188), .B(n14187), .Z(n14203) );
  XNOR U15046 ( .A(n14203), .B(sreg[1590]), .Z(n14204) );
  XOR U15047 ( .A(n14205), .B(n14204), .Z(c[1590]) );
  NANDN U15048 ( .A(n14186), .B(n14185), .Z(n14190) );
  NAND U15049 ( .A(n14188), .B(n14187), .Z(n14189) );
  NAND U15050 ( .A(n14190), .B(n14189), .Z(n14214) );
  AND U15051 ( .A(b[2]), .B(a[569]), .Z(n14220) );
  AND U15052 ( .A(a[570]), .B(b[1]), .Z(n14218) );
  AND U15053 ( .A(a[568]), .B(b[3]), .Z(n14217) );
  XOR U15054 ( .A(n14218), .B(n14217), .Z(n14219) );
  XOR U15055 ( .A(n14220), .B(n14219), .Z(n14223) );
  NAND U15056 ( .A(b[0]), .B(a[571]), .Z(n14224) );
  XOR U15057 ( .A(n14223), .B(n14224), .Z(n14226) );
  OR U15058 ( .A(n14192), .B(n14191), .Z(n14196) );
  NANDN U15059 ( .A(n14194), .B(n14193), .Z(n14195) );
  NAND U15060 ( .A(n14196), .B(n14195), .Z(n14225) );
  XNOR U15061 ( .A(n14226), .B(n14225), .Z(n14211) );
  NANDN U15062 ( .A(n14198), .B(n14197), .Z(n14202) );
  OR U15063 ( .A(n14200), .B(n14199), .Z(n14201) );
  NAND U15064 ( .A(n14202), .B(n14201), .Z(n14212) );
  XNOR U15065 ( .A(n14211), .B(n14212), .Z(n14213) );
  XNOR U15066 ( .A(n14214), .B(n14213), .Z(n14210) );
  NAND U15067 ( .A(n14203), .B(sreg[1590]), .Z(n14207) );
  OR U15068 ( .A(n14205), .B(n14204), .Z(n14206) );
  AND U15069 ( .A(n14207), .B(n14206), .Z(n14209) );
  XNOR U15070 ( .A(n14209), .B(sreg[1591]), .Z(n14208) );
  XOR U15071 ( .A(n14210), .B(n14208), .Z(c[1591]) );
  NANDN U15072 ( .A(n14212), .B(n14211), .Z(n14216) );
  NAND U15073 ( .A(n14214), .B(n14213), .Z(n14215) );
  NAND U15074 ( .A(n14216), .B(n14215), .Z(n14232) );
  AND U15075 ( .A(b[2]), .B(a[570]), .Z(n14238) );
  AND U15076 ( .A(a[571]), .B(b[1]), .Z(n14236) );
  AND U15077 ( .A(a[569]), .B(b[3]), .Z(n14235) );
  XOR U15078 ( .A(n14236), .B(n14235), .Z(n14237) );
  XOR U15079 ( .A(n14238), .B(n14237), .Z(n14241) );
  NAND U15080 ( .A(b[0]), .B(a[572]), .Z(n14242) );
  XOR U15081 ( .A(n14241), .B(n14242), .Z(n14244) );
  OR U15082 ( .A(n14218), .B(n14217), .Z(n14222) );
  NANDN U15083 ( .A(n14220), .B(n14219), .Z(n14221) );
  NAND U15084 ( .A(n14222), .B(n14221), .Z(n14243) );
  XNOR U15085 ( .A(n14244), .B(n14243), .Z(n14229) );
  NANDN U15086 ( .A(n14224), .B(n14223), .Z(n14228) );
  OR U15087 ( .A(n14226), .B(n14225), .Z(n14227) );
  NAND U15088 ( .A(n14228), .B(n14227), .Z(n14230) );
  XNOR U15089 ( .A(n14229), .B(n14230), .Z(n14231) );
  XNOR U15090 ( .A(n14232), .B(n14231), .Z(n14247) );
  XNOR U15091 ( .A(n14247), .B(sreg[1592]), .Z(n14249) );
  XNOR U15092 ( .A(n14248), .B(n14249), .Z(c[1592]) );
  NANDN U15093 ( .A(n14230), .B(n14229), .Z(n14234) );
  NAND U15094 ( .A(n14232), .B(n14231), .Z(n14233) );
  NAND U15095 ( .A(n14234), .B(n14233), .Z(n14258) );
  AND U15096 ( .A(b[2]), .B(a[571]), .Z(n14264) );
  AND U15097 ( .A(a[572]), .B(b[1]), .Z(n14262) );
  AND U15098 ( .A(a[570]), .B(b[3]), .Z(n14261) );
  XOR U15099 ( .A(n14262), .B(n14261), .Z(n14263) );
  XOR U15100 ( .A(n14264), .B(n14263), .Z(n14267) );
  NAND U15101 ( .A(b[0]), .B(a[573]), .Z(n14268) );
  XOR U15102 ( .A(n14267), .B(n14268), .Z(n14270) );
  OR U15103 ( .A(n14236), .B(n14235), .Z(n14240) );
  NANDN U15104 ( .A(n14238), .B(n14237), .Z(n14239) );
  NAND U15105 ( .A(n14240), .B(n14239), .Z(n14269) );
  XNOR U15106 ( .A(n14270), .B(n14269), .Z(n14255) );
  NANDN U15107 ( .A(n14242), .B(n14241), .Z(n14246) );
  OR U15108 ( .A(n14244), .B(n14243), .Z(n14245) );
  NAND U15109 ( .A(n14246), .B(n14245), .Z(n14256) );
  XNOR U15110 ( .A(n14255), .B(n14256), .Z(n14257) );
  XOR U15111 ( .A(n14258), .B(n14257), .Z(n14254) );
  NAND U15112 ( .A(n14247), .B(sreg[1592]), .Z(n14251) );
  NANDN U15113 ( .A(n14249), .B(n14248), .Z(n14250) );
  NAND U15114 ( .A(n14251), .B(n14250), .Z(n14253) );
  XNOR U15115 ( .A(sreg[1593]), .B(n14253), .Z(n14252) );
  XOR U15116 ( .A(n14254), .B(n14252), .Z(c[1593]) );
  NANDN U15117 ( .A(n14256), .B(n14255), .Z(n14260) );
  NAND U15118 ( .A(n14258), .B(n14257), .Z(n14259) );
  NAND U15119 ( .A(n14260), .B(n14259), .Z(n14276) );
  AND U15120 ( .A(b[2]), .B(a[572]), .Z(n14282) );
  AND U15121 ( .A(a[573]), .B(b[1]), .Z(n14280) );
  AND U15122 ( .A(a[571]), .B(b[3]), .Z(n14279) );
  XOR U15123 ( .A(n14280), .B(n14279), .Z(n14281) );
  XOR U15124 ( .A(n14282), .B(n14281), .Z(n14285) );
  NAND U15125 ( .A(b[0]), .B(a[574]), .Z(n14286) );
  XOR U15126 ( .A(n14285), .B(n14286), .Z(n14288) );
  OR U15127 ( .A(n14262), .B(n14261), .Z(n14266) );
  NANDN U15128 ( .A(n14264), .B(n14263), .Z(n14265) );
  NAND U15129 ( .A(n14266), .B(n14265), .Z(n14287) );
  XNOR U15130 ( .A(n14288), .B(n14287), .Z(n14273) );
  NANDN U15131 ( .A(n14268), .B(n14267), .Z(n14272) );
  OR U15132 ( .A(n14270), .B(n14269), .Z(n14271) );
  NAND U15133 ( .A(n14272), .B(n14271), .Z(n14274) );
  XNOR U15134 ( .A(n14273), .B(n14274), .Z(n14275) );
  XNOR U15135 ( .A(n14276), .B(n14275), .Z(n14291) );
  XNOR U15136 ( .A(n14291), .B(sreg[1594]), .Z(n14292) );
  XOR U15137 ( .A(n14293), .B(n14292), .Z(c[1594]) );
  NANDN U15138 ( .A(n14274), .B(n14273), .Z(n14278) );
  NAND U15139 ( .A(n14276), .B(n14275), .Z(n14277) );
  NAND U15140 ( .A(n14278), .B(n14277), .Z(n14302) );
  AND U15141 ( .A(b[2]), .B(a[573]), .Z(n14308) );
  AND U15142 ( .A(a[574]), .B(b[1]), .Z(n14306) );
  AND U15143 ( .A(a[572]), .B(b[3]), .Z(n14305) );
  XOR U15144 ( .A(n14306), .B(n14305), .Z(n14307) );
  XOR U15145 ( .A(n14308), .B(n14307), .Z(n14311) );
  NAND U15146 ( .A(b[0]), .B(a[575]), .Z(n14312) );
  XOR U15147 ( .A(n14311), .B(n14312), .Z(n14314) );
  OR U15148 ( .A(n14280), .B(n14279), .Z(n14284) );
  NANDN U15149 ( .A(n14282), .B(n14281), .Z(n14283) );
  NAND U15150 ( .A(n14284), .B(n14283), .Z(n14313) );
  XNOR U15151 ( .A(n14314), .B(n14313), .Z(n14299) );
  NANDN U15152 ( .A(n14286), .B(n14285), .Z(n14290) );
  OR U15153 ( .A(n14288), .B(n14287), .Z(n14289) );
  NAND U15154 ( .A(n14290), .B(n14289), .Z(n14300) );
  XNOR U15155 ( .A(n14299), .B(n14300), .Z(n14301) );
  XNOR U15156 ( .A(n14302), .B(n14301), .Z(n14298) );
  NAND U15157 ( .A(n14291), .B(sreg[1594]), .Z(n14295) );
  OR U15158 ( .A(n14293), .B(n14292), .Z(n14294) );
  AND U15159 ( .A(n14295), .B(n14294), .Z(n14297) );
  XNOR U15160 ( .A(n14297), .B(sreg[1595]), .Z(n14296) );
  XOR U15161 ( .A(n14298), .B(n14296), .Z(c[1595]) );
  NANDN U15162 ( .A(n14300), .B(n14299), .Z(n14304) );
  NAND U15163 ( .A(n14302), .B(n14301), .Z(n14303) );
  NAND U15164 ( .A(n14304), .B(n14303), .Z(n14320) );
  AND U15165 ( .A(b[2]), .B(a[574]), .Z(n14326) );
  AND U15166 ( .A(a[575]), .B(b[1]), .Z(n14324) );
  AND U15167 ( .A(a[573]), .B(b[3]), .Z(n14323) );
  XOR U15168 ( .A(n14324), .B(n14323), .Z(n14325) );
  XOR U15169 ( .A(n14326), .B(n14325), .Z(n14329) );
  NAND U15170 ( .A(b[0]), .B(a[576]), .Z(n14330) );
  XOR U15171 ( .A(n14329), .B(n14330), .Z(n14332) );
  OR U15172 ( .A(n14306), .B(n14305), .Z(n14310) );
  NANDN U15173 ( .A(n14308), .B(n14307), .Z(n14309) );
  NAND U15174 ( .A(n14310), .B(n14309), .Z(n14331) );
  XNOR U15175 ( .A(n14332), .B(n14331), .Z(n14317) );
  NANDN U15176 ( .A(n14312), .B(n14311), .Z(n14316) );
  OR U15177 ( .A(n14314), .B(n14313), .Z(n14315) );
  NAND U15178 ( .A(n14316), .B(n14315), .Z(n14318) );
  XNOR U15179 ( .A(n14317), .B(n14318), .Z(n14319) );
  XOR U15180 ( .A(n14320), .B(n14319), .Z(n14335) );
  XOR U15181 ( .A(sreg[1596]), .B(n14335), .Z(n14337) );
  XNOR U15182 ( .A(n14336), .B(n14337), .Z(c[1596]) );
  NANDN U15183 ( .A(n14318), .B(n14317), .Z(n14322) );
  NAND U15184 ( .A(n14320), .B(n14319), .Z(n14321) );
  NAND U15185 ( .A(n14322), .B(n14321), .Z(n14343) );
  AND U15186 ( .A(b[2]), .B(a[575]), .Z(n14349) );
  AND U15187 ( .A(a[576]), .B(b[1]), .Z(n14347) );
  AND U15188 ( .A(a[574]), .B(b[3]), .Z(n14346) );
  XOR U15189 ( .A(n14347), .B(n14346), .Z(n14348) );
  XOR U15190 ( .A(n14349), .B(n14348), .Z(n14352) );
  NAND U15191 ( .A(b[0]), .B(a[577]), .Z(n14353) );
  XOR U15192 ( .A(n14352), .B(n14353), .Z(n14355) );
  OR U15193 ( .A(n14324), .B(n14323), .Z(n14328) );
  NANDN U15194 ( .A(n14326), .B(n14325), .Z(n14327) );
  NAND U15195 ( .A(n14328), .B(n14327), .Z(n14354) );
  XNOR U15196 ( .A(n14355), .B(n14354), .Z(n14340) );
  NANDN U15197 ( .A(n14330), .B(n14329), .Z(n14334) );
  OR U15198 ( .A(n14332), .B(n14331), .Z(n14333) );
  NAND U15199 ( .A(n14334), .B(n14333), .Z(n14341) );
  XNOR U15200 ( .A(n14340), .B(n14341), .Z(n14342) );
  XNOR U15201 ( .A(n14343), .B(n14342), .Z(n14358) );
  XNOR U15202 ( .A(n14358), .B(sreg[1597]), .Z(n14360) );
  NANDN U15203 ( .A(n14335), .B(sreg[1596]), .Z(n14339) );
  NANDN U15204 ( .A(n14337), .B(n14336), .Z(n14338) );
  AND U15205 ( .A(n14339), .B(n14338), .Z(n14359) );
  XOR U15206 ( .A(n14360), .B(n14359), .Z(c[1597]) );
  NANDN U15207 ( .A(n14341), .B(n14340), .Z(n14345) );
  NAND U15208 ( .A(n14343), .B(n14342), .Z(n14344) );
  NAND U15209 ( .A(n14345), .B(n14344), .Z(n14369) );
  AND U15210 ( .A(b[2]), .B(a[576]), .Z(n14375) );
  AND U15211 ( .A(a[577]), .B(b[1]), .Z(n14373) );
  AND U15212 ( .A(a[575]), .B(b[3]), .Z(n14372) );
  XOR U15213 ( .A(n14373), .B(n14372), .Z(n14374) );
  XOR U15214 ( .A(n14375), .B(n14374), .Z(n14378) );
  NAND U15215 ( .A(b[0]), .B(a[578]), .Z(n14379) );
  XOR U15216 ( .A(n14378), .B(n14379), .Z(n14381) );
  OR U15217 ( .A(n14347), .B(n14346), .Z(n14351) );
  NANDN U15218 ( .A(n14349), .B(n14348), .Z(n14350) );
  NAND U15219 ( .A(n14351), .B(n14350), .Z(n14380) );
  XNOR U15220 ( .A(n14381), .B(n14380), .Z(n14366) );
  NANDN U15221 ( .A(n14353), .B(n14352), .Z(n14357) );
  OR U15222 ( .A(n14355), .B(n14354), .Z(n14356) );
  NAND U15223 ( .A(n14357), .B(n14356), .Z(n14367) );
  XNOR U15224 ( .A(n14366), .B(n14367), .Z(n14368) );
  XNOR U15225 ( .A(n14369), .B(n14368), .Z(n14365) );
  NAND U15226 ( .A(n14358), .B(sreg[1597]), .Z(n14362) );
  OR U15227 ( .A(n14360), .B(n14359), .Z(n14361) );
  AND U15228 ( .A(n14362), .B(n14361), .Z(n14364) );
  XNOR U15229 ( .A(n14364), .B(sreg[1598]), .Z(n14363) );
  XOR U15230 ( .A(n14365), .B(n14363), .Z(c[1598]) );
  NANDN U15231 ( .A(n14367), .B(n14366), .Z(n14371) );
  NAND U15232 ( .A(n14369), .B(n14368), .Z(n14370) );
  NAND U15233 ( .A(n14371), .B(n14370), .Z(n14387) );
  AND U15234 ( .A(b[2]), .B(a[577]), .Z(n14393) );
  AND U15235 ( .A(a[578]), .B(b[1]), .Z(n14391) );
  AND U15236 ( .A(a[576]), .B(b[3]), .Z(n14390) );
  XOR U15237 ( .A(n14391), .B(n14390), .Z(n14392) );
  XOR U15238 ( .A(n14393), .B(n14392), .Z(n14396) );
  NAND U15239 ( .A(b[0]), .B(a[579]), .Z(n14397) );
  XOR U15240 ( .A(n14396), .B(n14397), .Z(n14399) );
  OR U15241 ( .A(n14373), .B(n14372), .Z(n14377) );
  NANDN U15242 ( .A(n14375), .B(n14374), .Z(n14376) );
  NAND U15243 ( .A(n14377), .B(n14376), .Z(n14398) );
  XNOR U15244 ( .A(n14399), .B(n14398), .Z(n14384) );
  NANDN U15245 ( .A(n14379), .B(n14378), .Z(n14383) );
  OR U15246 ( .A(n14381), .B(n14380), .Z(n14382) );
  NAND U15247 ( .A(n14383), .B(n14382), .Z(n14385) );
  XNOR U15248 ( .A(n14384), .B(n14385), .Z(n14386) );
  XNOR U15249 ( .A(n14387), .B(n14386), .Z(n14402) );
  XNOR U15250 ( .A(n14402), .B(sreg[1599]), .Z(n14404) );
  XNOR U15251 ( .A(n14403), .B(n14404), .Z(c[1599]) );
  NANDN U15252 ( .A(n14385), .B(n14384), .Z(n14389) );
  NAND U15253 ( .A(n14387), .B(n14386), .Z(n14388) );
  NAND U15254 ( .A(n14389), .B(n14388), .Z(n14411) );
  AND U15255 ( .A(b[2]), .B(a[578]), .Z(n14417) );
  AND U15256 ( .A(a[579]), .B(b[1]), .Z(n14415) );
  AND U15257 ( .A(a[577]), .B(b[3]), .Z(n14414) );
  XOR U15258 ( .A(n14415), .B(n14414), .Z(n14416) );
  XOR U15259 ( .A(n14417), .B(n14416), .Z(n14420) );
  NAND U15260 ( .A(b[0]), .B(a[580]), .Z(n14421) );
  XOR U15261 ( .A(n14420), .B(n14421), .Z(n14423) );
  OR U15262 ( .A(n14391), .B(n14390), .Z(n14395) );
  NANDN U15263 ( .A(n14393), .B(n14392), .Z(n14394) );
  NAND U15264 ( .A(n14395), .B(n14394), .Z(n14422) );
  XNOR U15265 ( .A(n14423), .B(n14422), .Z(n14408) );
  NANDN U15266 ( .A(n14397), .B(n14396), .Z(n14401) );
  OR U15267 ( .A(n14399), .B(n14398), .Z(n14400) );
  NAND U15268 ( .A(n14401), .B(n14400), .Z(n14409) );
  XNOR U15269 ( .A(n14408), .B(n14409), .Z(n14410) );
  XOR U15270 ( .A(n14411), .B(n14410), .Z(n14427) );
  NAND U15271 ( .A(n14402), .B(sreg[1599]), .Z(n14406) );
  NANDN U15272 ( .A(n14404), .B(n14403), .Z(n14405) );
  NAND U15273 ( .A(n14406), .B(n14405), .Z(n14426) );
  XNOR U15274 ( .A(sreg[1600]), .B(n14426), .Z(n14407) );
  XOR U15275 ( .A(n14427), .B(n14407), .Z(c[1600]) );
  NANDN U15276 ( .A(n14409), .B(n14408), .Z(n14413) );
  NAND U15277 ( .A(n14411), .B(n14410), .Z(n14412) );
  NAND U15278 ( .A(n14413), .B(n14412), .Z(n14432) );
  AND U15279 ( .A(b[2]), .B(a[579]), .Z(n14438) );
  AND U15280 ( .A(a[580]), .B(b[1]), .Z(n14436) );
  AND U15281 ( .A(a[578]), .B(b[3]), .Z(n14435) );
  XOR U15282 ( .A(n14436), .B(n14435), .Z(n14437) );
  XOR U15283 ( .A(n14438), .B(n14437), .Z(n14441) );
  NAND U15284 ( .A(b[0]), .B(a[581]), .Z(n14442) );
  XOR U15285 ( .A(n14441), .B(n14442), .Z(n14444) );
  OR U15286 ( .A(n14415), .B(n14414), .Z(n14419) );
  NANDN U15287 ( .A(n14417), .B(n14416), .Z(n14418) );
  NAND U15288 ( .A(n14419), .B(n14418), .Z(n14443) );
  XNOR U15289 ( .A(n14444), .B(n14443), .Z(n14429) );
  NANDN U15290 ( .A(n14421), .B(n14420), .Z(n14425) );
  OR U15291 ( .A(n14423), .B(n14422), .Z(n14424) );
  NAND U15292 ( .A(n14425), .B(n14424), .Z(n14430) );
  XNOR U15293 ( .A(n14429), .B(n14430), .Z(n14431) );
  XNOR U15294 ( .A(n14432), .B(n14431), .Z(n14448) );
  XOR U15295 ( .A(n14447), .B(sreg[1601]), .Z(n14428) );
  XOR U15296 ( .A(n14448), .B(n14428), .Z(c[1601]) );
  NANDN U15297 ( .A(n14430), .B(n14429), .Z(n14434) );
  NAND U15298 ( .A(n14432), .B(n14431), .Z(n14433) );
  NAND U15299 ( .A(n14434), .B(n14433), .Z(n14455) );
  AND U15300 ( .A(b[2]), .B(a[580]), .Z(n14461) );
  AND U15301 ( .A(a[581]), .B(b[1]), .Z(n14459) );
  AND U15302 ( .A(a[579]), .B(b[3]), .Z(n14458) );
  XOR U15303 ( .A(n14459), .B(n14458), .Z(n14460) );
  XOR U15304 ( .A(n14461), .B(n14460), .Z(n14464) );
  NAND U15305 ( .A(b[0]), .B(a[582]), .Z(n14465) );
  XOR U15306 ( .A(n14464), .B(n14465), .Z(n14467) );
  OR U15307 ( .A(n14436), .B(n14435), .Z(n14440) );
  NANDN U15308 ( .A(n14438), .B(n14437), .Z(n14439) );
  NAND U15309 ( .A(n14440), .B(n14439), .Z(n14466) );
  XNOR U15310 ( .A(n14467), .B(n14466), .Z(n14452) );
  NANDN U15311 ( .A(n14442), .B(n14441), .Z(n14446) );
  OR U15312 ( .A(n14444), .B(n14443), .Z(n14445) );
  NAND U15313 ( .A(n14446), .B(n14445), .Z(n14453) );
  XNOR U15314 ( .A(n14452), .B(n14453), .Z(n14454) );
  XNOR U15315 ( .A(n14455), .B(n14454), .Z(n14451) );
  XOR U15316 ( .A(n14450), .B(sreg[1602]), .Z(n14449) );
  XOR U15317 ( .A(n14451), .B(n14449), .Z(c[1602]) );
  NANDN U15318 ( .A(n14453), .B(n14452), .Z(n14457) );
  NAND U15319 ( .A(n14455), .B(n14454), .Z(n14456) );
  NAND U15320 ( .A(n14457), .B(n14456), .Z(n14473) );
  AND U15321 ( .A(b[2]), .B(a[581]), .Z(n14479) );
  AND U15322 ( .A(a[582]), .B(b[1]), .Z(n14477) );
  AND U15323 ( .A(a[580]), .B(b[3]), .Z(n14476) );
  XOR U15324 ( .A(n14477), .B(n14476), .Z(n14478) );
  XOR U15325 ( .A(n14479), .B(n14478), .Z(n14482) );
  NAND U15326 ( .A(b[0]), .B(a[583]), .Z(n14483) );
  XOR U15327 ( .A(n14482), .B(n14483), .Z(n14485) );
  OR U15328 ( .A(n14459), .B(n14458), .Z(n14463) );
  NANDN U15329 ( .A(n14461), .B(n14460), .Z(n14462) );
  NAND U15330 ( .A(n14463), .B(n14462), .Z(n14484) );
  XNOR U15331 ( .A(n14485), .B(n14484), .Z(n14470) );
  NANDN U15332 ( .A(n14465), .B(n14464), .Z(n14469) );
  OR U15333 ( .A(n14467), .B(n14466), .Z(n14468) );
  NAND U15334 ( .A(n14469), .B(n14468), .Z(n14471) );
  XNOR U15335 ( .A(n14470), .B(n14471), .Z(n14472) );
  XNOR U15336 ( .A(n14473), .B(n14472), .Z(n14488) );
  XNOR U15337 ( .A(n14488), .B(sreg[1603]), .Z(n14490) );
  XNOR U15338 ( .A(n14489), .B(n14490), .Z(c[1603]) );
  NANDN U15339 ( .A(n14471), .B(n14470), .Z(n14475) );
  NAND U15340 ( .A(n14473), .B(n14472), .Z(n14474) );
  NAND U15341 ( .A(n14475), .B(n14474), .Z(n14499) );
  AND U15342 ( .A(b[2]), .B(a[582]), .Z(n14505) );
  AND U15343 ( .A(a[583]), .B(b[1]), .Z(n14503) );
  AND U15344 ( .A(a[581]), .B(b[3]), .Z(n14502) );
  XOR U15345 ( .A(n14503), .B(n14502), .Z(n14504) );
  XOR U15346 ( .A(n14505), .B(n14504), .Z(n14508) );
  NAND U15347 ( .A(b[0]), .B(a[584]), .Z(n14509) );
  XOR U15348 ( .A(n14508), .B(n14509), .Z(n14511) );
  OR U15349 ( .A(n14477), .B(n14476), .Z(n14481) );
  NANDN U15350 ( .A(n14479), .B(n14478), .Z(n14480) );
  NAND U15351 ( .A(n14481), .B(n14480), .Z(n14510) );
  XNOR U15352 ( .A(n14511), .B(n14510), .Z(n14496) );
  NANDN U15353 ( .A(n14483), .B(n14482), .Z(n14487) );
  OR U15354 ( .A(n14485), .B(n14484), .Z(n14486) );
  NAND U15355 ( .A(n14487), .B(n14486), .Z(n14497) );
  XNOR U15356 ( .A(n14496), .B(n14497), .Z(n14498) );
  XOR U15357 ( .A(n14499), .B(n14498), .Z(n14495) );
  NAND U15358 ( .A(n14488), .B(sreg[1603]), .Z(n14492) );
  NANDN U15359 ( .A(n14490), .B(n14489), .Z(n14491) );
  NAND U15360 ( .A(n14492), .B(n14491), .Z(n14494) );
  XNOR U15361 ( .A(sreg[1604]), .B(n14494), .Z(n14493) );
  XOR U15362 ( .A(n14495), .B(n14493), .Z(c[1604]) );
  NANDN U15363 ( .A(n14497), .B(n14496), .Z(n14501) );
  NAND U15364 ( .A(n14499), .B(n14498), .Z(n14500) );
  NAND U15365 ( .A(n14501), .B(n14500), .Z(n14517) );
  AND U15366 ( .A(b[2]), .B(a[583]), .Z(n14523) );
  AND U15367 ( .A(a[584]), .B(b[1]), .Z(n14521) );
  AND U15368 ( .A(a[582]), .B(b[3]), .Z(n14520) );
  XOR U15369 ( .A(n14521), .B(n14520), .Z(n14522) );
  XOR U15370 ( .A(n14523), .B(n14522), .Z(n14526) );
  NAND U15371 ( .A(b[0]), .B(a[585]), .Z(n14527) );
  XOR U15372 ( .A(n14526), .B(n14527), .Z(n14529) );
  OR U15373 ( .A(n14503), .B(n14502), .Z(n14507) );
  NANDN U15374 ( .A(n14505), .B(n14504), .Z(n14506) );
  NAND U15375 ( .A(n14507), .B(n14506), .Z(n14528) );
  XNOR U15376 ( .A(n14529), .B(n14528), .Z(n14514) );
  NANDN U15377 ( .A(n14509), .B(n14508), .Z(n14513) );
  OR U15378 ( .A(n14511), .B(n14510), .Z(n14512) );
  NAND U15379 ( .A(n14513), .B(n14512), .Z(n14515) );
  XNOR U15380 ( .A(n14514), .B(n14515), .Z(n14516) );
  XNOR U15381 ( .A(n14517), .B(n14516), .Z(n14532) );
  XNOR U15382 ( .A(n14532), .B(sreg[1605]), .Z(n14533) );
  XOR U15383 ( .A(n14534), .B(n14533), .Z(c[1605]) );
  NANDN U15384 ( .A(n14515), .B(n14514), .Z(n14519) );
  NAND U15385 ( .A(n14517), .B(n14516), .Z(n14518) );
  NAND U15386 ( .A(n14519), .B(n14518), .Z(n14540) );
  AND U15387 ( .A(b[2]), .B(a[584]), .Z(n14552) );
  AND U15388 ( .A(a[585]), .B(b[1]), .Z(n14550) );
  AND U15389 ( .A(a[583]), .B(b[3]), .Z(n14549) );
  XOR U15390 ( .A(n14550), .B(n14549), .Z(n14551) );
  XOR U15391 ( .A(n14552), .B(n14551), .Z(n14543) );
  NAND U15392 ( .A(b[0]), .B(a[586]), .Z(n14544) );
  XOR U15393 ( .A(n14543), .B(n14544), .Z(n14546) );
  OR U15394 ( .A(n14521), .B(n14520), .Z(n14525) );
  NANDN U15395 ( .A(n14523), .B(n14522), .Z(n14524) );
  NAND U15396 ( .A(n14525), .B(n14524), .Z(n14545) );
  XNOR U15397 ( .A(n14546), .B(n14545), .Z(n14537) );
  NANDN U15398 ( .A(n14527), .B(n14526), .Z(n14531) );
  OR U15399 ( .A(n14529), .B(n14528), .Z(n14530) );
  NAND U15400 ( .A(n14531), .B(n14530), .Z(n14538) );
  XNOR U15401 ( .A(n14537), .B(n14538), .Z(n14539) );
  XNOR U15402 ( .A(n14540), .B(n14539), .Z(n14555) );
  XOR U15403 ( .A(sreg[1606]), .B(n14555), .Z(n14556) );
  NAND U15404 ( .A(n14532), .B(sreg[1605]), .Z(n14536) );
  OR U15405 ( .A(n14534), .B(n14533), .Z(n14535) );
  NAND U15406 ( .A(n14536), .B(n14535), .Z(n14557) );
  XOR U15407 ( .A(n14556), .B(n14557), .Z(c[1606]) );
  NANDN U15408 ( .A(n14538), .B(n14537), .Z(n14542) );
  NAND U15409 ( .A(n14540), .B(n14539), .Z(n14541) );
  NAND U15410 ( .A(n14542), .B(n14541), .Z(n14564) );
  NANDN U15411 ( .A(n14544), .B(n14543), .Z(n14548) );
  OR U15412 ( .A(n14546), .B(n14545), .Z(n14547) );
  NAND U15413 ( .A(n14548), .B(n14547), .Z(n14561) );
  AND U15414 ( .A(b[2]), .B(a[585]), .Z(n14570) );
  AND U15415 ( .A(a[586]), .B(b[1]), .Z(n14568) );
  AND U15416 ( .A(a[584]), .B(b[3]), .Z(n14567) );
  XOR U15417 ( .A(n14568), .B(n14567), .Z(n14569) );
  XOR U15418 ( .A(n14570), .B(n14569), .Z(n14573) );
  NAND U15419 ( .A(b[0]), .B(a[587]), .Z(n14574) );
  XNOR U15420 ( .A(n14573), .B(n14574), .Z(n14575) );
  OR U15421 ( .A(n14550), .B(n14549), .Z(n14554) );
  NANDN U15422 ( .A(n14552), .B(n14551), .Z(n14553) );
  AND U15423 ( .A(n14554), .B(n14553), .Z(n14576) );
  XNOR U15424 ( .A(n14575), .B(n14576), .Z(n14562) );
  XNOR U15425 ( .A(n14561), .B(n14562), .Z(n14563) );
  XNOR U15426 ( .A(n14564), .B(n14563), .Z(n14580) );
  OR U15427 ( .A(n14555), .B(sreg[1606]), .Z(n14559) );
  NANDN U15428 ( .A(n14557), .B(n14556), .Z(n14558) );
  AND U15429 ( .A(n14559), .B(n14558), .Z(n14579) );
  XNOR U15430 ( .A(sreg[1607]), .B(n14579), .Z(n14560) );
  XNOR U15431 ( .A(n14580), .B(n14560), .Z(c[1607]) );
  NANDN U15432 ( .A(n14562), .B(n14561), .Z(n14566) );
  NANDN U15433 ( .A(n14564), .B(n14563), .Z(n14565) );
  NAND U15434 ( .A(n14566), .B(n14565), .Z(n14587) );
  AND U15435 ( .A(b[2]), .B(a[586]), .Z(n14593) );
  AND U15436 ( .A(a[587]), .B(b[1]), .Z(n14591) );
  AND U15437 ( .A(a[585]), .B(b[3]), .Z(n14590) );
  XOR U15438 ( .A(n14591), .B(n14590), .Z(n14592) );
  XOR U15439 ( .A(n14593), .B(n14592), .Z(n14596) );
  NAND U15440 ( .A(b[0]), .B(a[588]), .Z(n14597) );
  XOR U15441 ( .A(n14596), .B(n14597), .Z(n14599) );
  OR U15442 ( .A(n14568), .B(n14567), .Z(n14572) );
  NANDN U15443 ( .A(n14570), .B(n14569), .Z(n14571) );
  NAND U15444 ( .A(n14572), .B(n14571), .Z(n14598) );
  XNOR U15445 ( .A(n14599), .B(n14598), .Z(n14584) );
  NANDN U15446 ( .A(n14574), .B(n14573), .Z(n14578) );
  NAND U15447 ( .A(n14576), .B(n14575), .Z(n14577) );
  NAND U15448 ( .A(n14578), .B(n14577), .Z(n14585) );
  XNOR U15449 ( .A(n14584), .B(n14585), .Z(n14586) );
  XNOR U15450 ( .A(n14587), .B(n14586), .Z(n14583) );
  XOR U15451 ( .A(n14582), .B(sreg[1608]), .Z(n14581) );
  XNOR U15452 ( .A(n14583), .B(n14581), .Z(c[1608]) );
  NANDN U15453 ( .A(n14585), .B(n14584), .Z(n14589) );
  NANDN U15454 ( .A(n14587), .B(n14586), .Z(n14588) );
  NAND U15455 ( .A(n14589), .B(n14588), .Z(n14622) );
  AND U15456 ( .A(b[2]), .B(a[587]), .Z(n14616) );
  AND U15457 ( .A(a[588]), .B(b[1]), .Z(n14614) );
  AND U15458 ( .A(a[586]), .B(b[3]), .Z(n14613) );
  XOR U15459 ( .A(n14614), .B(n14613), .Z(n14615) );
  XOR U15460 ( .A(n14616), .B(n14615), .Z(n14607) );
  NAND U15461 ( .A(b[0]), .B(a[589]), .Z(n14608) );
  XOR U15462 ( .A(n14607), .B(n14608), .Z(n14610) );
  OR U15463 ( .A(n14591), .B(n14590), .Z(n14595) );
  NANDN U15464 ( .A(n14593), .B(n14592), .Z(n14594) );
  NAND U15465 ( .A(n14595), .B(n14594), .Z(n14609) );
  XNOR U15466 ( .A(n14610), .B(n14609), .Z(n14619) );
  NANDN U15467 ( .A(n14597), .B(n14596), .Z(n14601) );
  OR U15468 ( .A(n14599), .B(n14598), .Z(n14600) );
  NAND U15469 ( .A(n14601), .B(n14600), .Z(n14620) );
  XNOR U15470 ( .A(n14619), .B(n14620), .Z(n14621) );
  XNOR U15471 ( .A(n14622), .B(n14621), .Z(n14602) );
  XNOR U15472 ( .A(n14602), .B(sreg[1609]), .Z(n14604) );
  XNOR U15473 ( .A(n14603), .B(n14604), .Z(c[1609]) );
  NAND U15474 ( .A(n14602), .B(sreg[1609]), .Z(n14606) );
  NANDN U15475 ( .A(n14604), .B(n14603), .Z(n14605) );
  NAND U15476 ( .A(n14606), .B(n14605), .Z(n14626) );
  NANDN U15477 ( .A(n14608), .B(n14607), .Z(n14612) );
  OR U15478 ( .A(n14610), .B(n14609), .Z(n14611) );
  NAND U15479 ( .A(n14612), .B(n14611), .Z(n14628) );
  AND U15480 ( .A(b[2]), .B(a[588]), .Z(n14637) );
  AND U15481 ( .A(a[589]), .B(b[1]), .Z(n14635) );
  AND U15482 ( .A(a[587]), .B(b[3]), .Z(n14634) );
  XOR U15483 ( .A(n14635), .B(n14634), .Z(n14636) );
  XOR U15484 ( .A(n14637), .B(n14636), .Z(n14640) );
  NAND U15485 ( .A(b[0]), .B(a[590]), .Z(n14641) );
  XNOR U15486 ( .A(n14640), .B(n14641), .Z(n14642) );
  OR U15487 ( .A(n14614), .B(n14613), .Z(n14618) );
  NANDN U15488 ( .A(n14616), .B(n14615), .Z(n14617) );
  AND U15489 ( .A(n14618), .B(n14617), .Z(n14643) );
  XNOR U15490 ( .A(n14642), .B(n14643), .Z(n14629) );
  XNOR U15491 ( .A(n14628), .B(n14629), .Z(n14630) );
  NANDN U15492 ( .A(n14620), .B(n14619), .Z(n14624) );
  NAND U15493 ( .A(n14622), .B(n14621), .Z(n14623) );
  AND U15494 ( .A(n14624), .B(n14623), .Z(n14631) );
  XNOR U15495 ( .A(n14630), .B(n14631), .Z(n14627) );
  XOR U15496 ( .A(sreg[1610]), .B(n14627), .Z(n14625) );
  XNOR U15497 ( .A(n14626), .B(n14625), .Z(c[1610]) );
  NANDN U15498 ( .A(n14629), .B(n14628), .Z(n14633) );
  NAND U15499 ( .A(n14631), .B(n14630), .Z(n14632) );
  NAND U15500 ( .A(n14633), .B(n14632), .Z(n14649) );
  AND U15501 ( .A(b[2]), .B(a[589]), .Z(n14655) );
  AND U15502 ( .A(a[590]), .B(b[1]), .Z(n14653) );
  AND U15503 ( .A(a[588]), .B(b[3]), .Z(n14652) );
  XOR U15504 ( .A(n14653), .B(n14652), .Z(n14654) );
  XOR U15505 ( .A(n14655), .B(n14654), .Z(n14658) );
  NAND U15506 ( .A(b[0]), .B(a[591]), .Z(n14659) );
  XOR U15507 ( .A(n14658), .B(n14659), .Z(n14661) );
  OR U15508 ( .A(n14635), .B(n14634), .Z(n14639) );
  NANDN U15509 ( .A(n14637), .B(n14636), .Z(n14638) );
  NAND U15510 ( .A(n14639), .B(n14638), .Z(n14660) );
  XNOR U15511 ( .A(n14661), .B(n14660), .Z(n14646) );
  NANDN U15512 ( .A(n14641), .B(n14640), .Z(n14645) );
  NAND U15513 ( .A(n14643), .B(n14642), .Z(n14644) );
  NAND U15514 ( .A(n14645), .B(n14644), .Z(n14647) );
  XNOR U15515 ( .A(n14646), .B(n14647), .Z(n14648) );
  XOR U15516 ( .A(n14649), .B(n14648), .Z(n14664) );
  XNOR U15517 ( .A(n14664), .B(sreg[1611]), .Z(n14665) );
  XOR U15518 ( .A(n14666), .B(n14665), .Z(c[1611]) );
  NANDN U15519 ( .A(n14647), .B(n14646), .Z(n14651) );
  NANDN U15520 ( .A(n14649), .B(n14648), .Z(n14650) );
  NAND U15521 ( .A(n14651), .B(n14650), .Z(n14689) );
  AND U15522 ( .A(b[2]), .B(a[590]), .Z(n14683) );
  AND U15523 ( .A(a[591]), .B(b[1]), .Z(n14681) );
  AND U15524 ( .A(a[589]), .B(b[3]), .Z(n14680) );
  XOR U15525 ( .A(n14681), .B(n14680), .Z(n14682) );
  XOR U15526 ( .A(n14683), .B(n14682), .Z(n14674) );
  NAND U15527 ( .A(b[0]), .B(a[592]), .Z(n14675) );
  XOR U15528 ( .A(n14674), .B(n14675), .Z(n14677) );
  OR U15529 ( .A(n14653), .B(n14652), .Z(n14657) );
  NANDN U15530 ( .A(n14655), .B(n14654), .Z(n14656) );
  NAND U15531 ( .A(n14657), .B(n14656), .Z(n14676) );
  XNOR U15532 ( .A(n14677), .B(n14676), .Z(n14686) );
  NANDN U15533 ( .A(n14659), .B(n14658), .Z(n14663) );
  OR U15534 ( .A(n14661), .B(n14660), .Z(n14662) );
  NAND U15535 ( .A(n14663), .B(n14662), .Z(n14687) );
  XNOR U15536 ( .A(n14686), .B(n14687), .Z(n14688) );
  XNOR U15537 ( .A(n14689), .B(n14688), .Z(n14669) );
  XNOR U15538 ( .A(n14669), .B(sreg[1612]), .Z(n14671) );
  NAND U15539 ( .A(n14664), .B(sreg[1611]), .Z(n14668) );
  OR U15540 ( .A(n14666), .B(n14665), .Z(n14667) );
  AND U15541 ( .A(n14668), .B(n14667), .Z(n14670) );
  XOR U15542 ( .A(n14671), .B(n14670), .Z(c[1612]) );
  NAND U15543 ( .A(n14669), .B(sreg[1612]), .Z(n14673) );
  OR U15544 ( .A(n14671), .B(n14670), .Z(n14672) );
  NAND U15545 ( .A(n14673), .B(n14672), .Z(n14711) );
  NANDN U15546 ( .A(n14675), .B(n14674), .Z(n14679) );
  OR U15547 ( .A(n14677), .B(n14676), .Z(n14678) );
  NAND U15548 ( .A(n14679), .B(n14678), .Z(n14693) );
  AND U15549 ( .A(b[2]), .B(a[591]), .Z(n14702) );
  AND U15550 ( .A(a[592]), .B(b[1]), .Z(n14700) );
  AND U15551 ( .A(a[590]), .B(b[3]), .Z(n14699) );
  XOR U15552 ( .A(n14700), .B(n14699), .Z(n14701) );
  XOR U15553 ( .A(n14702), .B(n14701), .Z(n14705) );
  NAND U15554 ( .A(b[0]), .B(a[593]), .Z(n14706) );
  XNOR U15555 ( .A(n14705), .B(n14706), .Z(n14707) );
  OR U15556 ( .A(n14681), .B(n14680), .Z(n14685) );
  NANDN U15557 ( .A(n14683), .B(n14682), .Z(n14684) );
  AND U15558 ( .A(n14685), .B(n14684), .Z(n14708) );
  XNOR U15559 ( .A(n14707), .B(n14708), .Z(n14694) );
  XNOR U15560 ( .A(n14693), .B(n14694), .Z(n14695) );
  NANDN U15561 ( .A(n14687), .B(n14686), .Z(n14691) );
  NAND U15562 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15563 ( .A(n14691), .B(n14690), .Z(n14696) );
  XNOR U15564 ( .A(n14695), .B(n14696), .Z(n14712) );
  XOR U15565 ( .A(sreg[1613]), .B(n14712), .Z(n14692) );
  XNOR U15566 ( .A(n14711), .B(n14692), .Z(c[1613]) );
  NANDN U15567 ( .A(n14694), .B(n14693), .Z(n14698) );
  NAND U15568 ( .A(n14696), .B(n14695), .Z(n14697) );
  NAND U15569 ( .A(n14698), .B(n14697), .Z(n14719) );
  AND U15570 ( .A(b[2]), .B(a[592]), .Z(n14725) );
  AND U15571 ( .A(a[593]), .B(b[1]), .Z(n14723) );
  AND U15572 ( .A(a[591]), .B(b[3]), .Z(n14722) );
  XOR U15573 ( .A(n14723), .B(n14722), .Z(n14724) );
  XOR U15574 ( .A(n14725), .B(n14724), .Z(n14728) );
  NAND U15575 ( .A(b[0]), .B(a[594]), .Z(n14729) );
  XOR U15576 ( .A(n14728), .B(n14729), .Z(n14731) );
  OR U15577 ( .A(n14700), .B(n14699), .Z(n14704) );
  NANDN U15578 ( .A(n14702), .B(n14701), .Z(n14703) );
  NAND U15579 ( .A(n14704), .B(n14703), .Z(n14730) );
  XNOR U15580 ( .A(n14731), .B(n14730), .Z(n14716) );
  NANDN U15581 ( .A(n14706), .B(n14705), .Z(n14710) );
  NAND U15582 ( .A(n14708), .B(n14707), .Z(n14709) );
  NAND U15583 ( .A(n14710), .B(n14709), .Z(n14717) );
  XNOR U15584 ( .A(n14716), .B(n14717), .Z(n14718) );
  XOR U15585 ( .A(n14719), .B(n14718), .Z(n14715) );
  XNOR U15586 ( .A(sreg[1614]), .B(n14714), .Z(n14713) );
  XNOR U15587 ( .A(n14715), .B(n14713), .Z(c[1614]) );
  NANDN U15588 ( .A(n14717), .B(n14716), .Z(n14721) );
  NANDN U15589 ( .A(n14719), .B(n14718), .Z(n14720) );
  NAND U15590 ( .A(n14721), .B(n14720), .Z(n14754) );
  AND U15591 ( .A(b[2]), .B(a[593]), .Z(n14748) );
  AND U15592 ( .A(a[594]), .B(b[1]), .Z(n14746) );
  AND U15593 ( .A(a[592]), .B(b[3]), .Z(n14745) );
  XOR U15594 ( .A(n14746), .B(n14745), .Z(n14747) );
  XOR U15595 ( .A(n14748), .B(n14747), .Z(n14739) );
  NAND U15596 ( .A(b[0]), .B(a[595]), .Z(n14740) );
  XOR U15597 ( .A(n14739), .B(n14740), .Z(n14742) );
  OR U15598 ( .A(n14723), .B(n14722), .Z(n14727) );
  NANDN U15599 ( .A(n14725), .B(n14724), .Z(n14726) );
  NAND U15600 ( .A(n14727), .B(n14726), .Z(n14741) );
  XNOR U15601 ( .A(n14742), .B(n14741), .Z(n14751) );
  NANDN U15602 ( .A(n14729), .B(n14728), .Z(n14733) );
  OR U15603 ( .A(n14731), .B(n14730), .Z(n14732) );
  NAND U15604 ( .A(n14733), .B(n14732), .Z(n14752) );
  XNOR U15605 ( .A(n14751), .B(n14752), .Z(n14753) );
  XNOR U15606 ( .A(n14754), .B(n14753), .Z(n14734) );
  XNOR U15607 ( .A(n14734), .B(sreg[1615]), .Z(n14735) );
  XOR U15608 ( .A(n14736), .B(n14735), .Z(c[1615]) );
  NAND U15609 ( .A(n14734), .B(sreg[1615]), .Z(n14738) );
  OR U15610 ( .A(n14736), .B(n14735), .Z(n14737) );
  NAND U15611 ( .A(n14738), .B(n14737), .Z(n14758) );
  NANDN U15612 ( .A(n14740), .B(n14739), .Z(n14744) );
  OR U15613 ( .A(n14742), .B(n14741), .Z(n14743) );
  NAND U15614 ( .A(n14744), .B(n14743), .Z(n14760) );
  AND U15615 ( .A(b[2]), .B(a[594]), .Z(n14769) );
  AND U15616 ( .A(a[595]), .B(b[1]), .Z(n14767) );
  AND U15617 ( .A(a[593]), .B(b[3]), .Z(n14766) );
  XOR U15618 ( .A(n14767), .B(n14766), .Z(n14768) );
  XOR U15619 ( .A(n14769), .B(n14768), .Z(n14772) );
  NAND U15620 ( .A(b[0]), .B(a[596]), .Z(n14773) );
  XNOR U15621 ( .A(n14772), .B(n14773), .Z(n14774) );
  OR U15622 ( .A(n14746), .B(n14745), .Z(n14750) );
  NANDN U15623 ( .A(n14748), .B(n14747), .Z(n14749) );
  AND U15624 ( .A(n14750), .B(n14749), .Z(n14775) );
  XNOR U15625 ( .A(n14774), .B(n14775), .Z(n14761) );
  XNOR U15626 ( .A(n14760), .B(n14761), .Z(n14762) );
  NANDN U15627 ( .A(n14752), .B(n14751), .Z(n14756) );
  NAND U15628 ( .A(n14754), .B(n14753), .Z(n14755) );
  AND U15629 ( .A(n14756), .B(n14755), .Z(n14763) );
  XNOR U15630 ( .A(n14762), .B(n14763), .Z(n14759) );
  XOR U15631 ( .A(sreg[1616]), .B(n14759), .Z(n14757) );
  XNOR U15632 ( .A(n14758), .B(n14757), .Z(c[1616]) );
  NANDN U15633 ( .A(n14761), .B(n14760), .Z(n14765) );
  NAND U15634 ( .A(n14763), .B(n14762), .Z(n14764) );
  NAND U15635 ( .A(n14765), .B(n14764), .Z(n14781) );
  AND U15636 ( .A(b[2]), .B(a[595]), .Z(n14787) );
  AND U15637 ( .A(a[596]), .B(b[1]), .Z(n14785) );
  AND U15638 ( .A(a[594]), .B(b[3]), .Z(n14784) );
  XOR U15639 ( .A(n14785), .B(n14784), .Z(n14786) );
  XOR U15640 ( .A(n14787), .B(n14786), .Z(n14790) );
  NAND U15641 ( .A(b[0]), .B(a[597]), .Z(n14791) );
  XOR U15642 ( .A(n14790), .B(n14791), .Z(n14793) );
  OR U15643 ( .A(n14767), .B(n14766), .Z(n14771) );
  NANDN U15644 ( .A(n14769), .B(n14768), .Z(n14770) );
  NAND U15645 ( .A(n14771), .B(n14770), .Z(n14792) );
  XNOR U15646 ( .A(n14793), .B(n14792), .Z(n14778) );
  NANDN U15647 ( .A(n14773), .B(n14772), .Z(n14777) );
  NAND U15648 ( .A(n14775), .B(n14774), .Z(n14776) );
  NAND U15649 ( .A(n14777), .B(n14776), .Z(n14779) );
  XNOR U15650 ( .A(n14778), .B(n14779), .Z(n14780) );
  XOR U15651 ( .A(n14781), .B(n14780), .Z(n14796) );
  XNOR U15652 ( .A(n14796), .B(sreg[1617]), .Z(n14797) );
  XOR U15653 ( .A(n14798), .B(n14797), .Z(c[1617]) );
  NANDN U15654 ( .A(n14779), .B(n14778), .Z(n14783) );
  NANDN U15655 ( .A(n14781), .B(n14780), .Z(n14782) );
  NAND U15656 ( .A(n14783), .B(n14782), .Z(n14807) );
  AND U15657 ( .A(b[2]), .B(a[596]), .Z(n14813) );
  AND U15658 ( .A(a[597]), .B(b[1]), .Z(n14811) );
  AND U15659 ( .A(a[595]), .B(b[3]), .Z(n14810) );
  XOR U15660 ( .A(n14811), .B(n14810), .Z(n14812) );
  XOR U15661 ( .A(n14813), .B(n14812), .Z(n14816) );
  NAND U15662 ( .A(b[0]), .B(a[598]), .Z(n14817) );
  XOR U15663 ( .A(n14816), .B(n14817), .Z(n14819) );
  OR U15664 ( .A(n14785), .B(n14784), .Z(n14789) );
  NANDN U15665 ( .A(n14787), .B(n14786), .Z(n14788) );
  NAND U15666 ( .A(n14789), .B(n14788), .Z(n14818) );
  XNOR U15667 ( .A(n14819), .B(n14818), .Z(n14804) );
  NANDN U15668 ( .A(n14791), .B(n14790), .Z(n14795) );
  OR U15669 ( .A(n14793), .B(n14792), .Z(n14794) );
  NAND U15670 ( .A(n14795), .B(n14794), .Z(n14805) );
  XNOR U15671 ( .A(n14804), .B(n14805), .Z(n14806) );
  XOR U15672 ( .A(n14807), .B(n14806), .Z(n14803) );
  NAND U15673 ( .A(n14796), .B(sreg[1617]), .Z(n14800) );
  OR U15674 ( .A(n14798), .B(n14797), .Z(n14799) );
  NAND U15675 ( .A(n14800), .B(n14799), .Z(n14802) );
  XNOR U15676 ( .A(sreg[1618]), .B(n14802), .Z(n14801) );
  XOR U15677 ( .A(n14803), .B(n14801), .Z(c[1618]) );
  NANDN U15678 ( .A(n14805), .B(n14804), .Z(n14809) );
  NAND U15679 ( .A(n14807), .B(n14806), .Z(n14808) );
  NAND U15680 ( .A(n14809), .B(n14808), .Z(n14830) );
  AND U15681 ( .A(b[2]), .B(a[597]), .Z(n14836) );
  AND U15682 ( .A(a[598]), .B(b[1]), .Z(n14834) );
  AND U15683 ( .A(a[596]), .B(b[3]), .Z(n14833) );
  XOR U15684 ( .A(n14834), .B(n14833), .Z(n14835) );
  XOR U15685 ( .A(n14836), .B(n14835), .Z(n14839) );
  NAND U15686 ( .A(b[0]), .B(a[599]), .Z(n14840) );
  XOR U15687 ( .A(n14839), .B(n14840), .Z(n14842) );
  OR U15688 ( .A(n14811), .B(n14810), .Z(n14815) );
  NANDN U15689 ( .A(n14813), .B(n14812), .Z(n14814) );
  NAND U15690 ( .A(n14815), .B(n14814), .Z(n14841) );
  XNOR U15691 ( .A(n14842), .B(n14841), .Z(n14827) );
  NANDN U15692 ( .A(n14817), .B(n14816), .Z(n14821) );
  OR U15693 ( .A(n14819), .B(n14818), .Z(n14820) );
  NAND U15694 ( .A(n14821), .B(n14820), .Z(n14828) );
  XNOR U15695 ( .A(n14827), .B(n14828), .Z(n14829) );
  XNOR U15696 ( .A(n14830), .B(n14829), .Z(n14822) );
  XOR U15697 ( .A(sreg[1619]), .B(n14822), .Z(n14824) );
  XNOR U15698 ( .A(n14823), .B(n14824), .Z(c[1619]) );
  OR U15699 ( .A(n14822), .B(sreg[1619]), .Z(n14826) );
  NAND U15700 ( .A(n14824), .B(n14823), .Z(n14825) );
  AND U15701 ( .A(n14826), .B(n14825), .Z(n14864) );
  NANDN U15702 ( .A(n14828), .B(n14827), .Z(n14832) );
  NAND U15703 ( .A(n14830), .B(n14829), .Z(n14831) );
  NAND U15704 ( .A(n14832), .B(n14831), .Z(n14849) );
  AND U15705 ( .A(b[2]), .B(a[598]), .Z(n14855) );
  AND U15706 ( .A(a[599]), .B(b[1]), .Z(n14853) );
  AND U15707 ( .A(a[597]), .B(b[3]), .Z(n14852) );
  XOR U15708 ( .A(n14853), .B(n14852), .Z(n14854) );
  XOR U15709 ( .A(n14855), .B(n14854), .Z(n14858) );
  NAND U15710 ( .A(b[0]), .B(a[600]), .Z(n14859) );
  XOR U15711 ( .A(n14858), .B(n14859), .Z(n14861) );
  OR U15712 ( .A(n14834), .B(n14833), .Z(n14838) );
  NANDN U15713 ( .A(n14836), .B(n14835), .Z(n14837) );
  NAND U15714 ( .A(n14838), .B(n14837), .Z(n14860) );
  XNOR U15715 ( .A(n14861), .B(n14860), .Z(n14846) );
  NANDN U15716 ( .A(n14840), .B(n14839), .Z(n14844) );
  OR U15717 ( .A(n14842), .B(n14841), .Z(n14843) );
  NAND U15718 ( .A(n14844), .B(n14843), .Z(n14847) );
  XNOR U15719 ( .A(n14846), .B(n14847), .Z(n14848) );
  XNOR U15720 ( .A(n14849), .B(n14848), .Z(n14865) );
  XOR U15721 ( .A(sreg[1620]), .B(n14865), .Z(n14845) );
  XOR U15722 ( .A(n14864), .B(n14845), .Z(c[1620]) );
  NANDN U15723 ( .A(n14847), .B(n14846), .Z(n14851) );
  NAND U15724 ( .A(n14849), .B(n14848), .Z(n14850) );
  NAND U15725 ( .A(n14851), .B(n14850), .Z(n14870) );
  AND U15726 ( .A(b[2]), .B(a[599]), .Z(n14876) );
  AND U15727 ( .A(a[600]), .B(b[1]), .Z(n14874) );
  AND U15728 ( .A(a[598]), .B(b[3]), .Z(n14873) );
  XOR U15729 ( .A(n14874), .B(n14873), .Z(n14875) );
  XOR U15730 ( .A(n14876), .B(n14875), .Z(n14879) );
  NAND U15731 ( .A(b[0]), .B(a[601]), .Z(n14880) );
  XOR U15732 ( .A(n14879), .B(n14880), .Z(n14882) );
  OR U15733 ( .A(n14853), .B(n14852), .Z(n14857) );
  NANDN U15734 ( .A(n14855), .B(n14854), .Z(n14856) );
  NAND U15735 ( .A(n14857), .B(n14856), .Z(n14881) );
  XNOR U15736 ( .A(n14882), .B(n14881), .Z(n14867) );
  NANDN U15737 ( .A(n14859), .B(n14858), .Z(n14863) );
  OR U15738 ( .A(n14861), .B(n14860), .Z(n14862) );
  NAND U15739 ( .A(n14863), .B(n14862), .Z(n14868) );
  XNOR U15740 ( .A(n14867), .B(n14868), .Z(n14869) );
  XOR U15741 ( .A(n14870), .B(n14869), .Z(n14886) );
  XOR U15742 ( .A(sreg[1621]), .B(n14885), .Z(n14866) );
  XOR U15743 ( .A(n14886), .B(n14866), .Z(c[1621]) );
  NANDN U15744 ( .A(n14868), .B(n14867), .Z(n14872) );
  NAND U15745 ( .A(n14870), .B(n14869), .Z(n14871) );
  NAND U15746 ( .A(n14872), .B(n14871), .Z(n14893) );
  AND U15747 ( .A(b[2]), .B(a[600]), .Z(n14899) );
  AND U15748 ( .A(a[601]), .B(b[1]), .Z(n14897) );
  AND U15749 ( .A(a[599]), .B(b[3]), .Z(n14896) );
  XOR U15750 ( .A(n14897), .B(n14896), .Z(n14898) );
  XOR U15751 ( .A(n14899), .B(n14898), .Z(n14902) );
  NAND U15752 ( .A(b[0]), .B(a[602]), .Z(n14903) );
  XOR U15753 ( .A(n14902), .B(n14903), .Z(n14905) );
  OR U15754 ( .A(n14874), .B(n14873), .Z(n14878) );
  NANDN U15755 ( .A(n14876), .B(n14875), .Z(n14877) );
  NAND U15756 ( .A(n14878), .B(n14877), .Z(n14904) );
  XNOR U15757 ( .A(n14905), .B(n14904), .Z(n14890) );
  NANDN U15758 ( .A(n14880), .B(n14879), .Z(n14884) );
  OR U15759 ( .A(n14882), .B(n14881), .Z(n14883) );
  NAND U15760 ( .A(n14884), .B(n14883), .Z(n14891) );
  XNOR U15761 ( .A(n14890), .B(n14891), .Z(n14892) );
  XOR U15762 ( .A(n14893), .B(n14892), .Z(n14889) );
  XNOR U15763 ( .A(sreg[1622]), .B(n14888), .Z(n14887) );
  XOR U15764 ( .A(n14889), .B(n14887), .Z(c[1622]) );
  NANDN U15765 ( .A(n14891), .B(n14890), .Z(n14895) );
  NAND U15766 ( .A(n14893), .B(n14892), .Z(n14894) );
  NAND U15767 ( .A(n14895), .B(n14894), .Z(n14911) );
  AND U15768 ( .A(b[2]), .B(a[601]), .Z(n14917) );
  AND U15769 ( .A(a[602]), .B(b[1]), .Z(n14915) );
  AND U15770 ( .A(a[600]), .B(b[3]), .Z(n14914) );
  XOR U15771 ( .A(n14915), .B(n14914), .Z(n14916) );
  XOR U15772 ( .A(n14917), .B(n14916), .Z(n14920) );
  NAND U15773 ( .A(b[0]), .B(a[603]), .Z(n14921) );
  XOR U15774 ( .A(n14920), .B(n14921), .Z(n14923) );
  OR U15775 ( .A(n14897), .B(n14896), .Z(n14901) );
  NANDN U15776 ( .A(n14899), .B(n14898), .Z(n14900) );
  NAND U15777 ( .A(n14901), .B(n14900), .Z(n14922) );
  XNOR U15778 ( .A(n14923), .B(n14922), .Z(n14908) );
  NANDN U15779 ( .A(n14903), .B(n14902), .Z(n14907) );
  OR U15780 ( .A(n14905), .B(n14904), .Z(n14906) );
  NAND U15781 ( .A(n14907), .B(n14906), .Z(n14909) );
  XNOR U15782 ( .A(n14908), .B(n14909), .Z(n14910) );
  XNOR U15783 ( .A(n14911), .B(n14910), .Z(n14926) );
  XNOR U15784 ( .A(n14926), .B(sreg[1623]), .Z(n14927) );
  XOR U15785 ( .A(n14928), .B(n14927), .Z(c[1623]) );
  NANDN U15786 ( .A(n14909), .B(n14908), .Z(n14913) );
  NAND U15787 ( .A(n14911), .B(n14910), .Z(n14912) );
  NAND U15788 ( .A(n14913), .B(n14912), .Z(n14935) );
  AND U15789 ( .A(b[2]), .B(a[602]), .Z(n14941) );
  AND U15790 ( .A(a[603]), .B(b[1]), .Z(n14939) );
  AND U15791 ( .A(a[601]), .B(b[3]), .Z(n14938) );
  XOR U15792 ( .A(n14939), .B(n14938), .Z(n14940) );
  XOR U15793 ( .A(n14941), .B(n14940), .Z(n14944) );
  NAND U15794 ( .A(b[0]), .B(a[604]), .Z(n14945) );
  XOR U15795 ( .A(n14944), .B(n14945), .Z(n14947) );
  OR U15796 ( .A(n14915), .B(n14914), .Z(n14919) );
  NANDN U15797 ( .A(n14917), .B(n14916), .Z(n14918) );
  NAND U15798 ( .A(n14919), .B(n14918), .Z(n14946) );
  XNOR U15799 ( .A(n14947), .B(n14946), .Z(n14932) );
  NANDN U15800 ( .A(n14921), .B(n14920), .Z(n14925) );
  OR U15801 ( .A(n14923), .B(n14922), .Z(n14924) );
  NAND U15802 ( .A(n14925), .B(n14924), .Z(n14933) );
  XNOR U15803 ( .A(n14932), .B(n14933), .Z(n14934) );
  XOR U15804 ( .A(n14935), .B(n14934), .Z(n14951) );
  NAND U15805 ( .A(n14926), .B(sreg[1623]), .Z(n14930) );
  OR U15806 ( .A(n14928), .B(n14927), .Z(n14929) );
  NAND U15807 ( .A(n14930), .B(n14929), .Z(n14950) );
  XNOR U15808 ( .A(sreg[1624]), .B(n14950), .Z(n14931) );
  XOR U15809 ( .A(n14951), .B(n14931), .Z(c[1624]) );
  NANDN U15810 ( .A(n14933), .B(n14932), .Z(n14937) );
  NAND U15811 ( .A(n14935), .B(n14934), .Z(n14936) );
  NAND U15812 ( .A(n14937), .B(n14936), .Z(n14956) );
  AND U15813 ( .A(b[2]), .B(a[603]), .Z(n14962) );
  AND U15814 ( .A(a[604]), .B(b[1]), .Z(n14960) );
  AND U15815 ( .A(a[602]), .B(b[3]), .Z(n14959) );
  XOR U15816 ( .A(n14960), .B(n14959), .Z(n14961) );
  XOR U15817 ( .A(n14962), .B(n14961), .Z(n14965) );
  NAND U15818 ( .A(b[0]), .B(a[605]), .Z(n14966) );
  XOR U15819 ( .A(n14965), .B(n14966), .Z(n14968) );
  OR U15820 ( .A(n14939), .B(n14938), .Z(n14943) );
  NANDN U15821 ( .A(n14941), .B(n14940), .Z(n14942) );
  NAND U15822 ( .A(n14943), .B(n14942), .Z(n14967) );
  XNOR U15823 ( .A(n14968), .B(n14967), .Z(n14953) );
  NANDN U15824 ( .A(n14945), .B(n14944), .Z(n14949) );
  OR U15825 ( .A(n14947), .B(n14946), .Z(n14948) );
  NAND U15826 ( .A(n14949), .B(n14948), .Z(n14954) );
  XNOR U15827 ( .A(n14953), .B(n14954), .Z(n14955) );
  XOR U15828 ( .A(n14956), .B(n14955), .Z(n14972) );
  XNOR U15829 ( .A(sreg[1625]), .B(n14971), .Z(n14952) );
  XOR U15830 ( .A(n14972), .B(n14952), .Z(c[1625]) );
  NANDN U15831 ( .A(n14954), .B(n14953), .Z(n14958) );
  NAND U15832 ( .A(n14956), .B(n14955), .Z(n14957) );
  NAND U15833 ( .A(n14958), .B(n14957), .Z(n14979) );
  AND U15834 ( .A(b[2]), .B(a[604]), .Z(n14985) );
  AND U15835 ( .A(a[605]), .B(b[1]), .Z(n14983) );
  AND U15836 ( .A(a[603]), .B(b[3]), .Z(n14982) );
  XOR U15837 ( .A(n14983), .B(n14982), .Z(n14984) );
  XOR U15838 ( .A(n14985), .B(n14984), .Z(n14988) );
  NAND U15839 ( .A(b[0]), .B(a[606]), .Z(n14989) );
  XOR U15840 ( .A(n14988), .B(n14989), .Z(n14991) );
  OR U15841 ( .A(n14960), .B(n14959), .Z(n14964) );
  NANDN U15842 ( .A(n14962), .B(n14961), .Z(n14963) );
  NAND U15843 ( .A(n14964), .B(n14963), .Z(n14990) );
  XNOR U15844 ( .A(n14991), .B(n14990), .Z(n14976) );
  NANDN U15845 ( .A(n14966), .B(n14965), .Z(n14970) );
  OR U15846 ( .A(n14968), .B(n14967), .Z(n14969) );
  NAND U15847 ( .A(n14970), .B(n14969), .Z(n14977) );
  XNOR U15848 ( .A(n14976), .B(n14977), .Z(n14978) );
  XNOR U15849 ( .A(n14979), .B(n14978), .Z(n14975) );
  XOR U15850 ( .A(n14974), .B(sreg[1626]), .Z(n14973) );
  XOR U15851 ( .A(n14975), .B(n14973), .Z(c[1626]) );
  NANDN U15852 ( .A(n14977), .B(n14976), .Z(n14981) );
  NAND U15853 ( .A(n14979), .B(n14978), .Z(n14980) );
  NAND U15854 ( .A(n14981), .B(n14980), .Z(n14997) );
  AND U15855 ( .A(b[2]), .B(a[605]), .Z(n15003) );
  AND U15856 ( .A(a[606]), .B(b[1]), .Z(n15001) );
  AND U15857 ( .A(a[604]), .B(b[3]), .Z(n15000) );
  XOR U15858 ( .A(n15001), .B(n15000), .Z(n15002) );
  XOR U15859 ( .A(n15003), .B(n15002), .Z(n15006) );
  NAND U15860 ( .A(b[0]), .B(a[607]), .Z(n15007) );
  XOR U15861 ( .A(n15006), .B(n15007), .Z(n15009) );
  OR U15862 ( .A(n14983), .B(n14982), .Z(n14987) );
  NANDN U15863 ( .A(n14985), .B(n14984), .Z(n14986) );
  NAND U15864 ( .A(n14987), .B(n14986), .Z(n15008) );
  XNOR U15865 ( .A(n15009), .B(n15008), .Z(n14994) );
  NANDN U15866 ( .A(n14989), .B(n14988), .Z(n14993) );
  OR U15867 ( .A(n14991), .B(n14990), .Z(n14992) );
  NAND U15868 ( .A(n14993), .B(n14992), .Z(n14995) );
  XNOR U15869 ( .A(n14994), .B(n14995), .Z(n14996) );
  XNOR U15870 ( .A(n14997), .B(n14996), .Z(n15012) );
  XNOR U15871 ( .A(n15012), .B(sreg[1627]), .Z(n15014) );
  XNOR U15872 ( .A(n15013), .B(n15014), .Z(c[1627]) );
  NANDN U15873 ( .A(n14995), .B(n14994), .Z(n14999) );
  NAND U15874 ( .A(n14997), .B(n14996), .Z(n14998) );
  NAND U15875 ( .A(n14999), .B(n14998), .Z(n15023) );
  AND U15876 ( .A(b[2]), .B(a[606]), .Z(n15029) );
  AND U15877 ( .A(a[607]), .B(b[1]), .Z(n15027) );
  AND U15878 ( .A(a[605]), .B(b[3]), .Z(n15026) );
  XOR U15879 ( .A(n15027), .B(n15026), .Z(n15028) );
  XOR U15880 ( .A(n15029), .B(n15028), .Z(n15032) );
  NAND U15881 ( .A(b[0]), .B(a[608]), .Z(n15033) );
  XOR U15882 ( .A(n15032), .B(n15033), .Z(n15035) );
  OR U15883 ( .A(n15001), .B(n15000), .Z(n15005) );
  NANDN U15884 ( .A(n15003), .B(n15002), .Z(n15004) );
  NAND U15885 ( .A(n15005), .B(n15004), .Z(n15034) );
  XNOR U15886 ( .A(n15035), .B(n15034), .Z(n15020) );
  NANDN U15887 ( .A(n15007), .B(n15006), .Z(n15011) );
  OR U15888 ( .A(n15009), .B(n15008), .Z(n15010) );
  NAND U15889 ( .A(n15011), .B(n15010), .Z(n15021) );
  XNOR U15890 ( .A(n15020), .B(n15021), .Z(n15022) );
  XOR U15891 ( .A(n15023), .B(n15022), .Z(n15019) );
  NAND U15892 ( .A(n15012), .B(sreg[1627]), .Z(n15016) );
  NANDN U15893 ( .A(n15014), .B(n15013), .Z(n15015) );
  NAND U15894 ( .A(n15016), .B(n15015), .Z(n15018) );
  XNOR U15895 ( .A(sreg[1628]), .B(n15018), .Z(n15017) );
  XOR U15896 ( .A(n15019), .B(n15017), .Z(c[1628]) );
  NANDN U15897 ( .A(n15021), .B(n15020), .Z(n15025) );
  NAND U15898 ( .A(n15023), .B(n15022), .Z(n15024) );
  NAND U15899 ( .A(n15025), .B(n15024), .Z(n15041) );
  AND U15900 ( .A(b[2]), .B(a[607]), .Z(n15047) );
  AND U15901 ( .A(a[608]), .B(b[1]), .Z(n15045) );
  AND U15902 ( .A(a[606]), .B(b[3]), .Z(n15044) );
  XOR U15903 ( .A(n15045), .B(n15044), .Z(n15046) );
  XOR U15904 ( .A(n15047), .B(n15046), .Z(n15050) );
  NAND U15905 ( .A(b[0]), .B(a[609]), .Z(n15051) );
  XOR U15906 ( .A(n15050), .B(n15051), .Z(n15053) );
  OR U15907 ( .A(n15027), .B(n15026), .Z(n15031) );
  NANDN U15908 ( .A(n15029), .B(n15028), .Z(n15030) );
  NAND U15909 ( .A(n15031), .B(n15030), .Z(n15052) );
  XNOR U15910 ( .A(n15053), .B(n15052), .Z(n15038) );
  NANDN U15911 ( .A(n15033), .B(n15032), .Z(n15037) );
  OR U15912 ( .A(n15035), .B(n15034), .Z(n15036) );
  NAND U15913 ( .A(n15037), .B(n15036), .Z(n15039) );
  XNOR U15914 ( .A(n15038), .B(n15039), .Z(n15040) );
  XNOR U15915 ( .A(n15041), .B(n15040), .Z(n15056) );
  XNOR U15916 ( .A(n15056), .B(sreg[1629]), .Z(n15057) );
  XOR U15917 ( .A(n15058), .B(n15057), .Z(c[1629]) );
  NANDN U15918 ( .A(n15039), .B(n15038), .Z(n15043) );
  NAND U15919 ( .A(n15041), .B(n15040), .Z(n15042) );
  NAND U15920 ( .A(n15043), .B(n15042), .Z(n15065) );
  AND U15921 ( .A(b[2]), .B(a[608]), .Z(n15071) );
  AND U15922 ( .A(a[609]), .B(b[1]), .Z(n15069) );
  AND U15923 ( .A(a[607]), .B(b[3]), .Z(n15068) );
  XOR U15924 ( .A(n15069), .B(n15068), .Z(n15070) );
  XOR U15925 ( .A(n15071), .B(n15070), .Z(n15074) );
  NAND U15926 ( .A(b[0]), .B(a[610]), .Z(n15075) );
  XOR U15927 ( .A(n15074), .B(n15075), .Z(n15077) );
  OR U15928 ( .A(n15045), .B(n15044), .Z(n15049) );
  NANDN U15929 ( .A(n15047), .B(n15046), .Z(n15048) );
  NAND U15930 ( .A(n15049), .B(n15048), .Z(n15076) );
  XNOR U15931 ( .A(n15077), .B(n15076), .Z(n15062) );
  NANDN U15932 ( .A(n15051), .B(n15050), .Z(n15055) );
  OR U15933 ( .A(n15053), .B(n15052), .Z(n15054) );
  NAND U15934 ( .A(n15055), .B(n15054), .Z(n15063) );
  XNOR U15935 ( .A(n15062), .B(n15063), .Z(n15064) );
  XOR U15936 ( .A(n15065), .B(n15064), .Z(n15081) );
  NAND U15937 ( .A(n15056), .B(sreg[1629]), .Z(n15060) );
  OR U15938 ( .A(n15058), .B(n15057), .Z(n15059) );
  NAND U15939 ( .A(n15060), .B(n15059), .Z(n15080) );
  XNOR U15940 ( .A(sreg[1630]), .B(n15080), .Z(n15061) );
  XOR U15941 ( .A(n15081), .B(n15061), .Z(c[1630]) );
  NANDN U15942 ( .A(n15063), .B(n15062), .Z(n15067) );
  NAND U15943 ( .A(n15065), .B(n15064), .Z(n15066) );
  NAND U15944 ( .A(n15067), .B(n15066), .Z(n15086) );
  AND U15945 ( .A(b[2]), .B(a[609]), .Z(n15092) );
  AND U15946 ( .A(a[610]), .B(b[1]), .Z(n15090) );
  AND U15947 ( .A(a[608]), .B(b[3]), .Z(n15089) );
  XOR U15948 ( .A(n15090), .B(n15089), .Z(n15091) );
  XOR U15949 ( .A(n15092), .B(n15091), .Z(n15095) );
  NAND U15950 ( .A(b[0]), .B(a[611]), .Z(n15096) );
  XOR U15951 ( .A(n15095), .B(n15096), .Z(n15098) );
  OR U15952 ( .A(n15069), .B(n15068), .Z(n15073) );
  NANDN U15953 ( .A(n15071), .B(n15070), .Z(n15072) );
  NAND U15954 ( .A(n15073), .B(n15072), .Z(n15097) );
  XNOR U15955 ( .A(n15098), .B(n15097), .Z(n15083) );
  NANDN U15956 ( .A(n15075), .B(n15074), .Z(n15079) );
  OR U15957 ( .A(n15077), .B(n15076), .Z(n15078) );
  NAND U15958 ( .A(n15079), .B(n15078), .Z(n15084) );
  XNOR U15959 ( .A(n15083), .B(n15084), .Z(n15085) );
  XOR U15960 ( .A(n15086), .B(n15085), .Z(n15102) );
  XNOR U15961 ( .A(sreg[1631]), .B(n15101), .Z(n15082) );
  XOR U15962 ( .A(n15102), .B(n15082), .Z(c[1631]) );
  NANDN U15963 ( .A(n15084), .B(n15083), .Z(n15088) );
  NAND U15964 ( .A(n15086), .B(n15085), .Z(n15087) );
  NAND U15965 ( .A(n15088), .B(n15087), .Z(n15109) );
  AND U15966 ( .A(b[2]), .B(a[610]), .Z(n15121) );
  AND U15967 ( .A(a[611]), .B(b[1]), .Z(n15119) );
  AND U15968 ( .A(a[609]), .B(b[3]), .Z(n15118) );
  XOR U15969 ( .A(n15119), .B(n15118), .Z(n15120) );
  XOR U15970 ( .A(n15121), .B(n15120), .Z(n15112) );
  NAND U15971 ( .A(b[0]), .B(a[612]), .Z(n15113) );
  XOR U15972 ( .A(n15112), .B(n15113), .Z(n15115) );
  OR U15973 ( .A(n15090), .B(n15089), .Z(n15094) );
  NANDN U15974 ( .A(n15092), .B(n15091), .Z(n15093) );
  NAND U15975 ( .A(n15094), .B(n15093), .Z(n15114) );
  XNOR U15976 ( .A(n15115), .B(n15114), .Z(n15106) );
  NANDN U15977 ( .A(n15096), .B(n15095), .Z(n15100) );
  OR U15978 ( .A(n15098), .B(n15097), .Z(n15099) );
  NAND U15979 ( .A(n15100), .B(n15099), .Z(n15107) );
  XNOR U15980 ( .A(n15106), .B(n15107), .Z(n15108) );
  XNOR U15981 ( .A(n15109), .B(n15108), .Z(n15105) );
  XOR U15982 ( .A(n15104), .B(sreg[1632]), .Z(n15103) );
  XOR U15983 ( .A(n15105), .B(n15103), .Z(c[1632]) );
  NANDN U15984 ( .A(n15107), .B(n15106), .Z(n15111) );
  NAND U15985 ( .A(n15109), .B(n15108), .Z(n15110) );
  NAND U15986 ( .A(n15111), .B(n15110), .Z(n15139) );
  NANDN U15987 ( .A(n15113), .B(n15112), .Z(n15117) );
  OR U15988 ( .A(n15115), .B(n15114), .Z(n15116) );
  NAND U15989 ( .A(n15117), .B(n15116), .Z(n15136) );
  AND U15990 ( .A(b[2]), .B(a[611]), .Z(n15127) );
  AND U15991 ( .A(a[612]), .B(b[1]), .Z(n15125) );
  AND U15992 ( .A(a[610]), .B(b[3]), .Z(n15124) );
  XOR U15993 ( .A(n15125), .B(n15124), .Z(n15126) );
  XOR U15994 ( .A(n15127), .B(n15126), .Z(n15130) );
  NAND U15995 ( .A(b[0]), .B(a[613]), .Z(n15131) );
  XNOR U15996 ( .A(n15130), .B(n15131), .Z(n15132) );
  OR U15997 ( .A(n15119), .B(n15118), .Z(n15123) );
  NANDN U15998 ( .A(n15121), .B(n15120), .Z(n15122) );
  AND U15999 ( .A(n15123), .B(n15122), .Z(n15133) );
  XNOR U16000 ( .A(n15132), .B(n15133), .Z(n15137) );
  XNOR U16001 ( .A(n15136), .B(n15137), .Z(n15138) );
  XNOR U16002 ( .A(n15139), .B(n15138), .Z(n15142) );
  XNOR U16003 ( .A(sreg[1633]), .B(n15142), .Z(n15144) );
  XNOR U16004 ( .A(n15143), .B(n15144), .Z(c[1633]) );
  AND U16005 ( .A(b[2]), .B(a[612]), .Z(n15159) );
  AND U16006 ( .A(a[613]), .B(b[1]), .Z(n15157) );
  AND U16007 ( .A(a[611]), .B(b[3]), .Z(n15156) );
  XOR U16008 ( .A(n15157), .B(n15156), .Z(n15158) );
  XOR U16009 ( .A(n15159), .B(n15158), .Z(n15162) );
  NAND U16010 ( .A(b[0]), .B(a[614]), .Z(n15163) );
  XOR U16011 ( .A(n15162), .B(n15163), .Z(n15165) );
  OR U16012 ( .A(n15125), .B(n15124), .Z(n15129) );
  NANDN U16013 ( .A(n15127), .B(n15126), .Z(n15128) );
  NAND U16014 ( .A(n15129), .B(n15128), .Z(n15164) );
  XNOR U16015 ( .A(n15165), .B(n15164), .Z(n15150) );
  NANDN U16016 ( .A(n15131), .B(n15130), .Z(n15135) );
  NAND U16017 ( .A(n15133), .B(n15132), .Z(n15134) );
  NAND U16018 ( .A(n15135), .B(n15134), .Z(n15151) );
  XNOR U16019 ( .A(n15150), .B(n15151), .Z(n15152) );
  NANDN U16020 ( .A(n15137), .B(n15136), .Z(n15141) );
  NANDN U16021 ( .A(n15139), .B(n15138), .Z(n15140) );
  AND U16022 ( .A(n15141), .B(n15140), .Z(n15153) );
  XNOR U16023 ( .A(n15152), .B(n15153), .Z(n15149) );
  NAND U16024 ( .A(sreg[1633]), .B(n15142), .Z(n15146) );
  NANDN U16025 ( .A(n15144), .B(n15143), .Z(n15145) );
  AND U16026 ( .A(n15146), .B(n15145), .Z(n15148) );
  XNOR U16027 ( .A(n15148), .B(sreg[1634]), .Z(n15147) );
  XOR U16028 ( .A(n15149), .B(n15147), .Z(c[1634]) );
  NANDN U16029 ( .A(n15151), .B(n15150), .Z(n15155) );
  NAND U16030 ( .A(n15153), .B(n15152), .Z(n15154) );
  NAND U16031 ( .A(n15155), .B(n15154), .Z(n15183) );
  AND U16032 ( .A(b[2]), .B(a[613]), .Z(n15177) );
  AND U16033 ( .A(a[614]), .B(b[1]), .Z(n15175) );
  AND U16034 ( .A(a[612]), .B(b[3]), .Z(n15174) );
  XOR U16035 ( .A(n15175), .B(n15174), .Z(n15176) );
  XOR U16036 ( .A(n15177), .B(n15176), .Z(n15168) );
  NAND U16037 ( .A(b[0]), .B(a[615]), .Z(n15169) );
  XOR U16038 ( .A(n15168), .B(n15169), .Z(n15171) );
  OR U16039 ( .A(n15157), .B(n15156), .Z(n15161) );
  NANDN U16040 ( .A(n15159), .B(n15158), .Z(n15160) );
  NAND U16041 ( .A(n15161), .B(n15160), .Z(n15170) );
  XNOR U16042 ( .A(n15171), .B(n15170), .Z(n15180) );
  NANDN U16043 ( .A(n15163), .B(n15162), .Z(n15167) );
  OR U16044 ( .A(n15165), .B(n15164), .Z(n15166) );
  NAND U16045 ( .A(n15167), .B(n15166), .Z(n15181) );
  XNOR U16046 ( .A(n15180), .B(n15181), .Z(n15182) );
  XNOR U16047 ( .A(n15183), .B(n15182), .Z(n15186) );
  XNOR U16048 ( .A(n15186), .B(sreg[1635]), .Z(n15188) );
  XNOR U16049 ( .A(n15187), .B(n15188), .Z(c[1635]) );
  NANDN U16050 ( .A(n15169), .B(n15168), .Z(n15173) );
  OR U16051 ( .A(n15171), .B(n15170), .Z(n15172) );
  NAND U16052 ( .A(n15173), .B(n15172), .Z(n15206) );
  AND U16053 ( .A(b[2]), .B(a[614]), .Z(n15197) );
  AND U16054 ( .A(a[615]), .B(b[1]), .Z(n15195) );
  AND U16055 ( .A(a[613]), .B(b[3]), .Z(n15194) );
  XOR U16056 ( .A(n15195), .B(n15194), .Z(n15196) );
  XOR U16057 ( .A(n15197), .B(n15196), .Z(n15200) );
  NAND U16058 ( .A(b[0]), .B(a[616]), .Z(n15201) );
  XNOR U16059 ( .A(n15200), .B(n15201), .Z(n15202) );
  OR U16060 ( .A(n15175), .B(n15174), .Z(n15179) );
  NANDN U16061 ( .A(n15177), .B(n15176), .Z(n15178) );
  AND U16062 ( .A(n15179), .B(n15178), .Z(n15203) );
  XNOR U16063 ( .A(n15202), .B(n15203), .Z(n15207) );
  XNOR U16064 ( .A(n15206), .B(n15207), .Z(n15208) );
  NANDN U16065 ( .A(n15181), .B(n15180), .Z(n15185) );
  NAND U16066 ( .A(n15183), .B(n15182), .Z(n15184) );
  NAND U16067 ( .A(n15185), .B(n15184), .Z(n15209) );
  XOR U16068 ( .A(n15208), .B(n15209), .Z(n15193) );
  NAND U16069 ( .A(n15186), .B(sreg[1635]), .Z(n15190) );
  NANDN U16070 ( .A(n15188), .B(n15187), .Z(n15189) );
  AND U16071 ( .A(n15190), .B(n15189), .Z(n15192) );
  XNOR U16072 ( .A(n15192), .B(sreg[1636]), .Z(n15191) );
  XNOR U16073 ( .A(n15193), .B(n15191), .Z(c[1636]) );
  AND U16074 ( .A(b[2]), .B(a[615]), .Z(n15221) );
  AND U16075 ( .A(a[616]), .B(b[1]), .Z(n15219) );
  AND U16076 ( .A(a[614]), .B(b[3]), .Z(n15218) );
  XOR U16077 ( .A(n15219), .B(n15218), .Z(n15220) );
  XOR U16078 ( .A(n15221), .B(n15220), .Z(n15224) );
  NAND U16079 ( .A(b[0]), .B(a[617]), .Z(n15225) );
  XOR U16080 ( .A(n15224), .B(n15225), .Z(n15227) );
  OR U16081 ( .A(n15195), .B(n15194), .Z(n15199) );
  NANDN U16082 ( .A(n15197), .B(n15196), .Z(n15198) );
  NAND U16083 ( .A(n15199), .B(n15198), .Z(n15226) );
  XNOR U16084 ( .A(n15227), .B(n15226), .Z(n15212) );
  NANDN U16085 ( .A(n15201), .B(n15200), .Z(n15205) );
  NAND U16086 ( .A(n15203), .B(n15202), .Z(n15204) );
  NAND U16087 ( .A(n15205), .B(n15204), .Z(n15213) );
  XNOR U16088 ( .A(n15212), .B(n15213), .Z(n15214) );
  NANDN U16089 ( .A(n15207), .B(n15206), .Z(n15211) );
  NANDN U16090 ( .A(n15209), .B(n15208), .Z(n15210) );
  NAND U16091 ( .A(n15211), .B(n15210), .Z(n15215) );
  XOR U16092 ( .A(n15214), .B(n15215), .Z(n15230) );
  XNOR U16093 ( .A(n15230), .B(sreg[1637]), .Z(n15232) );
  XNOR U16094 ( .A(n15231), .B(n15232), .Z(c[1637]) );
  NANDN U16095 ( .A(n15213), .B(n15212), .Z(n15217) );
  NANDN U16096 ( .A(n15215), .B(n15214), .Z(n15216) );
  NAND U16097 ( .A(n15217), .B(n15216), .Z(n15255) );
  AND U16098 ( .A(b[2]), .B(a[616]), .Z(n15249) );
  AND U16099 ( .A(a[617]), .B(b[1]), .Z(n15247) );
  AND U16100 ( .A(a[615]), .B(b[3]), .Z(n15246) );
  XOR U16101 ( .A(n15247), .B(n15246), .Z(n15248) );
  XOR U16102 ( .A(n15249), .B(n15248), .Z(n15240) );
  NAND U16103 ( .A(b[0]), .B(a[618]), .Z(n15241) );
  XOR U16104 ( .A(n15240), .B(n15241), .Z(n15243) );
  OR U16105 ( .A(n15219), .B(n15218), .Z(n15223) );
  NANDN U16106 ( .A(n15221), .B(n15220), .Z(n15222) );
  NAND U16107 ( .A(n15223), .B(n15222), .Z(n15242) );
  XNOR U16108 ( .A(n15243), .B(n15242), .Z(n15252) );
  NANDN U16109 ( .A(n15225), .B(n15224), .Z(n15229) );
  OR U16110 ( .A(n15227), .B(n15226), .Z(n15228) );
  NAND U16111 ( .A(n15229), .B(n15228), .Z(n15253) );
  XNOR U16112 ( .A(n15252), .B(n15253), .Z(n15254) );
  XNOR U16113 ( .A(n15255), .B(n15254), .Z(n15235) );
  XNOR U16114 ( .A(n15235), .B(sreg[1638]), .Z(n15237) );
  NAND U16115 ( .A(n15230), .B(sreg[1637]), .Z(n15234) );
  NANDN U16116 ( .A(n15232), .B(n15231), .Z(n15233) );
  AND U16117 ( .A(n15234), .B(n15233), .Z(n15236) );
  XOR U16118 ( .A(n15237), .B(n15236), .Z(c[1638]) );
  NAND U16119 ( .A(n15235), .B(sreg[1638]), .Z(n15239) );
  OR U16120 ( .A(n15237), .B(n15236), .Z(n15238) );
  NAND U16121 ( .A(n15239), .B(n15238), .Z(n15260) );
  NANDN U16122 ( .A(n15241), .B(n15240), .Z(n15245) );
  OR U16123 ( .A(n15243), .B(n15242), .Z(n15244) );
  NAND U16124 ( .A(n15245), .B(n15244), .Z(n15275) );
  AND U16125 ( .A(b[2]), .B(a[617]), .Z(n15266) );
  AND U16126 ( .A(a[618]), .B(b[1]), .Z(n15264) );
  AND U16127 ( .A(a[616]), .B(b[3]), .Z(n15263) );
  XOR U16128 ( .A(n15264), .B(n15263), .Z(n15265) );
  XOR U16129 ( .A(n15266), .B(n15265), .Z(n15269) );
  NAND U16130 ( .A(b[0]), .B(a[619]), .Z(n15270) );
  XNOR U16131 ( .A(n15269), .B(n15270), .Z(n15271) );
  OR U16132 ( .A(n15247), .B(n15246), .Z(n15251) );
  NANDN U16133 ( .A(n15249), .B(n15248), .Z(n15250) );
  AND U16134 ( .A(n15251), .B(n15250), .Z(n15272) );
  XNOR U16135 ( .A(n15271), .B(n15272), .Z(n15276) );
  XNOR U16136 ( .A(n15275), .B(n15276), .Z(n15277) );
  NANDN U16137 ( .A(n15253), .B(n15252), .Z(n15257) );
  NAND U16138 ( .A(n15255), .B(n15254), .Z(n15256) );
  NAND U16139 ( .A(n15257), .B(n15256), .Z(n15278) );
  XNOR U16140 ( .A(n15277), .B(n15278), .Z(n15258) );
  XOR U16141 ( .A(sreg[1639]), .B(n15258), .Z(n15259) );
  XOR U16142 ( .A(n15260), .B(n15259), .Z(c[1639]) );
  OR U16143 ( .A(n15258), .B(sreg[1639]), .Z(n15262) );
  NANDN U16144 ( .A(n15260), .B(n15259), .Z(n15261) );
  NAND U16145 ( .A(n15262), .B(n15261), .Z(n15301) );
  AND U16146 ( .A(b[2]), .B(a[618]), .Z(n15290) );
  AND U16147 ( .A(a[619]), .B(b[1]), .Z(n15288) );
  AND U16148 ( .A(a[617]), .B(b[3]), .Z(n15287) );
  XOR U16149 ( .A(n15288), .B(n15287), .Z(n15289) );
  XOR U16150 ( .A(n15290), .B(n15289), .Z(n15293) );
  NAND U16151 ( .A(b[0]), .B(a[620]), .Z(n15294) );
  XOR U16152 ( .A(n15293), .B(n15294), .Z(n15296) );
  OR U16153 ( .A(n15264), .B(n15263), .Z(n15268) );
  NANDN U16154 ( .A(n15266), .B(n15265), .Z(n15267) );
  NAND U16155 ( .A(n15268), .B(n15267), .Z(n15295) );
  XNOR U16156 ( .A(n15296), .B(n15295), .Z(n15281) );
  NANDN U16157 ( .A(n15270), .B(n15269), .Z(n15274) );
  NAND U16158 ( .A(n15272), .B(n15271), .Z(n15273) );
  NAND U16159 ( .A(n15274), .B(n15273), .Z(n15282) );
  XNOR U16160 ( .A(n15281), .B(n15282), .Z(n15283) );
  NANDN U16161 ( .A(n15276), .B(n15275), .Z(n15280) );
  NANDN U16162 ( .A(n15278), .B(n15277), .Z(n15279) );
  NAND U16163 ( .A(n15280), .B(n15279), .Z(n15284) );
  XOR U16164 ( .A(n15283), .B(n15284), .Z(n15299) );
  XNOR U16165 ( .A(n15299), .B(sreg[1640]), .Z(n15300) );
  XOR U16166 ( .A(n15301), .B(n15300), .Z(c[1640]) );
  NANDN U16167 ( .A(n15282), .B(n15281), .Z(n15286) );
  NANDN U16168 ( .A(n15284), .B(n15283), .Z(n15285) );
  NAND U16169 ( .A(n15286), .B(n15285), .Z(n15324) );
  AND U16170 ( .A(b[2]), .B(a[619]), .Z(n15318) );
  AND U16171 ( .A(a[620]), .B(b[1]), .Z(n15316) );
  AND U16172 ( .A(a[618]), .B(b[3]), .Z(n15315) );
  XOR U16173 ( .A(n15316), .B(n15315), .Z(n15317) );
  XOR U16174 ( .A(n15318), .B(n15317), .Z(n15309) );
  NAND U16175 ( .A(b[0]), .B(a[621]), .Z(n15310) );
  XOR U16176 ( .A(n15309), .B(n15310), .Z(n15312) );
  OR U16177 ( .A(n15288), .B(n15287), .Z(n15292) );
  NANDN U16178 ( .A(n15290), .B(n15289), .Z(n15291) );
  NAND U16179 ( .A(n15292), .B(n15291), .Z(n15311) );
  XNOR U16180 ( .A(n15312), .B(n15311), .Z(n15321) );
  NANDN U16181 ( .A(n15294), .B(n15293), .Z(n15298) );
  OR U16182 ( .A(n15296), .B(n15295), .Z(n15297) );
  NAND U16183 ( .A(n15298), .B(n15297), .Z(n15322) );
  XNOR U16184 ( .A(n15321), .B(n15322), .Z(n15323) );
  XNOR U16185 ( .A(n15324), .B(n15323), .Z(n15304) );
  XNOR U16186 ( .A(n15304), .B(sreg[1641]), .Z(n15306) );
  NAND U16187 ( .A(n15299), .B(sreg[1640]), .Z(n15303) );
  OR U16188 ( .A(n15301), .B(n15300), .Z(n15302) );
  AND U16189 ( .A(n15303), .B(n15302), .Z(n15305) );
  XOR U16190 ( .A(n15306), .B(n15305), .Z(c[1641]) );
  NAND U16191 ( .A(n15304), .B(sreg[1641]), .Z(n15308) );
  OR U16192 ( .A(n15306), .B(n15305), .Z(n15307) );
  NAND U16193 ( .A(n15308), .B(n15307), .Z(n15346) );
  NANDN U16194 ( .A(n15310), .B(n15309), .Z(n15314) );
  OR U16195 ( .A(n15312), .B(n15311), .Z(n15313) );
  NAND U16196 ( .A(n15314), .B(n15313), .Z(n15328) );
  AND U16197 ( .A(b[2]), .B(a[620]), .Z(n15337) );
  AND U16198 ( .A(a[621]), .B(b[1]), .Z(n15335) );
  AND U16199 ( .A(a[619]), .B(b[3]), .Z(n15334) );
  XOR U16200 ( .A(n15335), .B(n15334), .Z(n15336) );
  XOR U16201 ( .A(n15337), .B(n15336), .Z(n15340) );
  NAND U16202 ( .A(b[0]), .B(a[622]), .Z(n15341) );
  XNOR U16203 ( .A(n15340), .B(n15341), .Z(n15342) );
  OR U16204 ( .A(n15316), .B(n15315), .Z(n15320) );
  NANDN U16205 ( .A(n15318), .B(n15317), .Z(n15319) );
  AND U16206 ( .A(n15320), .B(n15319), .Z(n15343) );
  XNOR U16207 ( .A(n15342), .B(n15343), .Z(n15329) );
  XNOR U16208 ( .A(n15328), .B(n15329), .Z(n15330) );
  NANDN U16209 ( .A(n15322), .B(n15321), .Z(n15326) );
  NAND U16210 ( .A(n15324), .B(n15323), .Z(n15325) );
  AND U16211 ( .A(n15326), .B(n15325), .Z(n15331) );
  XNOR U16212 ( .A(n15330), .B(n15331), .Z(n15347) );
  XOR U16213 ( .A(sreg[1642]), .B(n15347), .Z(n15327) );
  XNOR U16214 ( .A(n15346), .B(n15327), .Z(c[1642]) );
  NANDN U16215 ( .A(n15329), .B(n15328), .Z(n15333) );
  NAND U16216 ( .A(n15331), .B(n15330), .Z(n15332) );
  NAND U16217 ( .A(n15333), .B(n15332), .Z(n15354) );
  AND U16218 ( .A(b[2]), .B(a[621]), .Z(n15360) );
  AND U16219 ( .A(a[622]), .B(b[1]), .Z(n15358) );
  AND U16220 ( .A(a[620]), .B(b[3]), .Z(n15357) );
  XOR U16221 ( .A(n15358), .B(n15357), .Z(n15359) );
  XOR U16222 ( .A(n15360), .B(n15359), .Z(n15363) );
  NAND U16223 ( .A(b[0]), .B(a[623]), .Z(n15364) );
  XOR U16224 ( .A(n15363), .B(n15364), .Z(n15366) );
  OR U16225 ( .A(n15335), .B(n15334), .Z(n15339) );
  NANDN U16226 ( .A(n15337), .B(n15336), .Z(n15338) );
  NAND U16227 ( .A(n15339), .B(n15338), .Z(n15365) );
  XNOR U16228 ( .A(n15366), .B(n15365), .Z(n15351) );
  NANDN U16229 ( .A(n15341), .B(n15340), .Z(n15345) );
  NAND U16230 ( .A(n15343), .B(n15342), .Z(n15344) );
  NAND U16231 ( .A(n15345), .B(n15344), .Z(n15352) );
  XNOR U16232 ( .A(n15351), .B(n15352), .Z(n15353) );
  XNOR U16233 ( .A(n15354), .B(n15353), .Z(n15350) );
  XOR U16234 ( .A(n15349), .B(sreg[1643]), .Z(n15348) );
  XNOR U16235 ( .A(n15350), .B(n15348), .Z(c[1643]) );
  NANDN U16236 ( .A(n15352), .B(n15351), .Z(n15356) );
  NANDN U16237 ( .A(n15354), .B(n15353), .Z(n15355) );
  NAND U16238 ( .A(n15356), .B(n15355), .Z(n15377) );
  AND U16239 ( .A(b[2]), .B(a[622]), .Z(n15383) );
  AND U16240 ( .A(a[623]), .B(b[1]), .Z(n15381) );
  AND U16241 ( .A(a[621]), .B(b[3]), .Z(n15380) );
  XOR U16242 ( .A(n15381), .B(n15380), .Z(n15382) );
  XOR U16243 ( .A(n15383), .B(n15382), .Z(n15386) );
  NAND U16244 ( .A(b[0]), .B(a[624]), .Z(n15387) );
  XOR U16245 ( .A(n15386), .B(n15387), .Z(n15389) );
  OR U16246 ( .A(n15358), .B(n15357), .Z(n15362) );
  NANDN U16247 ( .A(n15360), .B(n15359), .Z(n15361) );
  NAND U16248 ( .A(n15362), .B(n15361), .Z(n15388) );
  XNOR U16249 ( .A(n15389), .B(n15388), .Z(n15374) );
  NANDN U16250 ( .A(n15364), .B(n15363), .Z(n15368) );
  OR U16251 ( .A(n15366), .B(n15365), .Z(n15367) );
  NAND U16252 ( .A(n15368), .B(n15367), .Z(n15375) );
  XNOR U16253 ( .A(n15374), .B(n15375), .Z(n15376) );
  XNOR U16254 ( .A(n15377), .B(n15376), .Z(n15369) );
  XOR U16255 ( .A(sreg[1644]), .B(n15369), .Z(n15370) );
  XOR U16256 ( .A(n15371), .B(n15370), .Z(c[1644]) );
  OR U16257 ( .A(n15369), .B(sreg[1644]), .Z(n15373) );
  NANDN U16258 ( .A(n15371), .B(n15370), .Z(n15372) );
  AND U16259 ( .A(n15373), .B(n15372), .Z(n15411) );
  NANDN U16260 ( .A(n15375), .B(n15374), .Z(n15379) );
  NAND U16261 ( .A(n15377), .B(n15376), .Z(n15378) );
  NAND U16262 ( .A(n15379), .B(n15378), .Z(n15396) );
  AND U16263 ( .A(b[2]), .B(a[623]), .Z(n15402) );
  AND U16264 ( .A(a[624]), .B(b[1]), .Z(n15400) );
  AND U16265 ( .A(a[622]), .B(b[3]), .Z(n15399) );
  XOR U16266 ( .A(n15400), .B(n15399), .Z(n15401) );
  XOR U16267 ( .A(n15402), .B(n15401), .Z(n15405) );
  NAND U16268 ( .A(b[0]), .B(a[625]), .Z(n15406) );
  XOR U16269 ( .A(n15405), .B(n15406), .Z(n15408) );
  OR U16270 ( .A(n15381), .B(n15380), .Z(n15385) );
  NANDN U16271 ( .A(n15383), .B(n15382), .Z(n15384) );
  NAND U16272 ( .A(n15385), .B(n15384), .Z(n15407) );
  XNOR U16273 ( .A(n15408), .B(n15407), .Z(n15393) );
  NANDN U16274 ( .A(n15387), .B(n15386), .Z(n15391) );
  OR U16275 ( .A(n15389), .B(n15388), .Z(n15390) );
  NAND U16276 ( .A(n15391), .B(n15390), .Z(n15394) );
  XNOR U16277 ( .A(n15393), .B(n15394), .Z(n15395) );
  XNOR U16278 ( .A(n15396), .B(n15395), .Z(n15412) );
  XOR U16279 ( .A(sreg[1645]), .B(n15412), .Z(n15392) );
  XOR U16280 ( .A(n15411), .B(n15392), .Z(c[1645]) );
  NANDN U16281 ( .A(n15394), .B(n15393), .Z(n15398) );
  NAND U16282 ( .A(n15396), .B(n15395), .Z(n15397) );
  NAND U16283 ( .A(n15398), .B(n15397), .Z(n15417) );
  AND U16284 ( .A(b[2]), .B(a[624]), .Z(n15423) );
  AND U16285 ( .A(a[625]), .B(b[1]), .Z(n15421) );
  AND U16286 ( .A(a[623]), .B(b[3]), .Z(n15420) );
  XOR U16287 ( .A(n15421), .B(n15420), .Z(n15422) );
  XOR U16288 ( .A(n15423), .B(n15422), .Z(n15426) );
  NAND U16289 ( .A(b[0]), .B(a[626]), .Z(n15427) );
  XOR U16290 ( .A(n15426), .B(n15427), .Z(n15429) );
  OR U16291 ( .A(n15400), .B(n15399), .Z(n15404) );
  NANDN U16292 ( .A(n15402), .B(n15401), .Z(n15403) );
  NAND U16293 ( .A(n15404), .B(n15403), .Z(n15428) );
  XNOR U16294 ( .A(n15429), .B(n15428), .Z(n15414) );
  NANDN U16295 ( .A(n15406), .B(n15405), .Z(n15410) );
  OR U16296 ( .A(n15408), .B(n15407), .Z(n15409) );
  NAND U16297 ( .A(n15410), .B(n15409), .Z(n15415) );
  XNOR U16298 ( .A(n15414), .B(n15415), .Z(n15416) );
  XNOR U16299 ( .A(n15417), .B(n15416), .Z(n15432) );
  XNOR U16300 ( .A(sreg[1646]), .B(n15433), .Z(n15413) );
  XNOR U16301 ( .A(n15432), .B(n15413), .Z(c[1646]) );
  NANDN U16302 ( .A(n15415), .B(n15414), .Z(n15419) );
  NAND U16303 ( .A(n15417), .B(n15416), .Z(n15418) );
  NAND U16304 ( .A(n15419), .B(n15418), .Z(n15440) );
  AND U16305 ( .A(b[2]), .B(a[625]), .Z(n15446) );
  AND U16306 ( .A(a[626]), .B(b[1]), .Z(n15444) );
  AND U16307 ( .A(a[624]), .B(b[3]), .Z(n15443) );
  XOR U16308 ( .A(n15444), .B(n15443), .Z(n15445) );
  XOR U16309 ( .A(n15446), .B(n15445), .Z(n15449) );
  NAND U16310 ( .A(b[0]), .B(a[627]), .Z(n15450) );
  XOR U16311 ( .A(n15449), .B(n15450), .Z(n15452) );
  OR U16312 ( .A(n15421), .B(n15420), .Z(n15425) );
  NANDN U16313 ( .A(n15423), .B(n15422), .Z(n15424) );
  NAND U16314 ( .A(n15425), .B(n15424), .Z(n15451) );
  XNOR U16315 ( .A(n15452), .B(n15451), .Z(n15437) );
  NANDN U16316 ( .A(n15427), .B(n15426), .Z(n15431) );
  OR U16317 ( .A(n15429), .B(n15428), .Z(n15430) );
  NAND U16318 ( .A(n15431), .B(n15430), .Z(n15438) );
  XNOR U16319 ( .A(n15437), .B(n15438), .Z(n15439) );
  XOR U16320 ( .A(n15440), .B(n15439), .Z(n15436) );
  XNOR U16321 ( .A(sreg[1647]), .B(n15435), .Z(n15434) );
  XOR U16322 ( .A(n15436), .B(n15434), .Z(c[1647]) );
  NANDN U16323 ( .A(n15438), .B(n15437), .Z(n15442) );
  NAND U16324 ( .A(n15440), .B(n15439), .Z(n15441) );
  NAND U16325 ( .A(n15442), .B(n15441), .Z(n15458) );
  AND U16326 ( .A(b[2]), .B(a[626]), .Z(n15464) );
  AND U16327 ( .A(a[627]), .B(b[1]), .Z(n15462) );
  AND U16328 ( .A(a[625]), .B(b[3]), .Z(n15461) );
  XOR U16329 ( .A(n15462), .B(n15461), .Z(n15463) );
  XOR U16330 ( .A(n15464), .B(n15463), .Z(n15467) );
  NAND U16331 ( .A(b[0]), .B(a[628]), .Z(n15468) );
  XOR U16332 ( .A(n15467), .B(n15468), .Z(n15470) );
  OR U16333 ( .A(n15444), .B(n15443), .Z(n15448) );
  NANDN U16334 ( .A(n15446), .B(n15445), .Z(n15447) );
  NAND U16335 ( .A(n15448), .B(n15447), .Z(n15469) );
  XNOR U16336 ( .A(n15470), .B(n15469), .Z(n15455) );
  NANDN U16337 ( .A(n15450), .B(n15449), .Z(n15454) );
  OR U16338 ( .A(n15452), .B(n15451), .Z(n15453) );
  NAND U16339 ( .A(n15454), .B(n15453), .Z(n15456) );
  XNOR U16340 ( .A(n15455), .B(n15456), .Z(n15457) );
  XNOR U16341 ( .A(n15458), .B(n15457), .Z(n15473) );
  XOR U16342 ( .A(sreg[1648]), .B(n15473), .Z(n15475) );
  XNOR U16343 ( .A(n15474), .B(n15475), .Z(c[1648]) );
  NANDN U16344 ( .A(n15456), .B(n15455), .Z(n15460) );
  NAND U16345 ( .A(n15458), .B(n15457), .Z(n15459) );
  NAND U16346 ( .A(n15460), .B(n15459), .Z(n15482) );
  AND U16347 ( .A(b[2]), .B(a[627]), .Z(n15488) );
  AND U16348 ( .A(a[628]), .B(b[1]), .Z(n15486) );
  AND U16349 ( .A(a[626]), .B(b[3]), .Z(n15485) );
  XOR U16350 ( .A(n15486), .B(n15485), .Z(n15487) );
  XOR U16351 ( .A(n15488), .B(n15487), .Z(n15491) );
  NAND U16352 ( .A(b[0]), .B(a[629]), .Z(n15492) );
  XOR U16353 ( .A(n15491), .B(n15492), .Z(n15494) );
  OR U16354 ( .A(n15462), .B(n15461), .Z(n15466) );
  NANDN U16355 ( .A(n15464), .B(n15463), .Z(n15465) );
  NAND U16356 ( .A(n15466), .B(n15465), .Z(n15493) );
  XNOR U16357 ( .A(n15494), .B(n15493), .Z(n15479) );
  NANDN U16358 ( .A(n15468), .B(n15467), .Z(n15472) );
  OR U16359 ( .A(n15470), .B(n15469), .Z(n15471) );
  NAND U16360 ( .A(n15472), .B(n15471), .Z(n15480) );
  XNOR U16361 ( .A(n15479), .B(n15480), .Z(n15481) );
  XOR U16362 ( .A(n15482), .B(n15481), .Z(n15498) );
  OR U16363 ( .A(n15473), .B(sreg[1648]), .Z(n15477) );
  NAND U16364 ( .A(n15475), .B(n15474), .Z(n15476) );
  AND U16365 ( .A(n15477), .B(n15476), .Z(n15497) );
  XNOR U16366 ( .A(sreg[1649]), .B(n15497), .Z(n15478) );
  XOR U16367 ( .A(n15498), .B(n15478), .Z(c[1649]) );
  NANDN U16368 ( .A(n15480), .B(n15479), .Z(n15484) );
  NAND U16369 ( .A(n15482), .B(n15481), .Z(n15483) );
  NAND U16370 ( .A(n15484), .B(n15483), .Z(n15505) );
  AND U16371 ( .A(b[2]), .B(a[628]), .Z(n15511) );
  AND U16372 ( .A(a[629]), .B(b[1]), .Z(n15509) );
  AND U16373 ( .A(a[627]), .B(b[3]), .Z(n15508) );
  XOR U16374 ( .A(n15509), .B(n15508), .Z(n15510) );
  XOR U16375 ( .A(n15511), .B(n15510), .Z(n15514) );
  NAND U16376 ( .A(b[0]), .B(a[630]), .Z(n15515) );
  XOR U16377 ( .A(n15514), .B(n15515), .Z(n15517) );
  OR U16378 ( .A(n15486), .B(n15485), .Z(n15490) );
  NANDN U16379 ( .A(n15488), .B(n15487), .Z(n15489) );
  NAND U16380 ( .A(n15490), .B(n15489), .Z(n15516) );
  XNOR U16381 ( .A(n15517), .B(n15516), .Z(n15502) );
  NANDN U16382 ( .A(n15492), .B(n15491), .Z(n15496) );
  OR U16383 ( .A(n15494), .B(n15493), .Z(n15495) );
  NAND U16384 ( .A(n15496), .B(n15495), .Z(n15503) );
  XNOR U16385 ( .A(n15502), .B(n15503), .Z(n15504) );
  XNOR U16386 ( .A(n15505), .B(n15504), .Z(n15501) );
  XOR U16387 ( .A(n15500), .B(sreg[1650]), .Z(n15499) );
  XOR U16388 ( .A(n15501), .B(n15499), .Z(c[1650]) );
  NANDN U16389 ( .A(n15503), .B(n15502), .Z(n15507) );
  NAND U16390 ( .A(n15505), .B(n15504), .Z(n15506) );
  NAND U16391 ( .A(n15507), .B(n15506), .Z(n15523) );
  AND U16392 ( .A(b[2]), .B(a[629]), .Z(n15529) );
  AND U16393 ( .A(a[630]), .B(b[1]), .Z(n15527) );
  AND U16394 ( .A(a[628]), .B(b[3]), .Z(n15526) );
  XOR U16395 ( .A(n15527), .B(n15526), .Z(n15528) );
  XOR U16396 ( .A(n15529), .B(n15528), .Z(n15532) );
  NAND U16397 ( .A(b[0]), .B(a[631]), .Z(n15533) );
  XOR U16398 ( .A(n15532), .B(n15533), .Z(n15535) );
  OR U16399 ( .A(n15509), .B(n15508), .Z(n15513) );
  NANDN U16400 ( .A(n15511), .B(n15510), .Z(n15512) );
  NAND U16401 ( .A(n15513), .B(n15512), .Z(n15534) );
  XNOR U16402 ( .A(n15535), .B(n15534), .Z(n15520) );
  NANDN U16403 ( .A(n15515), .B(n15514), .Z(n15519) );
  OR U16404 ( .A(n15517), .B(n15516), .Z(n15518) );
  NAND U16405 ( .A(n15519), .B(n15518), .Z(n15521) );
  XNOR U16406 ( .A(n15520), .B(n15521), .Z(n15522) );
  XNOR U16407 ( .A(n15523), .B(n15522), .Z(n15538) );
  XNOR U16408 ( .A(n15538), .B(sreg[1651]), .Z(n15540) );
  XNOR U16409 ( .A(n15539), .B(n15540), .Z(c[1651]) );
  NANDN U16410 ( .A(n15521), .B(n15520), .Z(n15525) );
  NAND U16411 ( .A(n15523), .B(n15522), .Z(n15524) );
  NAND U16412 ( .A(n15525), .B(n15524), .Z(n15546) );
  AND U16413 ( .A(b[2]), .B(a[630]), .Z(n15552) );
  AND U16414 ( .A(a[631]), .B(b[1]), .Z(n15550) );
  AND U16415 ( .A(a[629]), .B(b[3]), .Z(n15549) );
  XOR U16416 ( .A(n15550), .B(n15549), .Z(n15551) );
  XOR U16417 ( .A(n15552), .B(n15551), .Z(n15555) );
  NAND U16418 ( .A(b[0]), .B(a[632]), .Z(n15556) );
  XOR U16419 ( .A(n15555), .B(n15556), .Z(n15558) );
  OR U16420 ( .A(n15527), .B(n15526), .Z(n15531) );
  NANDN U16421 ( .A(n15529), .B(n15528), .Z(n15530) );
  NAND U16422 ( .A(n15531), .B(n15530), .Z(n15557) );
  XNOR U16423 ( .A(n15558), .B(n15557), .Z(n15543) );
  NANDN U16424 ( .A(n15533), .B(n15532), .Z(n15537) );
  OR U16425 ( .A(n15535), .B(n15534), .Z(n15536) );
  NAND U16426 ( .A(n15537), .B(n15536), .Z(n15544) );
  XNOR U16427 ( .A(n15543), .B(n15544), .Z(n15545) );
  XNOR U16428 ( .A(n15546), .B(n15545), .Z(n15561) );
  XNOR U16429 ( .A(n15561), .B(sreg[1652]), .Z(n15563) );
  NAND U16430 ( .A(n15538), .B(sreg[1651]), .Z(n15542) );
  NANDN U16431 ( .A(n15540), .B(n15539), .Z(n15541) );
  AND U16432 ( .A(n15542), .B(n15541), .Z(n15562) );
  XOR U16433 ( .A(n15563), .B(n15562), .Z(c[1652]) );
  NANDN U16434 ( .A(n15544), .B(n15543), .Z(n15548) );
  NAND U16435 ( .A(n15546), .B(n15545), .Z(n15547) );
  NAND U16436 ( .A(n15548), .B(n15547), .Z(n15572) );
  AND U16437 ( .A(b[2]), .B(a[631]), .Z(n15578) );
  AND U16438 ( .A(a[632]), .B(b[1]), .Z(n15576) );
  AND U16439 ( .A(a[630]), .B(b[3]), .Z(n15575) );
  XOR U16440 ( .A(n15576), .B(n15575), .Z(n15577) );
  XOR U16441 ( .A(n15578), .B(n15577), .Z(n15581) );
  NAND U16442 ( .A(b[0]), .B(a[633]), .Z(n15582) );
  XOR U16443 ( .A(n15581), .B(n15582), .Z(n15584) );
  OR U16444 ( .A(n15550), .B(n15549), .Z(n15554) );
  NANDN U16445 ( .A(n15552), .B(n15551), .Z(n15553) );
  NAND U16446 ( .A(n15554), .B(n15553), .Z(n15583) );
  XNOR U16447 ( .A(n15584), .B(n15583), .Z(n15569) );
  NANDN U16448 ( .A(n15556), .B(n15555), .Z(n15560) );
  OR U16449 ( .A(n15558), .B(n15557), .Z(n15559) );
  NAND U16450 ( .A(n15560), .B(n15559), .Z(n15570) );
  XNOR U16451 ( .A(n15569), .B(n15570), .Z(n15571) );
  XOR U16452 ( .A(n15572), .B(n15571), .Z(n15568) );
  NAND U16453 ( .A(n15561), .B(sreg[1652]), .Z(n15565) );
  OR U16454 ( .A(n15563), .B(n15562), .Z(n15564) );
  NAND U16455 ( .A(n15565), .B(n15564), .Z(n15567) );
  XNOR U16456 ( .A(sreg[1653]), .B(n15567), .Z(n15566) );
  XOR U16457 ( .A(n15568), .B(n15566), .Z(c[1653]) );
  NANDN U16458 ( .A(n15570), .B(n15569), .Z(n15574) );
  NAND U16459 ( .A(n15572), .B(n15571), .Z(n15573) );
  NAND U16460 ( .A(n15574), .B(n15573), .Z(n15590) );
  AND U16461 ( .A(b[2]), .B(a[632]), .Z(n15596) );
  AND U16462 ( .A(a[633]), .B(b[1]), .Z(n15594) );
  AND U16463 ( .A(a[631]), .B(b[3]), .Z(n15593) );
  XOR U16464 ( .A(n15594), .B(n15593), .Z(n15595) );
  XOR U16465 ( .A(n15596), .B(n15595), .Z(n15599) );
  NAND U16466 ( .A(b[0]), .B(a[634]), .Z(n15600) );
  XOR U16467 ( .A(n15599), .B(n15600), .Z(n15602) );
  OR U16468 ( .A(n15576), .B(n15575), .Z(n15580) );
  NANDN U16469 ( .A(n15578), .B(n15577), .Z(n15579) );
  NAND U16470 ( .A(n15580), .B(n15579), .Z(n15601) );
  XNOR U16471 ( .A(n15602), .B(n15601), .Z(n15587) );
  NANDN U16472 ( .A(n15582), .B(n15581), .Z(n15586) );
  OR U16473 ( .A(n15584), .B(n15583), .Z(n15585) );
  NAND U16474 ( .A(n15586), .B(n15585), .Z(n15588) );
  XNOR U16475 ( .A(n15587), .B(n15588), .Z(n15589) );
  XNOR U16476 ( .A(n15590), .B(n15589), .Z(n15605) );
  XNOR U16477 ( .A(n15605), .B(sreg[1654]), .Z(n15606) );
  XOR U16478 ( .A(n15607), .B(n15606), .Z(c[1654]) );
  NANDN U16479 ( .A(n15588), .B(n15587), .Z(n15592) );
  NAND U16480 ( .A(n15590), .B(n15589), .Z(n15591) );
  NAND U16481 ( .A(n15592), .B(n15591), .Z(n15614) );
  AND U16482 ( .A(b[2]), .B(a[633]), .Z(n15620) );
  AND U16483 ( .A(a[634]), .B(b[1]), .Z(n15618) );
  AND U16484 ( .A(a[632]), .B(b[3]), .Z(n15617) );
  XOR U16485 ( .A(n15618), .B(n15617), .Z(n15619) );
  XOR U16486 ( .A(n15620), .B(n15619), .Z(n15623) );
  NAND U16487 ( .A(b[0]), .B(a[635]), .Z(n15624) );
  XOR U16488 ( .A(n15623), .B(n15624), .Z(n15626) );
  OR U16489 ( .A(n15594), .B(n15593), .Z(n15598) );
  NANDN U16490 ( .A(n15596), .B(n15595), .Z(n15597) );
  NAND U16491 ( .A(n15598), .B(n15597), .Z(n15625) );
  XNOR U16492 ( .A(n15626), .B(n15625), .Z(n15611) );
  NANDN U16493 ( .A(n15600), .B(n15599), .Z(n15604) );
  OR U16494 ( .A(n15602), .B(n15601), .Z(n15603) );
  NAND U16495 ( .A(n15604), .B(n15603), .Z(n15612) );
  XNOR U16496 ( .A(n15611), .B(n15612), .Z(n15613) );
  XOR U16497 ( .A(n15614), .B(n15613), .Z(n15630) );
  NAND U16498 ( .A(n15605), .B(sreg[1654]), .Z(n15609) );
  OR U16499 ( .A(n15607), .B(n15606), .Z(n15608) );
  NAND U16500 ( .A(n15609), .B(n15608), .Z(n15629) );
  XNOR U16501 ( .A(sreg[1655]), .B(n15629), .Z(n15610) );
  XOR U16502 ( .A(n15630), .B(n15610), .Z(c[1655]) );
  NANDN U16503 ( .A(n15612), .B(n15611), .Z(n15616) );
  NAND U16504 ( .A(n15614), .B(n15613), .Z(n15615) );
  NAND U16505 ( .A(n15616), .B(n15615), .Z(n15635) );
  AND U16506 ( .A(b[2]), .B(a[634]), .Z(n15641) );
  AND U16507 ( .A(a[635]), .B(b[1]), .Z(n15639) );
  AND U16508 ( .A(a[633]), .B(b[3]), .Z(n15638) );
  XOR U16509 ( .A(n15639), .B(n15638), .Z(n15640) );
  XOR U16510 ( .A(n15641), .B(n15640), .Z(n15644) );
  NAND U16511 ( .A(b[0]), .B(a[636]), .Z(n15645) );
  XOR U16512 ( .A(n15644), .B(n15645), .Z(n15647) );
  OR U16513 ( .A(n15618), .B(n15617), .Z(n15622) );
  NANDN U16514 ( .A(n15620), .B(n15619), .Z(n15621) );
  NAND U16515 ( .A(n15622), .B(n15621), .Z(n15646) );
  XNOR U16516 ( .A(n15647), .B(n15646), .Z(n15632) );
  NANDN U16517 ( .A(n15624), .B(n15623), .Z(n15628) );
  OR U16518 ( .A(n15626), .B(n15625), .Z(n15627) );
  NAND U16519 ( .A(n15628), .B(n15627), .Z(n15633) );
  XNOR U16520 ( .A(n15632), .B(n15633), .Z(n15634) );
  XNOR U16521 ( .A(n15635), .B(n15634), .Z(n15651) );
  XOR U16522 ( .A(n15650), .B(sreg[1656]), .Z(n15631) );
  XOR U16523 ( .A(n15651), .B(n15631), .Z(c[1656]) );
  NANDN U16524 ( .A(n15633), .B(n15632), .Z(n15637) );
  NAND U16525 ( .A(n15635), .B(n15634), .Z(n15636) );
  NAND U16526 ( .A(n15637), .B(n15636), .Z(n15656) );
  AND U16527 ( .A(b[2]), .B(a[635]), .Z(n15662) );
  AND U16528 ( .A(a[636]), .B(b[1]), .Z(n15660) );
  AND U16529 ( .A(a[634]), .B(b[3]), .Z(n15659) );
  XOR U16530 ( .A(n15660), .B(n15659), .Z(n15661) );
  XOR U16531 ( .A(n15662), .B(n15661), .Z(n15665) );
  NAND U16532 ( .A(b[0]), .B(a[637]), .Z(n15666) );
  XOR U16533 ( .A(n15665), .B(n15666), .Z(n15668) );
  OR U16534 ( .A(n15639), .B(n15638), .Z(n15643) );
  NANDN U16535 ( .A(n15641), .B(n15640), .Z(n15642) );
  NAND U16536 ( .A(n15643), .B(n15642), .Z(n15667) );
  XNOR U16537 ( .A(n15668), .B(n15667), .Z(n15653) );
  NANDN U16538 ( .A(n15645), .B(n15644), .Z(n15649) );
  OR U16539 ( .A(n15647), .B(n15646), .Z(n15648) );
  NAND U16540 ( .A(n15649), .B(n15648), .Z(n15654) );
  XNOR U16541 ( .A(n15653), .B(n15654), .Z(n15655) );
  XOR U16542 ( .A(n15656), .B(n15655), .Z(n15672) );
  XOR U16543 ( .A(sreg[1657]), .B(n15671), .Z(n15652) );
  XOR U16544 ( .A(n15672), .B(n15652), .Z(c[1657]) );
  NANDN U16545 ( .A(n15654), .B(n15653), .Z(n15658) );
  NAND U16546 ( .A(n15656), .B(n15655), .Z(n15657) );
  NAND U16547 ( .A(n15658), .B(n15657), .Z(n15679) );
  AND U16548 ( .A(b[2]), .B(a[636]), .Z(n15685) );
  AND U16549 ( .A(a[637]), .B(b[1]), .Z(n15683) );
  AND U16550 ( .A(a[635]), .B(b[3]), .Z(n15682) );
  XOR U16551 ( .A(n15683), .B(n15682), .Z(n15684) );
  XOR U16552 ( .A(n15685), .B(n15684), .Z(n15688) );
  NAND U16553 ( .A(b[0]), .B(a[638]), .Z(n15689) );
  XOR U16554 ( .A(n15688), .B(n15689), .Z(n15691) );
  OR U16555 ( .A(n15660), .B(n15659), .Z(n15664) );
  NANDN U16556 ( .A(n15662), .B(n15661), .Z(n15663) );
  NAND U16557 ( .A(n15664), .B(n15663), .Z(n15690) );
  XNOR U16558 ( .A(n15691), .B(n15690), .Z(n15676) );
  NANDN U16559 ( .A(n15666), .B(n15665), .Z(n15670) );
  OR U16560 ( .A(n15668), .B(n15667), .Z(n15669) );
  NAND U16561 ( .A(n15670), .B(n15669), .Z(n15677) );
  XNOR U16562 ( .A(n15676), .B(n15677), .Z(n15678) );
  XOR U16563 ( .A(n15679), .B(n15678), .Z(n15675) );
  XNOR U16564 ( .A(sreg[1658]), .B(n15674), .Z(n15673) );
  XOR U16565 ( .A(n15675), .B(n15673), .Z(c[1658]) );
  NANDN U16566 ( .A(n15677), .B(n15676), .Z(n15681) );
  NAND U16567 ( .A(n15679), .B(n15678), .Z(n15680) );
  NAND U16568 ( .A(n15681), .B(n15680), .Z(n15697) );
  AND U16569 ( .A(b[2]), .B(a[637]), .Z(n15703) );
  AND U16570 ( .A(a[638]), .B(b[1]), .Z(n15701) );
  AND U16571 ( .A(a[636]), .B(b[3]), .Z(n15700) );
  XOR U16572 ( .A(n15701), .B(n15700), .Z(n15702) );
  XOR U16573 ( .A(n15703), .B(n15702), .Z(n15706) );
  NAND U16574 ( .A(b[0]), .B(a[639]), .Z(n15707) );
  XOR U16575 ( .A(n15706), .B(n15707), .Z(n15709) );
  OR U16576 ( .A(n15683), .B(n15682), .Z(n15687) );
  NANDN U16577 ( .A(n15685), .B(n15684), .Z(n15686) );
  NAND U16578 ( .A(n15687), .B(n15686), .Z(n15708) );
  XNOR U16579 ( .A(n15709), .B(n15708), .Z(n15694) );
  NANDN U16580 ( .A(n15689), .B(n15688), .Z(n15693) );
  OR U16581 ( .A(n15691), .B(n15690), .Z(n15692) );
  NAND U16582 ( .A(n15693), .B(n15692), .Z(n15695) );
  XNOR U16583 ( .A(n15694), .B(n15695), .Z(n15696) );
  XNOR U16584 ( .A(n15697), .B(n15696), .Z(n15712) );
  XNOR U16585 ( .A(n15712), .B(sreg[1659]), .Z(n15713) );
  XOR U16586 ( .A(n15714), .B(n15713), .Z(c[1659]) );
  NANDN U16587 ( .A(n15695), .B(n15694), .Z(n15699) );
  NAND U16588 ( .A(n15697), .B(n15696), .Z(n15698) );
  NAND U16589 ( .A(n15699), .B(n15698), .Z(n15720) );
  AND U16590 ( .A(b[2]), .B(a[638]), .Z(n15726) );
  AND U16591 ( .A(a[639]), .B(b[1]), .Z(n15724) );
  AND U16592 ( .A(a[637]), .B(b[3]), .Z(n15723) );
  XOR U16593 ( .A(n15724), .B(n15723), .Z(n15725) );
  XOR U16594 ( .A(n15726), .B(n15725), .Z(n15729) );
  NAND U16595 ( .A(b[0]), .B(a[640]), .Z(n15730) );
  XOR U16596 ( .A(n15729), .B(n15730), .Z(n15732) );
  OR U16597 ( .A(n15701), .B(n15700), .Z(n15705) );
  NANDN U16598 ( .A(n15703), .B(n15702), .Z(n15704) );
  NAND U16599 ( .A(n15705), .B(n15704), .Z(n15731) );
  XNOR U16600 ( .A(n15732), .B(n15731), .Z(n15717) );
  NANDN U16601 ( .A(n15707), .B(n15706), .Z(n15711) );
  OR U16602 ( .A(n15709), .B(n15708), .Z(n15710) );
  NAND U16603 ( .A(n15711), .B(n15710), .Z(n15718) );
  XNOR U16604 ( .A(n15717), .B(n15718), .Z(n15719) );
  XNOR U16605 ( .A(n15720), .B(n15719), .Z(n15735) );
  XOR U16606 ( .A(sreg[1660]), .B(n15735), .Z(n15736) );
  NAND U16607 ( .A(n15712), .B(sreg[1659]), .Z(n15716) );
  OR U16608 ( .A(n15714), .B(n15713), .Z(n15715) );
  NAND U16609 ( .A(n15716), .B(n15715), .Z(n15737) );
  XOR U16610 ( .A(n15736), .B(n15737), .Z(c[1660]) );
  NANDN U16611 ( .A(n15718), .B(n15717), .Z(n15722) );
  NAND U16612 ( .A(n15720), .B(n15719), .Z(n15721) );
  NAND U16613 ( .A(n15722), .B(n15721), .Z(n15758) );
  AND U16614 ( .A(b[2]), .B(a[639]), .Z(n15752) );
  AND U16615 ( .A(a[640]), .B(b[1]), .Z(n15750) );
  AND U16616 ( .A(a[638]), .B(b[3]), .Z(n15749) );
  XOR U16617 ( .A(n15750), .B(n15749), .Z(n15751) );
  XOR U16618 ( .A(n15752), .B(n15751), .Z(n15743) );
  NAND U16619 ( .A(b[0]), .B(a[641]), .Z(n15744) );
  XOR U16620 ( .A(n15743), .B(n15744), .Z(n15746) );
  OR U16621 ( .A(n15724), .B(n15723), .Z(n15728) );
  NANDN U16622 ( .A(n15726), .B(n15725), .Z(n15727) );
  NAND U16623 ( .A(n15728), .B(n15727), .Z(n15745) );
  XNOR U16624 ( .A(n15746), .B(n15745), .Z(n15755) );
  NANDN U16625 ( .A(n15730), .B(n15729), .Z(n15734) );
  OR U16626 ( .A(n15732), .B(n15731), .Z(n15733) );
  NAND U16627 ( .A(n15734), .B(n15733), .Z(n15756) );
  XNOR U16628 ( .A(n15755), .B(n15756), .Z(n15757) );
  XOR U16629 ( .A(n15758), .B(n15757), .Z(n15742) );
  OR U16630 ( .A(n15735), .B(sreg[1660]), .Z(n15739) );
  NANDN U16631 ( .A(n15737), .B(n15736), .Z(n15738) );
  AND U16632 ( .A(n15739), .B(n15738), .Z(n15741) );
  XNOR U16633 ( .A(sreg[1661]), .B(n15741), .Z(n15740) );
  XOR U16634 ( .A(n15742), .B(n15740), .Z(c[1661]) );
  NANDN U16635 ( .A(n15744), .B(n15743), .Z(n15748) );
  OR U16636 ( .A(n15746), .B(n15745), .Z(n15747) );
  NAND U16637 ( .A(n15748), .B(n15747), .Z(n15761) );
  AND U16638 ( .A(b[2]), .B(a[640]), .Z(n15770) );
  AND U16639 ( .A(a[641]), .B(b[1]), .Z(n15768) );
  AND U16640 ( .A(a[639]), .B(b[3]), .Z(n15767) );
  XOR U16641 ( .A(n15768), .B(n15767), .Z(n15769) );
  XOR U16642 ( .A(n15770), .B(n15769), .Z(n15773) );
  NAND U16643 ( .A(b[0]), .B(a[642]), .Z(n15774) );
  XNOR U16644 ( .A(n15773), .B(n15774), .Z(n15775) );
  OR U16645 ( .A(n15750), .B(n15749), .Z(n15754) );
  NANDN U16646 ( .A(n15752), .B(n15751), .Z(n15753) );
  AND U16647 ( .A(n15754), .B(n15753), .Z(n15776) );
  XNOR U16648 ( .A(n15775), .B(n15776), .Z(n15762) );
  XNOR U16649 ( .A(n15761), .B(n15762), .Z(n15763) );
  NANDN U16650 ( .A(n15756), .B(n15755), .Z(n15760) );
  NAND U16651 ( .A(n15758), .B(n15757), .Z(n15759) );
  AND U16652 ( .A(n15760), .B(n15759), .Z(n15764) );
  XOR U16653 ( .A(n15763), .B(n15764), .Z(n15779) );
  XNOR U16654 ( .A(sreg[1662]), .B(n15779), .Z(n15780) );
  XOR U16655 ( .A(n15781), .B(n15780), .Z(c[1662]) );
  NANDN U16656 ( .A(n15762), .B(n15761), .Z(n15766) );
  NAND U16657 ( .A(n15764), .B(n15763), .Z(n15765) );
  NAND U16658 ( .A(n15766), .B(n15765), .Z(n15790) );
  AND U16659 ( .A(b[2]), .B(a[641]), .Z(n15796) );
  AND U16660 ( .A(a[642]), .B(b[1]), .Z(n15794) );
  AND U16661 ( .A(a[640]), .B(b[3]), .Z(n15793) );
  XOR U16662 ( .A(n15794), .B(n15793), .Z(n15795) );
  XOR U16663 ( .A(n15796), .B(n15795), .Z(n15799) );
  NAND U16664 ( .A(b[0]), .B(a[643]), .Z(n15800) );
  XOR U16665 ( .A(n15799), .B(n15800), .Z(n15802) );
  OR U16666 ( .A(n15768), .B(n15767), .Z(n15772) );
  NANDN U16667 ( .A(n15770), .B(n15769), .Z(n15771) );
  NAND U16668 ( .A(n15772), .B(n15771), .Z(n15801) );
  XNOR U16669 ( .A(n15802), .B(n15801), .Z(n15787) );
  NANDN U16670 ( .A(n15774), .B(n15773), .Z(n15778) );
  NAND U16671 ( .A(n15776), .B(n15775), .Z(n15777) );
  NAND U16672 ( .A(n15778), .B(n15777), .Z(n15788) );
  XNOR U16673 ( .A(n15787), .B(n15788), .Z(n15789) );
  XOR U16674 ( .A(n15790), .B(n15789), .Z(n15786) );
  NAND U16675 ( .A(sreg[1662]), .B(n15779), .Z(n15783) );
  OR U16676 ( .A(n15781), .B(n15780), .Z(n15782) );
  NAND U16677 ( .A(n15783), .B(n15782), .Z(n15785) );
  XNOR U16678 ( .A(sreg[1663]), .B(n15785), .Z(n15784) );
  XNOR U16679 ( .A(n15786), .B(n15784), .Z(c[1663]) );
  NANDN U16680 ( .A(n15788), .B(n15787), .Z(n15792) );
  NANDN U16681 ( .A(n15790), .B(n15789), .Z(n15791) );
  NAND U16682 ( .A(n15792), .B(n15791), .Z(n15820) );
  AND U16683 ( .A(b[2]), .B(a[642]), .Z(n15814) );
  AND U16684 ( .A(a[643]), .B(b[1]), .Z(n15812) );
  AND U16685 ( .A(a[641]), .B(b[3]), .Z(n15811) );
  XOR U16686 ( .A(n15812), .B(n15811), .Z(n15813) );
  XOR U16687 ( .A(n15814), .B(n15813), .Z(n15805) );
  NAND U16688 ( .A(b[0]), .B(a[644]), .Z(n15806) );
  XOR U16689 ( .A(n15805), .B(n15806), .Z(n15808) );
  OR U16690 ( .A(n15794), .B(n15793), .Z(n15798) );
  NANDN U16691 ( .A(n15796), .B(n15795), .Z(n15797) );
  NAND U16692 ( .A(n15798), .B(n15797), .Z(n15807) );
  XNOR U16693 ( .A(n15808), .B(n15807), .Z(n15817) );
  NANDN U16694 ( .A(n15800), .B(n15799), .Z(n15804) );
  OR U16695 ( .A(n15802), .B(n15801), .Z(n15803) );
  NAND U16696 ( .A(n15804), .B(n15803), .Z(n15818) );
  XNOR U16697 ( .A(n15817), .B(n15818), .Z(n15819) );
  XNOR U16698 ( .A(n15820), .B(n15819), .Z(n15823) );
  XNOR U16699 ( .A(n15823), .B(sreg[1664]), .Z(n15824) );
  XOR U16700 ( .A(n15825), .B(n15824), .Z(c[1664]) );
  NANDN U16701 ( .A(n15806), .B(n15805), .Z(n15810) );
  OR U16702 ( .A(n15808), .B(n15807), .Z(n15809) );
  NAND U16703 ( .A(n15810), .B(n15809), .Z(n15828) );
  AND U16704 ( .A(b[2]), .B(a[643]), .Z(n15837) );
  AND U16705 ( .A(a[644]), .B(b[1]), .Z(n15835) );
  AND U16706 ( .A(a[642]), .B(b[3]), .Z(n15834) );
  XOR U16707 ( .A(n15835), .B(n15834), .Z(n15836) );
  XOR U16708 ( .A(n15837), .B(n15836), .Z(n15840) );
  NAND U16709 ( .A(b[0]), .B(a[645]), .Z(n15841) );
  XNOR U16710 ( .A(n15840), .B(n15841), .Z(n15842) );
  OR U16711 ( .A(n15812), .B(n15811), .Z(n15816) );
  NANDN U16712 ( .A(n15814), .B(n15813), .Z(n15815) );
  AND U16713 ( .A(n15816), .B(n15815), .Z(n15843) );
  XNOR U16714 ( .A(n15842), .B(n15843), .Z(n15829) );
  XNOR U16715 ( .A(n15828), .B(n15829), .Z(n15830) );
  NANDN U16716 ( .A(n15818), .B(n15817), .Z(n15822) );
  NAND U16717 ( .A(n15820), .B(n15819), .Z(n15821) );
  NAND U16718 ( .A(n15822), .B(n15821), .Z(n15831) );
  XNOR U16719 ( .A(n15830), .B(n15831), .Z(n15846) );
  XOR U16720 ( .A(sreg[1665]), .B(n15846), .Z(n15847) );
  NAND U16721 ( .A(n15823), .B(sreg[1664]), .Z(n15827) );
  OR U16722 ( .A(n15825), .B(n15824), .Z(n15826) );
  NAND U16723 ( .A(n15827), .B(n15826), .Z(n15848) );
  XOR U16724 ( .A(n15847), .B(n15848), .Z(c[1665]) );
  NANDN U16725 ( .A(n15829), .B(n15828), .Z(n15833) );
  NANDN U16726 ( .A(n15831), .B(n15830), .Z(n15832) );
  NAND U16727 ( .A(n15833), .B(n15832), .Z(n15857) );
  AND U16728 ( .A(b[2]), .B(a[644]), .Z(n15863) );
  AND U16729 ( .A(a[645]), .B(b[1]), .Z(n15861) );
  AND U16730 ( .A(a[643]), .B(b[3]), .Z(n15860) );
  XOR U16731 ( .A(n15861), .B(n15860), .Z(n15862) );
  XOR U16732 ( .A(n15863), .B(n15862), .Z(n15866) );
  NAND U16733 ( .A(b[0]), .B(a[646]), .Z(n15867) );
  XOR U16734 ( .A(n15866), .B(n15867), .Z(n15869) );
  OR U16735 ( .A(n15835), .B(n15834), .Z(n15839) );
  NANDN U16736 ( .A(n15837), .B(n15836), .Z(n15838) );
  NAND U16737 ( .A(n15839), .B(n15838), .Z(n15868) );
  XNOR U16738 ( .A(n15869), .B(n15868), .Z(n15854) );
  NANDN U16739 ( .A(n15841), .B(n15840), .Z(n15845) );
  NAND U16740 ( .A(n15843), .B(n15842), .Z(n15844) );
  NAND U16741 ( .A(n15845), .B(n15844), .Z(n15855) );
  XNOR U16742 ( .A(n15854), .B(n15855), .Z(n15856) );
  XOR U16743 ( .A(n15857), .B(n15856), .Z(n15853) );
  OR U16744 ( .A(n15846), .B(sreg[1665]), .Z(n15850) );
  NANDN U16745 ( .A(n15848), .B(n15847), .Z(n15849) );
  AND U16746 ( .A(n15850), .B(n15849), .Z(n15852) );
  XNOR U16747 ( .A(sreg[1666]), .B(n15852), .Z(n15851) );
  XNOR U16748 ( .A(n15853), .B(n15851), .Z(c[1666]) );
  NANDN U16749 ( .A(n15855), .B(n15854), .Z(n15859) );
  NANDN U16750 ( .A(n15857), .B(n15856), .Z(n15858) );
  NAND U16751 ( .A(n15859), .B(n15858), .Z(n15887) );
  AND U16752 ( .A(b[2]), .B(a[645]), .Z(n15881) );
  AND U16753 ( .A(a[646]), .B(b[1]), .Z(n15879) );
  AND U16754 ( .A(a[644]), .B(b[3]), .Z(n15878) );
  XOR U16755 ( .A(n15879), .B(n15878), .Z(n15880) );
  XOR U16756 ( .A(n15881), .B(n15880), .Z(n15872) );
  NAND U16757 ( .A(b[0]), .B(a[647]), .Z(n15873) );
  XOR U16758 ( .A(n15872), .B(n15873), .Z(n15875) );
  OR U16759 ( .A(n15861), .B(n15860), .Z(n15865) );
  NANDN U16760 ( .A(n15863), .B(n15862), .Z(n15864) );
  NAND U16761 ( .A(n15865), .B(n15864), .Z(n15874) );
  XNOR U16762 ( .A(n15875), .B(n15874), .Z(n15884) );
  NANDN U16763 ( .A(n15867), .B(n15866), .Z(n15871) );
  OR U16764 ( .A(n15869), .B(n15868), .Z(n15870) );
  NAND U16765 ( .A(n15871), .B(n15870), .Z(n15885) );
  XNOR U16766 ( .A(n15884), .B(n15885), .Z(n15886) );
  XNOR U16767 ( .A(n15887), .B(n15886), .Z(n15890) );
  XNOR U16768 ( .A(n15890), .B(sreg[1667]), .Z(n15891) );
  XOR U16769 ( .A(n15892), .B(n15891), .Z(c[1667]) );
  NANDN U16770 ( .A(n15873), .B(n15872), .Z(n15877) );
  OR U16771 ( .A(n15875), .B(n15874), .Z(n15876) );
  NAND U16772 ( .A(n15877), .B(n15876), .Z(n15895) );
  AND U16773 ( .A(b[2]), .B(a[646]), .Z(n15904) );
  AND U16774 ( .A(a[647]), .B(b[1]), .Z(n15902) );
  AND U16775 ( .A(a[645]), .B(b[3]), .Z(n15901) );
  XOR U16776 ( .A(n15902), .B(n15901), .Z(n15903) );
  XOR U16777 ( .A(n15904), .B(n15903), .Z(n15907) );
  NAND U16778 ( .A(b[0]), .B(a[648]), .Z(n15908) );
  XNOR U16779 ( .A(n15907), .B(n15908), .Z(n15909) );
  OR U16780 ( .A(n15879), .B(n15878), .Z(n15883) );
  NANDN U16781 ( .A(n15881), .B(n15880), .Z(n15882) );
  AND U16782 ( .A(n15883), .B(n15882), .Z(n15910) );
  XNOR U16783 ( .A(n15909), .B(n15910), .Z(n15896) );
  XNOR U16784 ( .A(n15895), .B(n15896), .Z(n15897) );
  NANDN U16785 ( .A(n15885), .B(n15884), .Z(n15889) );
  NAND U16786 ( .A(n15887), .B(n15886), .Z(n15888) );
  NAND U16787 ( .A(n15889), .B(n15888), .Z(n15898) );
  XNOR U16788 ( .A(n15897), .B(n15898), .Z(n15913) );
  XOR U16789 ( .A(sreg[1668]), .B(n15913), .Z(n15914) );
  NAND U16790 ( .A(n15890), .B(sreg[1667]), .Z(n15894) );
  OR U16791 ( .A(n15892), .B(n15891), .Z(n15893) );
  NAND U16792 ( .A(n15894), .B(n15893), .Z(n15915) );
  XOR U16793 ( .A(n15914), .B(n15915), .Z(c[1668]) );
  NANDN U16794 ( .A(n15896), .B(n15895), .Z(n15900) );
  NANDN U16795 ( .A(n15898), .B(n15897), .Z(n15899) );
  NAND U16796 ( .A(n15900), .B(n15899), .Z(n15924) );
  AND U16797 ( .A(b[2]), .B(a[647]), .Z(n15930) );
  AND U16798 ( .A(a[648]), .B(b[1]), .Z(n15928) );
  AND U16799 ( .A(a[646]), .B(b[3]), .Z(n15927) );
  XOR U16800 ( .A(n15928), .B(n15927), .Z(n15929) );
  XOR U16801 ( .A(n15930), .B(n15929), .Z(n15933) );
  NAND U16802 ( .A(b[0]), .B(a[649]), .Z(n15934) );
  XOR U16803 ( .A(n15933), .B(n15934), .Z(n15936) );
  OR U16804 ( .A(n15902), .B(n15901), .Z(n15906) );
  NANDN U16805 ( .A(n15904), .B(n15903), .Z(n15905) );
  NAND U16806 ( .A(n15906), .B(n15905), .Z(n15935) );
  XNOR U16807 ( .A(n15936), .B(n15935), .Z(n15921) );
  NANDN U16808 ( .A(n15908), .B(n15907), .Z(n15912) );
  NAND U16809 ( .A(n15910), .B(n15909), .Z(n15911) );
  NAND U16810 ( .A(n15912), .B(n15911), .Z(n15922) );
  XNOR U16811 ( .A(n15921), .B(n15922), .Z(n15923) );
  XOR U16812 ( .A(n15924), .B(n15923), .Z(n15920) );
  OR U16813 ( .A(n15913), .B(sreg[1668]), .Z(n15917) );
  NANDN U16814 ( .A(n15915), .B(n15914), .Z(n15916) );
  AND U16815 ( .A(n15917), .B(n15916), .Z(n15919) );
  XNOR U16816 ( .A(sreg[1669]), .B(n15919), .Z(n15918) );
  XNOR U16817 ( .A(n15920), .B(n15918), .Z(c[1669]) );
  NANDN U16818 ( .A(n15922), .B(n15921), .Z(n15926) );
  NANDN U16819 ( .A(n15924), .B(n15923), .Z(n15925) );
  NAND U16820 ( .A(n15926), .B(n15925), .Z(n15959) );
  AND U16821 ( .A(b[2]), .B(a[648]), .Z(n15953) );
  AND U16822 ( .A(a[649]), .B(b[1]), .Z(n15951) );
  AND U16823 ( .A(a[647]), .B(b[3]), .Z(n15950) );
  XOR U16824 ( .A(n15951), .B(n15950), .Z(n15952) );
  XOR U16825 ( .A(n15953), .B(n15952), .Z(n15944) );
  NAND U16826 ( .A(b[0]), .B(a[650]), .Z(n15945) );
  XOR U16827 ( .A(n15944), .B(n15945), .Z(n15947) );
  OR U16828 ( .A(n15928), .B(n15927), .Z(n15932) );
  NANDN U16829 ( .A(n15930), .B(n15929), .Z(n15931) );
  NAND U16830 ( .A(n15932), .B(n15931), .Z(n15946) );
  XNOR U16831 ( .A(n15947), .B(n15946), .Z(n15956) );
  NANDN U16832 ( .A(n15934), .B(n15933), .Z(n15938) );
  OR U16833 ( .A(n15936), .B(n15935), .Z(n15937) );
  NAND U16834 ( .A(n15938), .B(n15937), .Z(n15957) );
  XNOR U16835 ( .A(n15956), .B(n15957), .Z(n15958) );
  XNOR U16836 ( .A(n15959), .B(n15958), .Z(n15939) );
  XNOR U16837 ( .A(n15939), .B(sreg[1670]), .Z(n15940) );
  XOR U16838 ( .A(n15941), .B(n15940), .Z(c[1670]) );
  NAND U16839 ( .A(n15939), .B(sreg[1670]), .Z(n15943) );
  OR U16840 ( .A(n15941), .B(n15940), .Z(n15942) );
  NAND U16841 ( .A(n15943), .B(n15942), .Z(n15963) );
  NANDN U16842 ( .A(n15945), .B(n15944), .Z(n15949) );
  OR U16843 ( .A(n15947), .B(n15946), .Z(n15948) );
  NAND U16844 ( .A(n15949), .B(n15948), .Z(n15965) );
  AND U16845 ( .A(b[2]), .B(a[649]), .Z(n15974) );
  AND U16846 ( .A(a[650]), .B(b[1]), .Z(n15972) );
  AND U16847 ( .A(a[648]), .B(b[3]), .Z(n15971) );
  XOR U16848 ( .A(n15972), .B(n15971), .Z(n15973) );
  XOR U16849 ( .A(n15974), .B(n15973), .Z(n15977) );
  NAND U16850 ( .A(b[0]), .B(a[651]), .Z(n15978) );
  XNOR U16851 ( .A(n15977), .B(n15978), .Z(n15979) );
  OR U16852 ( .A(n15951), .B(n15950), .Z(n15955) );
  NANDN U16853 ( .A(n15953), .B(n15952), .Z(n15954) );
  AND U16854 ( .A(n15955), .B(n15954), .Z(n15980) );
  XNOR U16855 ( .A(n15979), .B(n15980), .Z(n15966) );
  XNOR U16856 ( .A(n15965), .B(n15966), .Z(n15967) );
  NANDN U16857 ( .A(n15957), .B(n15956), .Z(n15961) );
  NAND U16858 ( .A(n15959), .B(n15958), .Z(n15960) );
  AND U16859 ( .A(n15961), .B(n15960), .Z(n15968) );
  XNOR U16860 ( .A(n15967), .B(n15968), .Z(n15964) );
  XOR U16861 ( .A(sreg[1671]), .B(n15964), .Z(n15962) );
  XNOR U16862 ( .A(n15963), .B(n15962), .Z(c[1671]) );
  NANDN U16863 ( .A(n15966), .B(n15965), .Z(n15970) );
  NAND U16864 ( .A(n15968), .B(n15967), .Z(n15969) );
  NAND U16865 ( .A(n15970), .B(n15969), .Z(n15986) );
  AND U16866 ( .A(b[2]), .B(a[650]), .Z(n15992) );
  AND U16867 ( .A(a[651]), .B(b[1]), .Z(n15990) );
  AND U16868 ( .A(a[649]), .B(b[3]), .Z(n15989) );
  XOR U16869 ( .A(n15990), .B(n15989), .Z(n15991) );
  XOR U16870 ( .A(n15992), .B(n15991), .Z(n15995) );
  NAND U16871 ( .A(b[0]), .B(a[652]), .Z(n15996) );
  XOR U16872 ( .A(n15995), .B(n15996), .Z(n15998) );
  OR U16873 ( .A(n15972), .B(n15971), .Z(n15976) );
  NANDN U16874 ( .A(n15974), .B(n15973), .Z(n15975) );
  NAND U16875 ( .A(n15976), .B(n15975), .Z(n15997) );
  XNOR U16876 ( .A(n15998), .B(n15997), .Z(n15983) );
  NANDN U16877 ( .A(n15978), .B(n15977), .Z(n15982) );
  NAND U16878 ( .A(n15980), .B(n15979), .Z(n15981) );
  NAND U16879 ( .A(n15982), .B(n15981), .Z(n15984) );
  XNOR U16880 ( .A(n15983), .B(n15984), .Z(n15985) );
  XOR U16881 ( .A(n15986), .B(n15985), .Z(n16001) );
  XNOR U16882 ( .A(n16001), .B(sreg[1672]), .Z(n16002) );
  XOR U16883 ( .A(n16003), .B(n16002), .Z(c[1672]) );
  NANDN U16884 ( .A(n15984), .B(n15983), .Z(n15988) );
  NANDN U16885 ( .A(n15986), .B(n15985), .Z(n15987) );
  NAND U16886 ( .A(n15988), .B(n15987), .Z(n16009) );
  AND U16887 ( .A(b[2]), .B(a[651]), .Z(n16015) );
  AND U16888 ( .A(a[652]), .B(b[1]), .Z(n16013) );
  AND U16889 ( .A(a[650]), .B(b[3]), .Z(n16012) );
  XOR U16890 ( .A(n16013), .B(n16012), .Z(n16014) );
  XOR U16891 ( .A(n16015), .B(n16014), .Z(n16018) );
  NAND U16892 ( .A(b[0]), .B(a[653]), .Z(n16019) );
  XOR U16893 ( .A(n16018), .B(n16019), .Z(n16021) );
  OR U16894 ( .A(n15990), .B(n15989), .Z(n15994) );
  NANDN U16895 ( .A(n15992), .B(n15991), .Z(n15993) );
  NAND U16896 ( .A(n15994), .B(n15993), .Z(n16020) );
  XNOR U16897 ( .A(n16021), .B(n16020), .Z(n16006) );
  NANDN U16898 ( .A(n15996), .B(n15995), .Z(n16000) );
  OR U16899 ( .A(n15998), .B(n15997), .Z(n15999) );
  NAND U16900 ( .A(n16000), .B(n15999), .Z(n16007) );
  XNOR U16901 ( .A(n16006), .B(n16007), .Z(n16008) );
  XNOR U16902 ( .A(n16009), .B(n16008), .Z(n16025) );
  XNOR U16903 ( .A(n16025), .B(sreg[1673]), .Z(n16027) );
  NAND U16904 ( .A(n16001), .B(sreg[1672]), .Z(n16005) );
  OR U16905 ( .A(n16003), .B(n16002), .Z(n16004) );
  AND U16906 ( .A(n16005), .B(n16004), .Z(n16026) );
  XOR U16907 ( .A(n16027), .B(n16026), .Z(c[1673]) );
  NANDN U16908 ( .A(n16007), .B(n16006), .Z(n16011) );
  NAND U16909 ( .A(n16009), .B(n16008), .Z(n16010) );
  NAND U16910 ( .A(n16011), .B(n16010), .Z(n16035) );
  AND U16911 ( .A(b[2]), .B(a[652]), .Z(n16039) );
  AND U16912 ( .A(a[653]), .B(b[1]), .Z(n16037) );
  AND U16913 ( .A(a[651]), .B(b[3]), .Z(n16036) );
  XOR U16914 ( .A(n16037), .B(n16036), .Z(n16038) );
  XOR U16915 ( .A(n16039), .B(n16038), .Z(n16042) );
  NAND U16916 ( .A(b[0]), .B(a[654]), .Z(n16043) );
  XOR U16917 ( .A(n16042), .B(n16043), .Z(n16044) );
  OR U16918 ( .A(n16013), .B(n16012), .Z(n16017) );
  NANDN U16919 ( .A(n16015), .B(n16014), .Z(n16016) );
  AND U16920 ( .A(n16017), .B(n16016), .Z(n16045) );
  XOR U16921 ( .A(n16044), .B(n16045), .Z(n16033) );
  NANDN U16922 ( .A(n16019), .B(n16018), .Z(n16023) );
  OR U16923 ( .A(n16021), .B(n16020), .Z(n16022) );
  AND U16924 ( .A(n16023), .B(n16022), .Z(n16034) );
  XOR U16925 ( .A(n16033), .B(n16034), .Z(n16024) );
  XOR U16926 ( .A(n16035), .B(n16024), .Z(n16032) );
  NAND U16927 ( .A(n16025), .B(sreg[1673]), .Z(n16029) );
  OR U16928 ( .A(n16027), .B(n16026), .Z(n16028) );
  AND U16929 ( .A(n16029), .B(n16028), .Z(n16031) );
  XNOR U16930 ( .A(n16031), .B(sreg[1674]), .Z(n16030) );
  XNOR U16931 ( .A(n16032), .B(n16030), .Z(c[1674]) );
  AND U16932 ( .A(b[2]), .B(a[653]), .Z(n16055) );
  AND U16933 ( .A(a[654]), .B(b[1]), .Z(n16053) );
  AND U16934 ( .A(a[652]), .B(b[3]), .Z(n16052) );
  XOR U16935 ( .A(n16053), .B(n16052), .Z(n16054) );
  XOR U16936 ( .A(n16055), .B(n16054), .Z(n16046) );
  NAND U16937 ( .A(b[0]), .B(a[655]), .Z(n16047) );
  XOR U16938 ( .A(n16046), .B(n16047), .Z(n16049) );
  OR U16939 ( .A(n16037), .B(n16036), .Z(n16041) );
  NANDN U16940 ( .A(n16039), .B(n16038), .Z(n16040) );
  NAND U16941 ( .A(n16041), .B(n16040), .Z(n16048) );
  XNOR U16942 ( .A(n16049), .B(n16048), .Z(n16058) );
  XNOR U16943 ( .A(n16058), .B(n16059), .Z(n16061) );
  XOR U16944 ( .A(n16060), .B(n16061), .Z(n16064) );
  XOR U16945 ( .A(n16064), .B(sreg[1675]), .Z(n16066) );
  XNOR U16946 ( .A(n16065), .B(n16066), .Z(c[1675]) );
  NANDN U16947 ( .A(n16047), .B(n16046), .Z(n16051) );
  OR U16948 ( .A(n16049), .B(n16048), .Z(n16050) );
  NAND U16949 ( .A(n16051), .B(n16050), .Z(n16070) );
  AND U16950 ( .A(b[2]), .B(a[654]), .Z(n16085) );
  AND U16951 ( .A(a[655]), .B(b[1]), .Z(n16083) );
  AND U16952 ( .A(a[653]), .B(b[3]), .Z(n16082) );
  XOR U16953 ( .A(n16083), .B(n16082), .Z(n16084) );
  XOR U16954 ( .A(n16085), .B(n16084), .Z(n16076) );
  NAND U16955 ( .A(b[0]), .B(a[656]), .Z(n16077) );
  XNOR U16956 ( .A(n16076), .B(n16077), .Z(n16078) );
  OR U16957 ( .A(n16053), .B(n16052), .Z(n16057) );
  NANDN U16958 ( .A(n16055), .B(n16054), .Z(n16056) );
  AND U16959 ( .A(n16057), .B(n16056), .Z(n16079) );
  XNOR U16960 ( .A(n16078), .B(n16079), .Z(n16071) );
  XNOR U16961 ( .A(n16070), .B(n16071), .Z(n16072) );
  NANDN U16962 ( .A(n16059), .B(n16058), .Z(n16063) );
  NAND U16963 ( .A(n16061), .B(n16060), .Z(n16062) );
  NAND U16964 ( .A(n16063), .B(n16062), .Z(n16073) );
  XOR U16965 ( .A(n16072), .B(n16073), .Z(n16090) );
  NANDN U16966 ( .A(n16064), .B(sreg[1675]), .Z(n16068) );
  NANDN U16967 ( .A(n16066), .B(n16065), .Z(n16067) );
  AND U16968 ( .A(n16068), .B(n16067), .Z(n16089) );
  XNOR U16969 ( .A(n16089), .B(sreg[1676]), .Z(n16069) );
  XNOR U16970 ( .A(n16090), .B(n16069), .Z(c[1676]) );
  NANDN U16971 ( .A(n16071), .B(n16070), .Z(n16075) );
  NANDN U16972 ( .A(n16073), .B(n16072), .Z(n16074) );
  NAND U16973 ( .A(n16075), .B(n16074), .Z(n16094) );
  NANDN U16974 ( .A(n16077), .B(n16076), .Z(n16081) );
  NAND U16975 ( .A(n16079), .B(n16078), .Z(n16080) );
  AND U16976 ( .A(n16081), .B(n16080), .Z(n16093) );
  AND U16977 ( .A(b[2]), .B(a[655]), .Z(n16098) );
  AND U16978 ( .A(a[656]), .B(b[1]), .Z(n16096) );
  AND U16979 ( .A(a[654]), .B(b[3]), .Z(n16095) );
  XOR U16980 ( .A(n16096), .B(n16095), .Z(n16097) );
  XOR U16981 ( .A(n16098), .B(n16097), .Z(n16101) );
  NAND U16982 ( .A(b[0]), .B(a[657]), .Z(n16102) );
  XOR U16983 ( .A(n16101), .B(n16102), .Z(n16104) );
  OR U16984 ( .A(n16083), .B(n16082), .Z(n16087) );
  NANDN U16985 ( .A(n16085), .B(n16084), .Z(n16086) );
  NAND U16986 ( .A(n16087), .B(n16086), .Z(n16103) );
  XOR U16987 ( .A(n16104), .B(n16103), .Z(n16092) );
  XNOR U16988 ( .A(n16093), .B(n16092), .Z(n16088) );
  XOR U16989 ( .A(n16094), .B(n16088), .Z(n16108) );
  XOR U16990 ( .A(sreg[1677]), .B(n16107), .Z(n16091) );
  XNOR U16991 ( .A(n16108), .B(n16091), .Z(c[1677]) );
  AND U16992 ( .A(b[2]), .B(a[656]), .Z(n16121) );
  AND U16993 ( .A(a[657]), .B(b[1]), .Z(n16119) );
  AND U16994 ( .A(a[655]), .B(b[3]), .Z(n16118) );
  XOR U16995 ( .A(n16119), .B(n16118), .Z(n16120) );
  XOR U16996 ( .A(n16121), .B(n16120), .Z(n16124) );
  NAND U16997 ( .A(b[0]), .B(a[658]), .Z(n16125) );
  XOR U16998 ( .A(n16124), .B(n16125), .Z(n16127) );
  OR U16999 ( .A(n16096), .B(n16095), .Z(n16100) );
  NANDN U17000 ( .A(n16098), .B(n16097), .Z(n16099) );
  NAND U17001 ( .A(n16100), .B(n16099), .Z(n16126) );
  XNOR U17002 ( .A(n16127), .B(n16126), .Z(n16112) );
  NANDN U17003 ( .A(n16102), .B(n16101), .Z(n16106) );
  OR U17004 ( .A(n16104), .B(n16103), .Z(n16105) );
  NAND U17005 ( .A(n16106), .B(n16105), .Z(n16113) );
  XNOR U17006 ( .A(n16112), .B(n16113), .Z(n16114) );
  XNOR U17007 ( .A(n16115), .B(n16114), .Z(n16111) );
  XOR U17008 ( .A(n16110), .B(sreg[1678]), .Z(n16109) );
  XNOR U17009 ( .A(n16111), .B(n16109), .Z(c[1678]) );
  NANDN U17010 ( .A(n16113), .B(n16112), .Z(n16117) );
  NANDN U17011 ( .A(n16115), .B(n16114), .Z(n16116) );
  NAND U17012 ( .A(n16117), .B(n16116), .Z(n16133) );
  AND U17013 ( .A(b[2]), .B(a[657]), .Z(n16139) );
  AND U17014 ( .A(a[658]), .B(b[1]), .Z(n16137) );
  AND U17015 ( .A(a[656]), .B(b[3]), .Z(n16136) );
  XOR U17016 ( .A(n16137), .B(n16136), .Z(n16138) );
  XOR U17017 ( .A(n16139), .B(n16138), .Z(n16142) );
  NAND U17018 ( .A(b[0]), .B(a[659]), .Z(n16143) );
  XOR U17019 ( .A(n16142), .B(n16143), .Z(n16145) );
  OR U17020 ( .A(n16119), .B(n16118), .Z(n16123) );
  NANDN U17021 ( .A(n16121), .B(n16120), .Z(n16122) );
  NAND U17022 ( .A(n16123), .B(n16122), .Z(n16144) );
  XNOR U17023 ( .A(n16145), .B(n16144), .Z(n16130) );
  NANDN U17024 ( .A(n16125), .B(n16124), .Z(n16129) );
  OR U17025 ( .A(n16127), .B(n16126), .Z(n16128) );
  NAND U17026 ( .A(n16129), .B(n16128), .Z(n16131) );
  XNOR U17027 ( .A(n16130), .B(n16131), .Z(n16132) );
  XNOR U17028 ( .A(n16133), .B(n16132), .Z(n16149) );
  XOR U17029 ( .A(sreg[1679]), .B(n16149), .Z(n16150) );
  XOR U17030 ( .A(n16151), .B(n16150), .Z(c[1679]) );
  NANDN U17031 ( .A(n16131), .B(n16130), .Z(n16135) );
  NAND U17032 ( .A(n16133), .B(n16132), .Z(n16134) );
  AND U17033 ( .A(n16135), .B(n16134), .Z(n16159) );
  AND U17034 ( .A(b[2]), .B(a[658]), .Z(n16167) );
  AND U17035 ( .A(a[659]), .B(b[1]), .Z(n16165) );
  AND U17036 ( .A(a[657]), .B(b[3]), .Z(n16164) );
  XOR U17037 ( .A(n16165), .B(n16164), .Z(n16166) );
  XOR U17038 ( .A(n16167), .B(n16166), .Z(n16160) );
  NAND U17039 ( .A(b[0]), .B(a[660]), .Z(n16161) );
  XOR U17040 ( .A(n16160), .B(n16161), .Z(n16162) );
  OR U17041 ( .A(n16137), .B(n16136), .Z(n16141) );
  NANDN U17042 ( .A(n16139), .B(n16138), .Z(n16140) );
  AND U17043 ( .A(n16141), .B(n16140), .Z(n16163) );
  XOR U17044 ( .A(n16162), .B(n16163), .Z(n16157) );
  NANDN U17045 ( .A(n16143), .B(n16142), .Z(n16147) );
  OR U17046 ( .A(n16145), .B(n16144), .Z(n16146) );
  AND U17047 ( .A(n16147), .B(n16146), .Z(n16158) );
  XOR U17048 ( .A(n16157), .B(n16158), .Z(n16148) );
  XNOR U17049 ( .A(n16159), .B(n16148), .Z(n16156) );
  OR U17050 ( .A(n16149), .B(sreg[1679]), .Z(n16153) );
  NANDN U17051 ( .A(n16151), .B(n16150), .Z(n16152) );
  AND U17052 ( .A(n16153), .B(n16152), .Z(n16155) );
  XNOR U17053 ( .A(sreg[1680]), .B(n16155), .Z(n16154) );
  XOR U17054 ( .A(n16156), .B(n16154), .Z(c[1680]) );
  AND U17055 ( .A(b[2]), .B(a[659]), .Z(n16173) );
  AND U17056 ( .A(a[660]), .B(b[1]), .Z(n16171) );
  AND U17057 ( .A(a[658]), .B(b[3]), .Z(n16170) );
  XOR U17058 ( .A(n16171), .B(n16170), .Z(n16172) );
  XOR U17059 ( .A(n16173), .B(n16172), .Z(n16176) );
  NAND U17060 ( .A(b[0]), .B(a[661]), .Z(n16177) );
  XNOR U17061 ( .A(n16176), .B(n16177), .Z(n16178) );
  OR U17062 ( .A(n16165), .B(n16164), .Z(n16169) );
  NANDN U17063 ( .A(n16167), .B(n16166), .Z(n16168) );
  AND U17064 ( .A(n16169), .B(n16168), .Z(n16179) );
  XNOR U17065 ( .A(n16178), .B(n16179), .Z(n16183) );
  XNOR U17066 ( .A(n16182), .B(n16183), .Z(n16184) );
  XNOR U17067 ( .A(n16185), .B(n16184), .Z(n16188) );
  XNOR U17068 ( .A(sreg[1681]), .B(n16188), .Z(n16189) );
  XOR U17069 ( .A(n16190), .B(n16189), .Z(c[1681]) );
  AND U17070 ( .A(b[2]), .B(a[660]), .Z(n16205) );
  AND U17071 ( .A(a[661]), .B(b[1]), .Z(n16203) );
  AND U17072 ( .A(a[659]), .B(b[3]), .Z(n16202) );
  XOR U17073 ( .A(n16203), .B(n16202), .Z(n16204) );
  XOR U17074 ( .A(n16205), .B(n16204), .Z(n16208) );
  NAND U17075 ( .A(b[0]), .B(a[662]), .Z(n16209) );
  XOR U17076 ( .A(n16208), .B(n16209), .Z(n16211) );
  OR U17077 ( .A(n16171), .B(n16170), .Z(n16175) );
  NANDN U17078 ( .A(n16173), .B(n16172), .Z(n16174) );
  NAND U17079 ( .A(n16175), .B(n16174), .Z(n16210) );
  XNOR U17080 ( .A(n16211), .B(n16210), .Z(n16196) );
  NANDN U17081 ( .A(n16177), .B(n16176), .Z(n16181) );
  NAND U17082 ( .A(n16179), .B(n16178), .Z(n16180) );
  NAND U17083 ( .A(n16181), .B(n16180), .Z(n16197) );
  XNOR U17084 ( .A(n16196), .B(n16197), .Z(n16198) );
  NANDN U17085 ( .A(n16183), .B(n16182), .Z(n16187) );
  NANDN U17086 ( .A(n16185), .B(n16184), .Z(n16186) );
  NAND U17087 ( .A(n16187), .B(n16186), .Z(n16199) );
  XOR U17088 ( .A(n16198), .B(n16199), .Z(n16195) );
  NAND U17089 ( .A(sreg[1681]), .B(n16188), .Z(n16192) );
  OR U17090 ( .A(n16190), .B(n16189), .Z(n16191) );
  NAND U17091 ( .A(n16192), .B(n16191), .Z(n16194) );
  XNOR U17092 ( .A(sreg[1682]), .B(n16194), .Z(n16193) );
  XNOR U17093 ( .A(n16195), .B(n16193), .Z(c[1682]) );
  NANDN U17094 ( .A(n16197), .B(n16196), .Z(n16201) );
  NANDN U17095 ( .A(n16199), .B(n16198), .Z(n16200) );
  NAND U17096 ( .A(n16201), .B(n16200), .Z(n16234) );
  AND U17097 ( .A(b[2]), .B(a[661]), .Z(n16228) );
  AND U17098 ( .A(a[662]), .B(b[1]), .Z(n16226) );
  AND U17099 ( .A(a[660]), .B(b[3]), .Z(n16225) );
  XOR U17100 ( .A(n16226), .B(n16225), .Z(n16227) );
  XOR U17101 ( .A(n16228), .B(n16227), .Z(n16219) );
  NAND U17102 ( .A(b[0]), .B(a[663]), .Z(n16220) );
  XOR U17103 ( .A(n16219), .B(n16220), .Z(n16222) );
  OR U17104 ( .A(n16203), .B(n16202), .Z(n16207) );
  NANDN U17105 ( .A(n16205), .B(n16204), .Z(n16206) );
  NAND U17106 ( .A(n16207), .B(n16206), .Z(n16221) );
  XNOR U17107 ( .A(n16222), .B(n16221), .Z(n16231) );
  NANDN U17108 ( .A(n16209), .B(n16208), .Z(n16213) );
  OR U17109 ( .A(n16211), .B(n16210), .Z(n16212) );
  NAND U17110 ( .A(n16213), .B(n16212), .Z(n16232) );
  XNOR U17111 ( .A(n16231), .B(n16232), .Z(n16233) );
  XNOR U17112 ( .A(n16234), .B(n16233), .Z(n16214) );
  XNOR U17113 ( .A(n16214), .B(sreg[1683]), .Z(n16215) );
  XOR U17114 ( .A(n16216), .B(n16215), .Z(c[1683]) );
  NAND U17115 ( .A(n16214), .B(sreg[1683]), .Z(n16218) );
  OR U17116 ( .A(n16216), .B(n16215), .Z(n16217) );
  NAND U17117 ( .A(n16218), .B(n16217), .Z(n16256) );
  NANDN U17118 ( .A(n16220), .B(n16219), .Z(n16224) );
  OR U17119 ( .A(n16222), .B(n16221), .Z(n16223) );
  NAND U17120 ( .A(n16224), .B(n16223), .Z(n16238) );
  AND U17121 ( .A(b[2]), .B(a[662]), .Z(n16247) );
  AND U17122 ( .A(a[663]), .B(b[1]), .Z(n16245) );
  AND U17123 ( .A(a[661]), .B(b[3]), .Z(n16244) );
  XOR U17124 ( .A(n16245), .B(n16244), .Z(n16246) );
  XOR U17125 ( .A(n16247), .B(n16246), .Z(n16250) );
  NAND U17126 ( .A(b[0]), .B(a[664]), .Z(n16251) );
  XNOR U17127 ( .A(n16250), .B(n16251), .Z(n16252) );
  OR U17128 ( .A(n16226), .B(n16225), .Z(n16230) );
  NANDN U17129 ( .A(n16228), .B(n16227), .Z(n16229) );
  AND U17130 ( .A(n16230), .B(n16229), .Z(n16253) );
  XNOR U17131 ( .A(n16252), .B(n16253), .Z(n16239) );
  XNOR U17132 ( .A(n16238), .B(n16239), .Z(n16240) );
  NANDN U17133 ( .A(n16232), .B(n16231), .Z(n16236) );
  NAND U17134 ( .A(n16234), .B(n16233), .Z(n16235) );
  AND U17135 ( .A(n16236), .B(n16235), .Z(n16241) );
  XNOR U17136 ( .A(n16240), .B(n16241), .Z(n16257) );
  XOR U17137 ( .A(sreg[1684]), .B(n16257), .Z(n16237) );
  XNOR U17138 ( .A(n16256), .B(n16237), .Z(c[1684]) );
  NANDN U17139 ( .A(n16239), .B(n16238), .Z(n16243) );
  NAND U17140 ( .A(n16241), .B(n16240), .Z(n16242) );
  NAND U17141 ( .A(n16243), .B(n16242), .Z(n16262) );
  AND U17142 ( .A(b[2]), .B(a[663]), .Z(n16268) );
  AND U17143 ( .A(a[664]), .B(b[1]), .Z(n16266) );
  AND U17144 ( .A(a[662]), .B(b[3]), .Z(n16265) );
  XOR U17145 ( .A(n16266), .B(n16265), .Z(n16267) );
  XOR U17146 ( .A(n16268), .B(n16267), .Z(n16271) );
  NAND U17147 ( .A(b[0]), .B(a[665]), .Z(n16272) );
  XOR U17148 ( .A(n16271), .B(n16272), .Z(n16274) );
  OR U17149 ( .A(n16245), .B(n16244), .Z(n16249) );
  NANDN U17150 ( .A(n16247), .B(n16246), .Z(n16248) );
  NAND U17151 ( .A(n16249), .B(n16248), .Z(n16273) );
  XNOR U17152 ( .A(n16274), .B(n16273), .Z(n16259) );
  NANDN U17153 ( .A(n16251), .B(n16250), .Z(n16255) );
  NAND U17154 ( .A(n16253), .B(n16252), .Z(n16254) );
  NAND U17155 ( .A(n16255), .B(n16254), .Z(n16260) );
  XNOR U17156 ( .A(n16259), .B(n16260), .Z(n16261) );
  XOR U17157 ( .A(n16262), .B(n16261), .Z(n16278) );
  XNOR U17158 ( .A(sreg[1685]), .B(n16277), .Z(n16258) );
  XNOR U17159 ( .A(n16278), .B(n16258), .Z(c[1685]) );
  NANDN U17160 ( .A(n16260), .B(n16259), .Z(n16264) );
  NANDN U17161 ( .A(n16262), .B(n16261), .Z(n16263) );
  NAND U17162 ( .A(n16264), .B(n16263), .Z(n16283) );
  AND U17163 ( .A(b[2]), .B(a[664]), .Z(n16289) );
  AND U17164 ( .A(a[665]), .B(b[1]), .Z(n16287) );
  AND U17165 ( .A(a[663]), .B(b[3]), .Z(n16286) );
  XOR U17166 ( .A(n16287), .B(n16286), .Z(n16288) );
  XOR U17167 ( .A(n16289), .B(n16288), .Z(n16292) );
  NAND U17168 ( .A(b[0]), .B(a[666]), .Z(n16293) );
  XOR U17169 ( .A(n16292), .B(n16293), .Z(n16295) );
  OR U17170 ( .A(n16266), .B(n16265), .Z(n16270) );
  NANDN U17171 ( .A(n16268), .B(n16267), .Z(n16269) );
  NAND U17172 ( .A(n16270), .B(n16269), .Z(n16294) );
  XNOR U17173 ( .A(n16295), .B(n16294), .Z(n16280) );
  NANDN U17174 ( .A(n16272), .B(n16271), .Z(n16276) );
  OR U17175 ( .A(n16274), .B(n16273), .Z(n16275) );
  NAND U17176 ( .A(n16276), .B(n16275), .Z(n16281) );
  XNOR U17177 ( .A(n16280), .B(n16281), .Z(n16282) );
  XNOR U17178 ( .A(n16283), .B(n16282), .Z(n16299) );
  XOR U17179 ( .A(n16298), .B(sreg[1686]), .Z(n16279) );
  XOR U17180 ( .A(n16299), .B(n16279), .Z(c[1686]) );
  NANDN U17181 ( .A(n16281), .B(n16280), .Z(n16285) );
  NAND U17182 ( .A(n16283), .B(n16282), .Z(n16284) );
  NAND U17183 ( .A(n16285), .B(n16284), .Z(n16306) );
  AND U17184 ( .A(b[2]), .B(a[665]), .Z(n16312) );
  AND U17185 ( .A(a[666]), .B(b[1]), .Z(n16310) );
  AND U17186 ( .A(a[664]), .B(b[3]), .Z(n16309) );
  XOR U17187 ( .A(n16310), .B(n16309), .Z(n16311) );
  XOR U17188 ( .A(n16312), .B(n16311), .Z(n16315) );
  NAND U17189 ( .A(b[0]), .B(a[667]), .Z(n16316) );
  XOR U17190 ( .A(n16315), .B(n16316), .Z(n16318) );
  OR U17191 ( .A(n16287), .B(n16286), .Z(n16291) );
  NANDN U17192 ( .A(n16289), .B(n16288), .Z(n16290) );
  NAND U17193 ( .A(n16291), .B(n16290), .Z(n16317) );
  XNOR U17194 ( .A(n16318), .B(n16317), .Z(n16303) );
  NANDN U17195 ( .A(n16293), .B(n16292), .Z(n16297) );
  OR U17196 ( .A(n16295), .B(n16294), .Z(n16296) );
  NAND U17197 ( .A(n16297), .B(n16296), .Z(n16304) );
  XNOR U17198 ( .A(n16303), .B(n16304), .Z(n16305) );
  XNOR U17199 ( .A(n16306), .B(n16305), .Z(n16302) );
  XOR U17200 ( .A(n16301), .B(sreg[1687]), .Z(n16300) );
  XOR U17201 ( .A(n16302), .B(n16300), .Z(c[1687]) );
  NANDN U17202 ( .A(n16304), .B(n16303), .Z(n16308) );
  NAND U17203 ( .A(n16306), .B(n16305), .Z(n16307) );
  NAND U17204 ( .A(n16308), .B(n16307), .Z(n16324) );
  AND U17205 ( .A(b[2]), .B(a[666]), .Z(n16330) );
  AND U17206 ( .A(a[667]), .B(b[1]), .Z(n16328) );
  AND U17207 ( .A(a[665]), .B(b[3]), .Z(n16327) );
  XOR U17208 ( .A(n16328), .B(n16327), .Z(n16329) );
  XOR U17209 ( .A(n16330), .B(n16329), .Z(n16333) );
  NAND U17210 ( .A(b[0]), .B(a[668]), .Z(n16334) );
  XOR U17211 ( .A(n16333), .B(n16334), .Z(n16336) );
  OR U17212 ( .A(n16310), .B(n16309), .Z(n16314) );
  NANDN U17213 ( .A(n16312), .B(n16311), .Z(n16313) );
  NAND U17214 ( .A(n16314), .B(n16313), .Z(n16335) );
  XNOR U17215 ( .A(n16336), .B(n16335), .Z(n16321) );
  NANDN U17216 ( .A(n16316), .B(n16315), .Z(n16320) );
  OR U17217 ( .A(n16318), .B(n16317), .Z(n16319) );
  NAND U17218 ( .A(n16320), .B(n16319), .Z(n16322) );
  XNOR U17219 ( .A(n16321), .B(n16322), .Z(n16323) );
  XNOR U17220 ( .A(n16324), .B(n16323), .Z(n16339) );
  XNOR U17221 ( .A(n16339), .B(sreg[1688]), .Z(n16341) );
  XNOR U17222 ( .A(n16340), .B(n16341), .Z(c[1688]) );
  NANDN U17223 ( .A(n16322), .B(n16321), .Z(n16326) );
  NAND U17224 ( .A(n16324), .B(n16323), .Z(n16325) );
  NAND U17225 ( .A(n16326), .B(n16325), .Z(n16352) );
  AND U17226 ( .A(b[2]), .B(a[667]), .Z(n16358) );
  AND U17227 ( .A(a[668]), .B(b[1]), .Z(n16356) );
  AND U17228 ( .A(a[666]), .B(b[3]), .Z(n16355) );
  XOR U17229 ( .A(n16356), .B(n16355), .Z(n16357) );
  XOR U17230 ( .A(n16358), .B(n16357), .Z(n16361) );
  NAND U17231 ( .A(b[0]), .B(a[669]), .Z(n16362) );
  XOR U17232 ( .A(n16361), .B(n16362), .Z(n16364) );
  OR U17233 ( .A(n16328), .B(n16327), .Z(n16332) );
  NANDN U17234 ( .A(n16330), .B(n16329), .Z(n16331) );
  NAND U17235 ( .A(n16332), .B(n16331), .Z(n16363) );
  XNOR U17236 ( .A(n16364), .B(n16363), .Z(n16349) );
  NANDN U17237 ( .A(n16334), .B(n16333), .Z(n16338) );
  OR U17238 ( .A(n16336), .B(n16335), .Z(n16337) );
  NAND U17239 ( .A(n16338), .B(n16337), .Z(n16350) );
  XNOR U17240 ( .A(n16349), .B(n16350), .Z(n16351) );
  XNOR U17241 ( .A(n16352), .B(n16351), .Z(n16344) );
  XNOR U17242 ( .A(n16344), .B(sreg[1689]), .Z(n16346) );
  NAND U17243 ( .A(n16339), .B(sreg[1688]), .Z(n16343) );
  NANDN U17244 ( .A(n16341), .B(n16340), .Z(n16342) );
  AND U17245 ( .A(n16343), .B(n16342), .Z(n16345) );
  XOR U17246 ( .A(n16346), .B(n16345), .Z(c[1689]) );
  NAND U17247 ( .A(n16344), .B(sreg[1689]), .Z(n16348) );
  OR U17248 ( .A(n16346), .B(n16345), .Z(n16347) );
  AND U17249 ( .A(n16348), .B(n16347), .Z(n16387) );
  NANDN U17250 ( .A(n16350), .B(n16349), .Z(n16354) );
  NAND U17251 ( .A(n16352), .B(n16351), .Z(n16353) );
  NAND U17252 ( .A(n16354), .B(n16353), .Z(n16371) );
  AND U17253 ( .A(b[2]), .B(a[668]), .Z(n16377) );
  AND U17254 ( .A(a[669]), .B(b[1]), .Z(n16375) );
  AND U17255 ( .A(a[667]), .B(b[3]), .Z(n16374) );
  XOR U17256 ( .A(n16375), .B(n16374), .Z(n16376) );
  XOR U17257 ( .A(n16377), .B(n16376), .Z(n16380) );
  NAND U17258 ( .A(b[0]), .B(a[670]), .Z(n16381) );
  XOR U17259 ( .A(n16380), .B(n16381), .Z(n16383) );
  OR U17260 ( .A(n16356), .B(n16355), .Z(n16360) );
  NANDN U17261 ( .A(n16358), .B(n16357), .Z(n16359) );
  NAND U17262 ( .A(n16360), .B(n16359), .Z(n16382) );
  XNOR U17263 ( .A(n16383), .B(n16382), .Z(n16368) );
  NANDN U17264 ( .A(n16362), .B(n16361), .Z(n16366) );
  OR U17265 ( .A(n16364), .B(n16363), .Z(n16365) );
  NAND U17266 ( .A(n16366), .B(n16365), .Z(n16369) );
  XNOR U17267 ( .A(n16368), .B(n16369), .Z(n16370) );
  XNOR U17268 ( .A(n16371), .B(n16370), .Z(n16386) );
  XNOR U17269 ( .A(sreg[1690]), .B(n16386), .Z(n16367) );
  XOR U17270 ( .A(n16387), .B(n16367), .Z(c[1690]) );
  NANDN U17271 ( .A(n16369), .B(n16368), .Z(n16373) );
  NAND U17272 ( .A(n16371), .B(n16370), .Z(n16372) );
  NAND U17273 ( .A(n16373), .B(n16372), .Z(n16394) );
  AND U17274 ( .A(b[2]), .B(a[669]), .Z(n16400) );
  AND U17275 ( .A(a[670]), .B(b[1]), .Z(n16398) );
  AND U17276 ( .A(a[668]), .B(b[3]), .Z(n16397) );
  XOR U17277 ( .A(n16398), .B(n16397), .Z(n16399) );
  XOR U17278 ( .A(n16400), .B(n16399), .Z(n16403) );
  NAND U17279 ( .A(b[0]), .B(a[671]), .Z(n16404) );
  XOR U17280 ( .A(n16403), .B(n16404), .Z(n16406) );
  OR U17281 ( .A(n16375), .B(n16374), .Z(n16379) );
  NANDN U17282 ( .A(n16377), .B(n16376), .Z(n16378) );
  NAND U17283 ( .A(n16379), .B(n16378), .Z(n16405) );
  XNOR U17284 ( .A(n16406), .B(n16405), .Z(n16391) );
  NANDN U17285 ( .A(n16381), .B(n16380), .Z(n16385) );
  OR U17286 ( .A(n16383), .B(n16382), .Z(n16384) );
  NAND U17287 ( .A(n16385), .B(n16384), .Z(n16392) );
  XNOR U17288 ( .A(n16391), .B(n16392), .Z(n16393) );
  XOR U17289 ( .A(n16394), .B(n16393), .Z(n16390) );
  XNOR U17290 ( .A(sreg[1691]), .B(n16389), .Z(n16388) );
  XOR U17291 ( .A(n16390), .B(n16388), .Z(c[1691]) );
  NANDN U17292 ( .A(n16392), .B(n16391), .Z(n16396) );
  NAND U17293 ( .A(n16394), .B(n16393), .Z(n16395) );
  NAND U17294 ( .A(n16396), .B(n16395), .Z(n16412) );
  AND U17295 ( .A(b[2]), .B(a[670]), .Z(n16418) );
  AND U17296 ( .A(a[671]), .B(b[1]), .Z(n16416) );
  AND U17297 ( .A(a[669]), .B(b[3]), .Z(n16415) );
  XOR U17298 ( .A(n16416), .B(n16415), .Z(n16417) );
  XOR U17299 ( .A(n16418), .B(n16417), .Z(n16421) );
  NAND U17300 ( .A(b[0]), .B(a[672]), .Z(n16422) );
  XOR U17301 ( .A(n16421), .B(n16422), .Z(n16424) );
  OR U17302 ( .A(n16398), .B(n16397), .Z(n16402) );
  NANDN U17303 ( .A(n16400), .B(n16399), .Z(n16401) );
  NAND U17304 ( .A(n16402), .B(n16401), .Z(n16423) );
  XNOR U17305 ( .A(n16424), .B(n16423), .Z(n16409) );
  NANDN U17306 ( .A(n16404), .B(n16403), .Z(n16408) );
  OR U17307 ( .A(n16406), .B(n16405), .Z(n16407) );
  NAND U17308 ( .A(n16408), .B(n16407), .Z(n16410) );
  XNOR U17309 ( .A(n16409), .B(n16410), .Z(n16411) );
  XNOR U17310 ( .A(n16412), .B(n16411), .Z(n16427) );
  XNOR U17311 ( .A(n16427), .B(sreg[1692]), .Z(n16428) );
  XOR U17312 ( .A(n16429), .B(n16428), .Z(c[1692]) );
  NANDN U17313 ( .A(n16410), .B(n16409), .Z(n16414) );
  NAND U17314 ( .A(n16412), .B(n16411), .Z(n16413) );
  NAND U17315 ( .A(n16414), .B(n16413), .Z(n16440) );
  AND U17316 ( .A(b[2]), .B(a[671]), .Z(n16446) );
  AND U17317 ( .A(a[672]), .B(b[1]), .Z(n16444) );
  AND U17318 ( .A(a[670]), .B(b[3]), .Z(n16443) );
  XOR U17319 ( .A(n16444), .B(n16443), .Z(n16445) );
  XOR U17320 ( .A(n16446), .B(n16445), .Z(n16449) );
  NAND U17321 ( .A(b[0]), .B(a[673]), .Z(n16450) );
  XOR U17322 ( .A(n16449), .B(n16450), .Z(n16452) );
  OR U17323 ( .A(n16416), .B(n16415), .Z(n16420) );
  NANDN U17324 ( .A(n16418), .B(n16417), .Z(n16419) );
  NAND U17325 ( .A(n16420), .B(n16419), .Z(n16451) );
  XNOR U17326 ( .A(n16452), .B(n16451), .Z(n16437) );
  NANDN U17327 ( .A(n16422), .B(n16421), .Z(n16426) );
  OR U17328 ( .A(n16424), .B(n16423), .Z(n16425) );
  NAND U17329 ( .A(n16426), .B(n16425), .Z(n16438) );
  XNOR U17330 ( .A(n16437), .B(n16438), .Z(n16439) );
  XNOR U17331 ( .A(n16440), .B(n16439), .Z(n16432) );
  XOR U17332 ( .A(sreg[1693]), .B(n16432), .Z(n16433) );
  NAND U17333 ( .A(n16427), .B(sreg[1692]), .Z(n16431) );
  OR U17334 ( .A(n16429), .B(n16428), .Z(n16430) );
  NAND U17335 ( .A(n16431), .B(n16430), .Z(n16434) );
  XOR U17336 ( .A(n16433), .B(n16434), .Z(c[1693]) );
  OR U17337 ( .A(n16432), .B(sreg[1693]), .Z(n16436) );
  NANDN U17338 ( .A(n16434), .B(n16433), .Z(n16435) );
  AND U17339 ( .A(n16436), .B(n16435), .Z(n16456) );
  NANDN U17340 ( .A(n16438), .B(n16437), .Z(n16442) );
  NAND U17341 ( .A(n16440), .B(n16439), .Z(n16441) );
  NAND U17342 ( .A(n16442), .B(n16441), .Z(n16461) );
  AND U17343 ( .A(b[2]), .B(a[672]), .Z(n16467) );
  AND U17344 ( .A(a[673]), .B(b[1]), .Z(n16465) );
  AND U17345 ( .A(a[671]), .B(b[3]), .Z(n16464) );
  XOR U17346 ( .A(n16465), .B(n16464), .Z(n16466) );
  XOR U17347 ( .A(n16467), .B(n16466), .Z(n16470) );
  NAND U17348 ( .A(b[0]), .B(a[674]), .Z(n16471) );
  XOR U17349 ( .A(n16470), .B(n16471), .Z(n16473) );
  OR U17350 ( .A(n16444), .B(n16443), .Z(n16448) );
  NANDN U17351 ( .A(n16446), .B(n16445), .Z(n16447) );
  NAND U17352 ( .A(n16448), .B(n16447), .Z(n16472) );
  XNOR U17353 ( .A(n16473), .B(n16472), .Z(n16458) );
  NANDN U17354 ( .A(n16450), .B(n16449), .Z(n16454) );
  OR U17355 ( .A(n16452), .B(n16451), .Z(n16453) );
  NAND U17356 ( .A(n16454), .B(n16453), .Z(n16459) );
  XNOR U17357 ( .A(n16458), .B(n16459), .Z(n16460) );
  XNOR U17358 ( .A(n16461), .B(n16460), .Z(n16457) );
  XOR U17359 ( .A(sreg[1694]), .B(n16457), .Z(n16455) );
  XOR U17360 ( .A(n16456), .B(n16455), .Z(c[1694]) );
  NANDN U17361 ( .A(n16459), .B(n16458), .Z(n16463) );
  NAND U17362 ( .A(n16461), .B(n16460), .Z(n16462) );
  NAND U17363 ( .A(n16463), .B(n16462), .Z(n16479) );
  AND U17364 ( .A(b[2]), .B(a[673]), .Z(n16485) );
  AND U17365 ( .A(a[674]), .B(b[1]), .Z(n16483) );
  AND U17366 ( .A(a[672]), .B(b[3]), .Z(n16482) );
  XOR U17367 ( .A(n16483), .B(n16482), .Z(n16484) );
  XOR U17368 ( .A(n16485), .B(n16484), .Z(n16488) );
  NAND U17369 ( .A(b[0]), .B(a[675]), .Z(n16489) );
  XOR U17370 ( .A(n16488), .B(n16489), .Z(n16491) );
  OR U17371 ( .A(n16465), .B(n16464), .Z(n16469) );
  NANDN U17372 ( .A(n16467), .B(n16466), .Z(n16468) );
  NAND U17373 ( .A(n16469), .B(n16468), .Z(n16490) );
  XNOR U17374 ( .A(n16491), .B(n16490), .Z(n16476) );
  NANDN U17375 ( .A(n16471), .B(n16470), .Z(n16475) );
  OR U17376 ( .A(n16473), .B(n16472), .Z(n16474) );
  NAND U17377 ( .A(n16475), .B(n16474), .Z(n16477) );
  XNOR U17378 ( .A(n16476), .B(n16477), .Z(n16478) );
  XNOR U17379 ( .A(n16479), .B(n16478), .Z(n16494) );
  XNOR U17380 ( .A(n16494), .B(sreg[1695]), .Z(n16496) );
  XNOR U17381 ( .A(n16495), .B(n16496), .Z(c[1695]) );
  NANDN U17382 ( .A(n16477), .B(n16476), .Z(n16481) );
  NAND U17383 ( .A(n16479), .B(n16478), .Z(n16480) );
  NAND U17384 ( .A(n16481), .B(n16480), .Z(n16502) );
  AND U17385 ( .A(b[2]), .B(a[674]), .Z(n16508) );
  AND U17386 ( .A(a[675]), .B(b[1]), .Z(n16506) );
  AND U17387 ( .A(a[673]), .B(b[3]), .Z(n16505) );
  XOR U17388 ( .A(n16506), .B(n16505), .Z(n16507) );
  XOR U17389 ( .A(n16508), .B(n16507), .Z(n16511) );
  NAND U17390 ( .A(b[0]), .B(a[676]), .Z(n16512) );
  XOR U17391 ( .A(n16511), .B(n16512), .Z(n16514) );
  OR U17392 ( .A(n16483), .B(n16482), .Z(n16487) );
  NANDN U17393 ( .A(n16485), .B(n16484), .Z(n16486) );
  NAND U17394 ( .A(n16487), .B(n16486), .Z(n16513) );
  XNOR U17395 ( .A(n16514), .B(n16513), .Z(n16499) );
  NANDN U17396 ( .A(n16489), .B(n16488), .Z(n16493) );
  OR U17397 ( .A(n16491), .B(n16490), .Z(n16492) );
  NAND U17398 ( .A(n16493), .B(n16492), .Z(n16500) );
  XNOR U17399 ( .A(n16499), .B(n16500), .Z(n16501) );
  XNOR U17400 ( .A(n16502), .B(n16501), .Z(n16517) );
  XOR U17401 ( .A(sreg[1696]), .B(n16517), .Z(n16518) );
  NAND U17402 ( .A(n16494), .B(sreg[1695]), .Z(n16498) );
  NANDN U17403 ( .A(n16496), .B(n16495), .Z(n16497) );
  NAND U17404 ( .A(n16498), .B(n16497), .Z(n16519) );
  XOR U17405 ( .A(n16518), .B(n16519), .Z(c[1696]) );
  NANDN U17406 ( .A(n16500), .B(n16499), .Z(n16504) );
  NAND U17407 ( .A(n16502), .B(n16501), .Z(n16503) );
  NAND U17408 ( .A(n16504), .B(n16503), .Z(n16526) );
  AND U17409 ( .A(b[2]), .B(a[675]), .Z(n16532) );
  AND U17410 ( .A(a[676]), .B(b[1]), .Z(n16530) );
  AND U17411 ( .A(a[674]), .B(b[3]), .Z(n16529) );
  XOR U17412 ( .A(n16530), .B(n16529), .Z(n16531) );
  XOR U17413 ( .A(n16532), .B(n16531), .Z(n16535) );
  NAND U17414 ( .A(b[0]), .B(a[677]), .Z(n16536) );
  XOR U17415 ( .A(n16535), .B(n16536), .Z(n16538) );
  OR U17416 ( .A(n16506), .B(n16505), .Z(n16510) );
  NANDN U17417 ( .A(n16508), .B(n16507), .Z(n16509) );
  NAND U17418 ( .A(n16510), .B(n16509), .Z(n16537) );
  XNOR U17419 ( .A(n16538), .B(n16537), .Z(n16523) );
  NANDN U17420 ( .A(n16512), .B(n16511), .Z(n16516) );
  OR U17421 ( .A(n16514), .B(n16513), .Z(n16515) );
  NAND U17422 ( .A(n16516), .B(n16515), .Z(n16524) );
  XNOR U17423 ( .A(n16523), .B(n16524), .Z(n16525) );
  XOR U17424 ( .A(n16526), .B(n16525), .Z(n16542) );
  OR U17425 ( .A(n16517), .B(sreg[1696]), .Z(n16521) );
  NANDN U17426 ( .A(n16519), .B(n16518), .Z(n16520) );
  AND U17427 ( .A(n16521), .B(n16520), .Z(n16541) );
  XNOR U17428 ( .A(sreg[1697]), .B(n16541), .Z(n16522) );
  XOR U17429 ( .A(n16542), .B(n16522), .Z(c[1697]) );
  NANDN U17430 ( .A(n16524), .B(n16523), .Z(n16528) );
  NAND U17431 ( .A(n16526), .B(n16525), .Z(n16527) );
  NAND U17432 ( .A(n16528), .B(n16527), .Z(n16549) );
  AND U17433 ( .A(b[2]), .B(a[676]), .Z(n16555) );
  AND U17434 ( .A(a[677]), .B(b[1]), .Z(n16553) );
  AND U17435 ( .A(a[675]), .B(b[3]), .Z(n16552) );
  XOR U17436 ( .A(n16553), .B(n16552), .Z(n16554) );
  XOR U17437 ( .A(n16555), .B(n16554), .Z(n16558) );
  NAND U17438 ( .A(b[0]), .B(a[678]), .Z(n16559) );
  XOR U17439 ( .A(n16558), .B(n16559), .Z(n16561) );
  OR U17440 ( .A(n16530), .B(n16529), .Z(n16534) );
  NANDN U17441 ( .A(n16532), .B(n16531), .Z(n16533) );
  NAND U17442 ( .A(n16534), .B(n16533), .Z(n16560) );
  XNOR U17443 ( .A(n16561), .B(n16560), .Z(n16546) );
  NANDN U17444 ( .A(n16536), .B(n16535), .Z(n16540) );
  OR U17445 ( .A(n16538), .B(n16537), .Z(n16539) );
  NAND U17446 ( .A(n16540), .B(n16539), .Z(n16547) );
  XNOR U17447 ( .A(n16546), .B(n16547), .Z(n16548) );
  XNOR U17448 ( .A(n16549), .B(n16548), .Z(n16545) );
  XOR U17449 ( .A(n16544), .B(sreg[1698]), .Z(n16543) );
  XOR U17450 ( .A(n16545), .B(n16543), .Z(c[1698]) );
  NANDN U17451 ( .A(n16547), .B(n16546), .Z(n16551) );
  NAND U17452 ( .A(n16549), .B(n16548), .Z(n16550) );
  NAND U17453 ( .A(n16551), .B(n16550), .Z(n16567) );
  AND U17454 ( .A(b[2]), .B(a[677]), .Z(n16573) );
  AND U17455 ( .A(a[678]), .B(b[1]), .Z(n16571) );
  AND U17456 ( .A(a[676]), .B(b[3]), .Z(n16570) );
  XOR U17457 ( .A(n16571), .B(n16570), .Z(n16572) );
  XOR U17458 ( .A(n16573), .B(n16572), .Z(n16576) );
  NAND U17459 ( .A(b[0]), .B(a[679]), .Z(n16577) );
  XOR U17460 ( .A(n16576), .B(n16577), .Z(n16579) );
  OR U17461 ( .A(n16553), .B(n16552), .Z(n16557) );
  NANDN U17462 ( .A(n16555), .B(n16554), .Z(n16556) );
  NAND U17463 ( .A(n16557), .B(n16556), .Z(n16578) );
  XNOR U17464 ( .A(n16579), .B(n16578), .Z(n16564) );
  NANDN U17465 ( .A(n16559), .B(n16558), .Z(n16563) );
  OR U17466 ( .A(n16561), .B(n16560), .Z(n16562) );
  NAND U17467 ( .A(n16563), .B(n16562), .Z(n16565) );
  XNOR U17468 ( .A(n16564), .B(n16565), .Z(n16566) );
  XNOR U17469 ( .A(n16567), .B(n16566), .Z(n16582) );
  XNOR U17470 ( .A(n16582), .B(sreg[1699]), .Z(n16584) );
  XNOR U17471 ( .A(n16583), .B(n16584), .Z(c[1699]) );
  NANDN U17472 ( .A(n16565), .B(n16564), .Z(n16569) );
  NAND U17473 ( .A(n16567), .B(n16566), .Z(n16568) );
  NAND U17474 ( .A(n16569), .B(n16568), .Z(n16590) );
  AND U17475 ( .A(b[2]), .B(a[678]), .Z(n16596) );
  AND U17476 ( .A(a[679]), .B(b[1]), .Z(n16594) );
  AND U17477 ( .A(a[677]), .B(b[3]), .Z(n16593) );
  XOR U17478 ( .A(n16594), .B(n16593), .Z(n16595) );
  XOR U17479 ( .A(n16596), .B(n16595), .Z(n16599) );
  NAND U17480 ( .A(b[0]), .B(a[680]), .Z(n16600) );
  XOR U17481 ( .A(n16599), .B(n16600), .Z(n16602) );
  OR U17482 ( .A(n16571), .B(n16570), .Z(n16575) );
  NANDN U17483 ( .A(n16573), .B(n16572), .Z(n16574) );
  NAND U17484 ( .A(n16575), .B(n16574), .Z(n16601) );
  XNOR U17485 ( .A(n16602), .B(n16601), .Z(n16587) );
  NANDN U17486 ( .A(n16577), .B(n16576), .Z(n16581) );
  OR U17487 ( .A(n16579), .B(n16578), .Z(n16580) );
  NAND U17488 ( .A(n16581), .B(n16580), .Z(n16588) );
  XNOR U17489 ( .A(n16587), .B(n16588), .Z(n16589) );
  XNOR U17490 ( .A(n16590), .B(n16589), .Z(n16605) );
  XNOR U17491 ( .A(n16605), .B(sreg[1700]), .Z(n16607) );
  NAND U17492 ( .A(n16582), .B(sreg[1699]), .Z(n16586) );
  NANDN U17493 ( .A(n16584), .B(n16583), .Z(n16585) );
  AND U17494 ( .A(n16586), .B(n16585), .Z(n16606) );
  XOR U17495 ( .A(n16607), .B(n16606), .Z(c[1700]) );
  NANDN U17496 ( .A(n16588), .B(n16587), .Z(n16592) );
  NAND U17497 ( .A(n16590), .B(n16589), .Z(n16591) );
  NAND U17498 ( .A(n16592), .B(n16591), .Z(n16614) );
  AND U17499 ( .A(b[2]), .B(a[679]), .Z(n16620) );
  AND U17500 ( .A(a[680]), .B(b[1]), .Z(n16618) );
  AND U17501 ( .A(a[678]), .B(b[3]), .Z(n16617) );
  XOR U17502 ( .A(n16618), .B(n16617), .Z(n16619) );
  XOR U17503 ( .A(n16620), .B(n16619), .Z(n16623) );
  NAND U17504 ( .A(b[0]), .B(a[681]), .Z(n16624) );
  XOR U17505 ( .A(n16623), .B(n16624), .Z(n16626) );
  OR U17506 ( .A(n16594), .B(n16593), .Z(n16598) );
  NANDN U17507 ( .A(n16596), .B(n16595), .Z(n16597) );
  NAND U17508 ( .A(n16598), .B(n16597), .Z(n16625) );
  XNOR U17509 ( .A(n16626), .B(n16625), .Z(n16611) );
  NANDN U17510 ( .A(n16600), .B(n16599), .Z(n16604) );
  OR U17511 ( .A(n16602), .B(n16601), .Z(n16603) );
  NAND U17512 ( .A(n16604), .B(n16603), .Z(n16612) );
  XNOR U17513 ( .A(n16611), .B(n16612), .Z(n16613) );
  XOR U17514 ( .A(n16614), .B(n16613), .Z(n16630) );
  NAND U17515 ( .A(n16605), .B(sreg[1700]), .Z(n16609) );
  OR U17516 ( .A(n16607), .B(n16606), .Z(n16608) );
  NAND U17517 ( .A(n16609), .B(n16608), .Z(n16629) );
  XNOR U17518 ( .A(sreg[1701]), .B(n16629), .Z(n16610) );
  XOR U17519 ( .A(n16630), .B(n16610), .Z(c[1701]) );
  NANDN U17520 ( .A(n16612), .B(n16611), .Z(n16616) );
  NAND U17521 ( .A(n16614), .B(n16613), .Z(n16615) );
  NAND U17522 ( .A(n16616), .B(n16615), .Z(n16635) );
  AND U17523 ( .A(b[2]), .B(a[680]), .Z(n16641) );
  AND U17524 ( .A(a[681]), .B(b[1]), .Z(n16639) );
  AND U17525 ( .A(a[679]), .B(b[3]), .Z(n16638) );
  XOR U17526 ( .A(n16639), .B(n16638), .Z(n16640) );
  XOR U17527 ( .A(n16641), .B(n16640), .Z(n16644) );
  NAND U17528 ( .A(b[0]), .B(a[682]), .Z(n16645) );
  XOR U17529 ( .A(n16644), .B(n16645), .Z(n16647) );
  OR U17530 ( .A(n16618), .B(n16617), .Z(n16622) );
  NANDN U17531 ( .A(n16620), .B(n16619), .Z(n16621) );
  NAND U17532 ( .A(n16622), .B(n16621), .Z(n16646) );
  XNOR U17533 ( .A(n16647), .B(n16646), .Z(n16632) );
  NANDN U17534 ( .A(n16624), .B(n16623), .Z(n16628) );
  OR U17535 ( .A(n16626), .B(n16625), .Z(n16627) );
  NAND U17536 ( .A(n16628), .B(n16627), .Z(n16633) );
  XNOR U17537 ( .A(n16632), .B(n16633), .Z(n16634) );
  XNOR U17538 ( .A(n16635), .B(n16634), .Z(n16651) );
  XOR U17539 ( .A(n16650), .B(sreg[1702]), .Z(n16631) );
  XOR U17540 ( .A(n16651), .B(n16631), .Z(c[1702]) );
  NANDN U17541 ( .A(n16633), .B(n16632), .Z(n16637) );
  NAND U17542 ( .A(n16635), .B(n16634), .Z(n16636) );
  NAND U17543 ( .A(n16637), .B(n16636), .Z(n16658) );
  AND U17544 ( .A(b[2]), .B(a[681]), .Z(n16664) );
  AND U17545 ( .A(a[682]), .B(b[1]), .Z(n16662) );
  AND U17546 ( .A(a[680]), .B(b[3]), .Z(n16661) );
  XOR U17547 ( .A(n16662), .B(n16661), .Z(n16663) );
  XOR U17548 ( .A(n16664), .B(n16663), .Z(n16667) );
  NAND U17549 ( .A(b[0]), .B(a[683]), .Z(n16668) );
  XOR U17550 ( .A(n16667), .B(n16668), .Z(n16670) );
  OR U17551 ( .A(n16639), .B(n16638), .Z(n16643) );
  NANDN U17552 ( .A(n16641), .B(n16640), .Z(n16642) );
  NAND U17553 ( .A(n16643), .B(n16642), .Z(n16669) );
  XNOR U17554 ( .A(n16670), .B(n16669), .Z(n16655) );
  NANDN U17555 ( .A(n16645), .B(n16644), .Z(n16649) );
  OR U17556 ( .A(n16647), .B(n16646), .Z(n16648) );
  NAND U17557 ( .A(n16649), .B(n16648), .Z(n16656) );
  XNOR U17558 ( .A(n16655), .B(n16656), .Z(n16657) );
  XNOR U17559 ( .A(n16658), .B(n16657), .Z(n16654) );
  XOR U17560 ( .A(n16653), .B(sreg[1703]), .Z(n16652) );
  XOR U17561 ( .A(n16654), .B(n16652), .Z(c[1703]) );
  NANDN U17562 ( .A(n16656), .B(n16655), .Z(n16660) );
  NAND U17563 ( .A(n16658), .B(n16657), .Z(n16659) );
  NAND U17564 ( .A(n16660), .B(n16659), .Z(n16676) );
  AND U17565 ( .A(b[2]), .B(a[682]), .Z(n16682) );
  AND U17566 ( .A(a[683]), .B(b[1]), .Z(n16680) );
  AND U17567 ( .A(a[681]), .B(b[3]), .Z(n16679) );
  XOR U17568 ( .A(n16680), .B(n16679), .Z(n16681) );
  XOR U17569 ( .A(n16682), .B(n16681), .Z(n16685) );
  NAND U17570 ( .A(b[0]), .B(a[684]), .Z(n16686) );
  XOR U17571 ( .A(n16685), .B(n16686), .Z(n16688) );
  OR U17572 ( .A(n16662), .B(n16661), .Z(n16666) );
  NANDN U17573 ( .A(n16664), .B(n16663), .Z(n16665) );
  NAND U17574 ( .A(n16666), .B(n16665), .Z(n16687) );
  XNOR U17575 ( .A(n16688), .B(n16687), .Z(n16673) );
  NANDN U17576 ( .A(n16668), .B(n16667), .Z(n16672) );
  OR U17577 ( .A(n16670), .B(n16669), .Z(n16671) );
  NAND U17578 ( .A(n16672), .B(n16671), .Z(n16674) );
  XNOR U17579 ( .A(n16673), .B(n16674), .Z(n16675) );
  XNOR U17580 ( .A(n16676), .B(n16675), .Z(n16691) );
  XNOR U17581 ( .A(n16691), .B(sreg[1704]), .Z(n16693) );
  XNOR U17582 ( .A(n16692), .B(n16693), .Z(c[1704]) );
  NANDN U17583 ( .A(n16674), .B(n16673), .Z(n16678) );
  NAND U17584 ( .A(n16676), .B(n16675), .Z(n16677) );
  NAND U17585 ( .A(n16678), .B(n16677), .Z(n16702) );
  AND U17586 ( .A(b[2]), .B(a[683]), .Z(n16708) );
  AND U17587 ( .A(a[684]), .B(b[1]), .Z(n16706) );
  AND U17588 ( .A(a[682]), .B(b[3]), .Z(n16705) );
  XOR U17589 ( .A(n16706), .B(n16705), .Z(n16707) );
  XOR U17590 ( .A(n16708), .B(n16707), .Z(n16711) );
  NAND U17591 ( .A(b[0]), .B(a[685]), .Z(n16712) );
  XOR U17592 ( .A(n16711), .B(n16712), .Z(n16714) );
  OR U17593 ( .A(n16680), .B(n16679), .Z(n16684) );
  NANDN U17594 ( .A(n16682), .B(n16681), .Z(n16683) );
  NAND U17595 ( .A(n16684), .B(n16683), .Z(n16713) );
  XNOR U17596 ( .A(n16714), .B(n16713), .Z(n16699) );
  NANDN U17597 ( .A(n16686), .B(n16685), .Z(n16690) );
  OR U17598 ( .A(n16688), .B(n16687), .Z(n16689) );
  NAND U17599 ( .A(n16690), .B(n16689), .Z(n16700) );
  XNOR U17600 ( .A(n16699), .B(n16700), .Z(n16701) );
  XOR U17601 ( .A(n16702), .B(n16701), .Z(n16698) );
  NAND U17602 ( .A(n16691), .B(sreg[1704]), .Z(n16695) );
  NANDN U17603 ( .A(n16693), .B(n16692), .Z(n16694) );
  NAND U17604 ( .A(n16695), .B(n16694), .Z(n16697) );
  XNOR U17605 ( .A(sreg[1705]), .B(n16697), .Z(n16696) );
  XOR U17606 ( .A(n16698), .B(n16696), .Z(c[1705]) );
  NANDN U17607 ( .A(n16700), .B(n16699), .Z(n16704) );
  NAND U17608 ( .A(n16702), .B(n16701), .Z(n16703) );
  NAND U17609 ( .A(n16704), .B(n16703), .Z(n16720) );
  AND U17610 ( .A(b[2]), .B(a[684]), .Z(n16726) );
  AND U17611 ( .A(a[685]), .B(b[1]), .Z(n16724) );
  AND U17612 ( .A(a[683]), .B(b[3]), .Z(n16723) );
  XOR U17613 ( .A(n16724), .B(n16723), .Z(n16725) );
  XOR U17614 ( .A(n16726), .B(n16725), .Z(n16729) );
  NAND U17615 ( .A(b[0]), .B(a[686]), .Z(n16730) );
  XOR U17616 ( .A(n16729), .B(n16730), .Z(n16732) );
  OR U17617 ( .A(n16706), .B(n16705), .Z(n16710) );
  NANDN U17618 ( .A(n16708), .B(n16707), .Z(n16709) );
  NAND U17619 ( .A(n16710), .B(n16709), .Z(n16731) );
  XNOR U17620 ( .A(n16732), .B(n16731), .Z(n16717) );
  NANDN U17621 ( .A(n16712), .B(n16711), .Z(n16716) );
  OR U17622 ( .A(n16714), .B(n16713), .Z(n16715) );
  NAND U17623 ( .A(n16716), .B(n16715), .Z(n16718) );
  XNOR U17624 ( .A(n16717), .B(n16718), .Z(n16719) );
  XNOR U17625 ( .A(n16720), .B(n16719), .Z(n16735) );
  XNOR U17626 ( .A(n16735), .B(sreg[1706]), .Z(n16736) );
  XOR U17627 ( .A(n16737), .B(n16736), .Z(c[1706]) );
  NANDN U17628 ( .A(n16718), .B(n16717), .Z(n16722) );
  NAND U17629 ( .A(n16720), .B(n16719), .Z(n16721) );
  NAND U17630 ( .A(n16722), .B(n16721), .Z(n16746) );
  AND U17631 ( .A(b[2]), .B(a[685]), .Z(n16752) );
  AND U17632 ( .A(a[686]), .B(b[1]), .Z(n16750) );
  AND U17633 ( .A(a[684]), .B(b[3]), .Z(n16749) );
  XOR U17634 ( .A(n16750), .B(n16749), .Z(n16751) );
  XOR U17635 ( .A(n16752), .B(n16751), .Z(n16755) );
  NAND U17636 ( .A(b[0]), .B(a[687]), .Z(n16756) );
  XOR U17637 ( .A(n16755), .B(n16756), .Z(n16758) );
  OR U17638 ( .A(n16724), .B(n16723), .Z(n16728) );
  NANDN U17639 ( .A(n16726), .B(n16725), .Z(n16727) );
  NAND U17640 ( .A(n16728), .B(n16727), .Z(n16757) );
  XNOR U17641 ( .A(n16758), .B(n16757), .Z(n16743) );
  NANDN U17642 ( .A(n16730), .B(n16729), .Z(n16734) );
  OR U17643 ( .A(n16732), .B(n16731), .Z(n16733) );
  NAND U17644 ( .A(n16734), .B(n16733), .Z(n16744) );
  XNOR U17645 ( .A(n16743), .B(n16744), .Z(n16745) );
  XOR U17646 ( .A(n16746), .B(n16745), .Z(n16742) );
  NAND U17647 ( .A(n16735), .B(sreg[1706]), .Z(n16739) );
  OR U17648 ( .A(n16737), .B(n16736), .Z(n16738) );
  NAND U17649 ( .A(n16739), .B(n16738), .Z(n16741) );
  XNOR U17650 ( .A(sreg[1707]), .B(n16741), .Z(n16740) );
  XOR U17651 ( .A(n16742), .B(n16740), .Z(c[1707]) );
  NANDN U17652 ( .A(n16744), .B(n16743), .Z(n16748) );
  NAND U17653 ( .A(n16746), .B(n16745), .Z(n16747) );
  NAND U17654 ( .A(n16748), .B(n16747), .Z(n16764) );
  AND U17655 ( .A(b[2]), .B(a[686]), .Z(n16776) );
  AND U17656 ( .A(a[687]), .B(b[1]), .Z(n16774) );
  AND U17657 ( .A(a[685]), .B(b[3]), .Z(n16773) );
  XOR U17658 ( .A(n16774), .B(n16773), .Z(n16775) );
  XOR U17659 ( .A(n16776), .B(n16775), .Z(n16767) );
  NAND U17660 ( .A(b[0]), .B(a[688]), .Z(n16768) );
  XOR U17661 ( .A(n16767), .B(n16768), .Z(n16770) );
  OR U17662 ( .A(n16750), .B(n16749), .Z(n16754) );
  NANDN U17663 ( .A(n16752), .B(n16751), .Z(n16753) );
  NAND U17664 ( .A(n16754), .B(n16753), .Z(n16769) );
  XNOR U17665 ( .A(n16770), .B(n16769), .Z(n16761) );
  NANDN U17666 ( .A(n16756), .B(n16755), .Z(n16760) );
  OR U17667 ( .A(n16758), .B(n16757), .Z(n16759) );
  NAND U17668 ( .A(n16760), .B(n16759), .Z(n16762) );
  XNOR U17669 ( .A(n16761), .B(n16762), .Z(n16763) );
  XOR U17670 ( .A(n16764), .B(n16763), .Z(n16780) );
  XNOR U17671 ( .A(sreg[1708]), .B(n16780), .Z(n16781) );
  XNOR U17672 ( .A(n16782), .B(n16781), .Z(c[1708]) );
  NANDN U17673 ( .A(n16762), .B(n16761), .Z(n16766) );
  NAND U17674 ( .A(n16764), .B(n16763), .Z(n16765) );
  AND U17675 ( .A(n16766), .B(n16765), .Z(n16788) );
  NANDN U17676 ( .A(n16768), .B(n16767), .Z(n16772) );
  OR U17677 ( .A(n16770), .B(n16769), .Z(n16771) );
  AND U17678 ( .A(n16772), .B(n16771), .Z(n16787) );
  AND U17679 ( .A(b[2]), .B(a[687]), .Z(n16792) );
  AND U17680 ( .A(a[688]), .B(b[1]), .Z(n16790) );
  AND U17681 ( .A(a[686]), .B(b[3]), .Z(n16789) );
  XOR U17682 ( .A(n16790), .B(n16789), .Z(n16791) );
  XOR U17683 ( .A(n16792), .B(n16791), .Z(n16795) );
  NAND U17684 ( .A(b[0]), .B(a[689]), .Z(n16796) );
  XOR U17685 ( .A(n16795), .B(n16796), .Z(n16798) );
  OR U17686 ( .A(n16774), .B(n16773), .Z(n16778) );
  NANDN U17687 ( .A(n16776), .B(n16775), .Z(n16777) );
  NAND U17688 ( .A(n16778), .B(n16777), .Z(n16797) );
  XOR U17689 ( .A(n16798), .B(n16797), .Z(n16786) );
  XNOR U17690 ( .A(n16787), .B(n16786), .Z(n16779) );
  XOR U17691 ( .A(n16788), .B(n16779), .Z(n16802) );
  NANDN U17692 ( .A(sreg[1708]), .B(n16780), .Z(n16784) );
  NAND U17693 ( .A(n16782), .B(n16781), .Z(n16783) );
  AND U17694 ( .A(n16784), .B(n16783), .Z(n16801) );
  XNOR U17695 ( .A(sreg[1709]), .B(n16801), .Z(n16785) );
  XNOR U17696 ( .A(n16802), .B(n16785), .Z(c[1709]) );
  AND U17697 ( .A(b[2]), .B(a[688]), .Z(n16813) );
  AND U17698 ( .A(a[689]), .B(b[1]), .Z(n16811) );
  AND U17699 ( .A(a[687]), .B(b[3]), .Z(n16810) );
  XOR U17700 ( .A(n16811), .B(n16810), .Z(n16812) );
  XOR U17701 ( .A(n16813), .B(n16812), .Z(n16816) );
  NAND U17702 ( .A(b[0]), .B(a[690]), .Z(n16817) );
  XOR U17703 ( .A(n16816), .B(n16817), .Z(n16819) );
  OR U17704 ( .A(n16790), .B(n16789), .Z(n16794) );
  NANDN U17705 ( .A(n16792), .B(n16791), .Z(n16793) );
  NAND U17706 ( .A(n16794), .B(n16793), .Z(n16818) );
  XNOR U17707 ( .A(n16819), .B(n16818), .Z(n16804) );
  NANDN U17708 ( .A(n16796), .B(n16795), .Z(n16800) );
  OR U17709 ( .A(n16798), .B(n16797), .Z(n16799) );
  NAND U17710 ( .A(n16800), .B(n16799), .Z(n16805) );
  XNOR U17711 ( .A(n16804), .B(n16805), .Z(n16806) );
  XNOR U17712 ( .A(n16807), .B(n16806), .Z(n16823) );
  XOR U17713 ( .A(n16822), .B(sreg[1710]), .Z(n16803) );
  XNOR U17714 ( .A(n16823), .B(n16803), .Z(c[1710]) );
  NANDN U17715 ( .A(n16805), .B(n16804), .Z(n16809) );
  NANDN U17716 ( .A(n16807), .B(n16806), .Z(n16808) );
  NAND U17717 ( .A(n16809), .B(n16808), .Z(n16830) );
  AND U17718 ( .A(b[2]), .B(a[689]), .Z(n16836) );
  AND U17719 ( .A(a[690]), .B(b[1]), .Z(n16834) );
  AND U17720 ( .A(a[688]), .B(b[3]), .Z(n16833) );
  XOR U17721 ( .A(n16834), .B(n16833), .Z(n16835) );
  XOR U17722 ( .A(n16836), .B(n16835), .Z(n16839) );
  NAND U17723 ( .A(b[0]), .B(a[691]), .Z(n16840) );
  XOR U17724 ( .A(n16839), .B(n16840), .Z(n16842) );
  OR U17725 ( .A(n16811), .B(n16810), .Z(n16815) );
  NANDN U17726 ( .A(n16813), .B(n16812), .Z(n16814) );
  NAND U17727 ( .A(n16815), .B(n16814), .Z(n16841) );
  XNOR U17728 ( .A(n16842), .B(n16841), .Z(n16827) );
  NANDN U17729 ( .A(n16817), .B(n16816), .Z(n16821) );
  OR U17730 ( .A(n16819), .B(n16818), .Z(n16820) );
  NAND U17731 ( .A(n16821), .B(n16820), .Z(n16828) );
  XNOR U17732 ( .A(n16827), .B(n16828), .Z(n16829) );
  XOR U17733 ( .A(n16830), .B(n16829), .Z(n16826) );
  XOR U17734 ( .A(sreg[1711]), .B(n16825), .Z(n16824) );
  XOR U17735 ( .A(n16826), .B(n16824), .Z(c[1711]) );
  NANDN U17736 ( .A(n16828), .B(n16827), .Z(n16832) );
  NAND U17737 ( .A(n16830), .B(n16829), .Z(n16831) );
  AND U17738 ( .A(n16832), .B(n16831), .Z(n16848) );
  AND U17739 ( .A(b[2]), .B(a[690]), .Z(n16852) );
  AND U17740 ( .A(a[691]), .B(b[1]), .Z(n16850) );
  AND U17741 ( .A(a[689]), .B(b[3]), .Z(n16849) );
  XOR U17742 ( .A(n16850), .B(n16849), .Z(n16851) );
  XOR U17743 ( .A(n16852), .B(n16851), .Z(n16855) );
  NAND U17744 ( .A(b[0]), .B(a[692]), .Z(n16856) );
  XOR U17745 ( .A(n16855), .B(n16856), .Z(n16857) );
  OR U17746 ( .A(n16834), .B(n16833), .Z(n16838) );
  NANDN U17747 ( .A(n16836), .B(n16835), .Z(n16837) );
  AND U17748 ( .A(n16838), .B(n16837), .Z(n16858) );
  XOR U17749 ( .A(n16857), .B(n16858), .Z(n16846) );
  NANDN U17750 ( .A(n16840), .B(n16839), .Z(n16844) );
  OR U17751 ( .A(n16842), .B(n16841), .Z(n16843) );
  AND U17752 ( .A(n16844), .B(n16843), .Z(n16847) );
  XOR U17753 ( .A(n16846), .B(n16847), .Z(n16845) );
  XOR U17754 ( .A(n16848), .B(n16845), .Z(n16859) );
  XNOR U17755 ( .A(sreg[1712]), .B(n16859), .Z(n16860) );
  XOR U17756 ( .A(n16861), .B(n16860), .Z(c[1712]) );
  AND U17757 ( .A(b[2]), .B(a[691]), .Z(n16874) );
  AND U17758 ( .A(a[692]), .B(b[1]), .Z(n16872) );
  AND U17759 ( .A(a[690]), .B(b[3]), .Z(n16871) );
  XOR U17760 ( .A(n16872), .B(n16871), .Z(n16873) );
  XOR U17761 ( .A(n16874), .B(n16873), .Z(n16877) );
  NAND U17762 ( .A(b[0]), .B(a[693]), .Z(n16878) );
  XOR U17763 ( .A(n16877), .B(n16878), .Z(n16880) );
  OR U17764 ( .A(n16850), .B(n16849), .Z(n16854) );
  NANDN U17765 ( .A(n16852), .B(n16851), .Z(n16853) );
  NAND U17766 ( .A(n16854), .B(n16853), .Z(n16879) );
  XNOR U17767 ( .A(n16880), .B(n16879), .Z(n16865) );
  XNOR U17768 ( .A(n16865), .B(n16866), .Z(n16868) );
  XOR U17769 ( .A(n16867), .B(n16868), .Z(n16884) );
  NAND U17770 ( .A(sreg[1712]), .B(n16859), .Z(n16863) );
  OR U17771 ( .A(n16861), .B(n16860), .Z(n16862) );
  NAND U17772 ( .A(n16863), .B(n16862), .Z(n16883) );
  XNOR U17773 ( .A(sreg[1713]), .B(n16883), .Z(n16864) );
  XOR U17774 ( .A(n16884), .B(n16864), .Z(c[1713]) );
  NANDN U17775 ( .A(n16866), .B(n16865), .Z(n16870) );
  NAND U17776 ( .A(n16868), .B(n16867), .Z(n16869) );
  NAND U17777 ( .A(n16870), .B(n16869), .Z(n16891) );
  AND U17778 ( .A(b[2]), .B(a[692]), .Z(n16897) );
  AND U17779 ( .A(a[693]), .B(b[1]), .Z(n16895) );
  AND U17780 ( .A(a[691]), .B(b[3]), .Z(n16894) );
  XOR U17781 ( .A(n16895), .B(n16894), .Z(n16896) );
  XOR U17782 ( .A(n16897), .B(n16896), .Z(n16900) );
  NAND U17783 ( .A(b[0]), .B(a[694]), .Z(n16901) );
  XOR U17784 ( .A(n16900), .B(n16901), .Z(n16903) );
  OR U17785 ( .A(n16872), .B(n16871), .Z(n16876) );
  NANDN U17786 ( .A(n16874), .B(n16873), .Z(n16875) );
  NAND U17787 ( .A(n16876), .B(n16875), .Z(n16902) );
  XNOR U17788 ( .A(n16903), .B(n16902), .Z(n16888) );
  NANDN U17789 ( .A(n16878), .B(n16877), .Z(n16882) );
  OR U17790 ( .A(n16880), .B(n16879), .Z(n16881) );
  NAND U17791 ( .A(n16882), .B(n16881), .Z(n16889) );
  XNOR U17792 ( .A(n16888), .B(n16889), .Z(n16890) );
  XOR U17793 ( .A(n16891), .B(n16890), .Z(n16887) );
  XNOR U17794 ( .A(sreg[1714]), .B(n16886), .Z(n16885) );
  XOR U17795 ( .A(n16887), .B(n16885), .Z(c[1714]) );
  NANDN U17796 ( .A(n16889), .B(n16888), .Z(n16893) );
  NAND U17797 ( .A(n16891), .B(n16890), .Z(n16892) );
  NAND U17798 ( .A(n16893), .B(n16892), .Z(n16909) );
  AND U17799 ( .A(b[2]), .B(a[693]), .Z(n16915) );
  AND U17800 ( .A(a[694]), .B(b[1]), .Z(n16913) );
  AND U17801 ( .A(a[692]), .B(b[3]), .Z(n16912) );
  XOR U17802 ( .A(n16913), .B(n16912), .Z(n16914) );
  XOR U17803 ( .A(n16915), .B(n16914), .Z(n16918) );
  NAND U17804 ( .A(b[0]), .B(a[695]), .Z(n16919) );
  XOR U17805 ( .A(n16918), .B(n16919), .Z(n16921) );
  OR U17806 ( .A(n16895), .B(n16894), .Z(n16899) );
  NANDN U17807 ( .A(n16897), .B(n16896), .Z(n16898) );
  NAND U17808 ( .A(n16899), .B(n16898), .Z(n16920) );
  XNOR U17809 ( .A(n16921), .B(n16920), .Z(n16906) );
  NANDN U17810 ( .A(n16901), .B(n16900), .Z(n16905) );
  OR U17811 ( .A(n16903), .B(n16902), .Z(n16904) );
  NAND U17812 ( .A(n16905), .B(n16904), .Z(n16907) );
  XNOR U17813 ( .A(n16906), .B(n16907), .Z(n16908) );
  XNOR U17814 ( .A(n16909), .B(n16908), .Z(n16924) );
  XNOR U17815 ( .A(n16924), .B(sreg[1715]), .Z(n16925) );
  XOR U17816 ( .A(n16926), .B(n16925), .Z(c[1715]) );
  NANDN U17817 ( .A(n16907), .B(n16906), .Z(n16911) );
  NAND U17818 ( .A(n16909), .B(n16908), .Z(n16910) );
  NAND U17819 ( .A(n16911), .B(n16910), .Z(n16935) );
  AND U17820 ( .A(b[2]), .B(a[694]), .Z(n16941) );
  AND U17821 ( .A(a[695]), .B(b[1]), .Z(n16939) );
  AND U17822 ( .A(a[693]), .B(b[3]), .Z(n16938) );
  XOR U17823 ( .A(n16939), .B(n16938), .Z(n16940) );
  XOR U17824 ( .A(n16941), .B(n16940), .Z(n16944) );
  NAND U17825 ( .A(b[0]), .B(a[696]), .Z(n16945) );
  XOR U17826 ( .A(n16944), .B(n16945), .Z(n16947) );
  OR U17827 ( .A(n16913), .B(n16912), .Z(n16917) );
  NANDN U17828 ( .A(n16915), .B(n16914), .Z(n16916) );
  NAND U17829 ( .A(n16917), .B(n16916), .Z(n16946) );
  XNOR U17830 ( .A(n16947), .B(n16946), .Z(n16932) );
  NANDN U17831 ( .A(n16919), .B(n16918), .Z(n16923) );
  OR U17832 ( .A(n16921), .B(n16920), .Z(n16922) );
  NAND U17833 ( .A(n16923), .B(n16922), .Z(n16933) );
  XNOR U17834 ( .A(n16932), .B(n16933), .Z(n16934) );
  XOR U17835 ( .A(n16935), .B(n16934), .Z(n16931) );
  NAND U17836 ( .A(n16924), .B(sreg[1715]), .Z(n16928) );
  OR U17837 ( .A(n16926), .B(n16925), .Z(n16927) );
  NAND U17838 ( .A(n16928), .B(n16927), .Z(n16930) );
  XNOR U17839 ( .A(sreg[1716]), .B(n16930), .Z(n16929) );
  XOR U17840 ( .A(n16931), .B(n16929), .Z(c[1716]) );
  NANDN U17841 ( .A(n16933), .B(n16932), .Z(n16937) );
  NAND U17842 ( .A(n16935), .B(n16934), .Z(n16936) );
  NAND U17843 ( .A(n16937), .B(n16936), .Z(n16953) );
  AND U17844 ( .A(b[2]), .B(a[695]), .Z(n16959) );
  AND U17845 ( .A(a[696]), .B(b[1]), .Z(n16957) );
  AND U17846 ( .A(a[694]), .B(b[3]), .Z(n16956) );
  XOR U17847 ( .A(n16957), .B(n16956), .Z(n16958) );
  XOR U17848 ( .A(n16959), .B(n16958), .Z(n16962) );
  NAND U17849 ( .A(b[0]), .B(a[697]), .Z(n16963) );
  XOR U17850 ( .A(n16962), .B(n16963), .Z(n16965) );
  OR U17851 ( .A(n16939), .B(n16938), .Z(n16943) );
  NANDN U17852 ( .A(n16941), .B(n16940), .Z(n16942) );
  NAND U17853 ( .A(n16943), .B(n16942), .Z(n16964) );
  XNOR U17854 ( .A(n16965), .B(n16964), .Z(n16950) );
  NANDN U17855 ( .A(n16945), .B(n16944), .Z(n16949) );
  OR U17856 ( .A(n16947), .B(n16946), .Z(n16948) );
  NAND U17857 ( .A(n16949), .B(n16948), .Z(n16951) );
  XNOR U17858 ( .A(n16950), .B(n16951), .Z(n16952) );
  XNOR U17859 ( .A(n16953), .B(n16952), .Z(n16968) );
  XOR U17860 ( .A(sreg[1717]), .B(n16968), .Z(n16970) );
  XNOR U17861 ( .A(n16969), .B(n16970), .Z(c[1717]) );
  NANDN U17862 ( .A(n16951), .B(n16950), .Z(n16955) );
  NAND U17863 ( .A(n16953), .B(n16952), .Z(n16954) );
  NAND U17864 ( .A(n16955), .B(n16954), .Z(n16977) );
  AND U17865 ( .A(b[2]), .B(a[696]), .Z(n16983) );
  AND U17866 ( .A(a[697]), .B(b[1]), .Z(n16981) );
  AND U17867 ( .A(a[695]), .B(b[3]), .Z(n16980) );
  XOR U17868 ( .A(n16981), .B(n16980), .Z(n16982) );
  XOR U17869 ( .A(n16983), .B(n16982), .Z(n16986) );
  NAND U17870 ( .A(b[0]), .B(a[698]), .Z(n16987) );
  XOR U17871 ( .A(n16986), .B(n16987), .Z(n16989) );
  OR U17872 ( .A(n16957), .B(n16956), .Z(n16961) );
  NANDN U17873 ( .A(n16959), .B(n16958), .Z(n16960) );
  NAND U17874 ( .A(n16961), .B(n16960), .Z(n16988) );
  XNOR U17875 ( .A(n16989), .B(n16988), .Z(n16974) );
  NANDN U17876 ( .A(n16963), .B(n16962), .Z(n16967) );
  OR U17877 ( .A(n16965), .B(n16964), .Z(n16966) );
  NAND U17878 ( .A(n16967), .B(n16966), .Z(n16975) );
  XNOR U17879 ( .A(n16974), .B(n16975), .Z(n16976) );
  XOR U17880 ( .A(n16977), .B(n16976), .Z(n16993) );
  OR U17881 ( .A(n16968), .B(sreg[1717]), .Z(n16972) );
  NAND U17882 ( .A(n16970), .B(n16969), .Z(n16971) );
  AND U17883 ( .A(n16972), .B(n16971), .Z(n16992) );
  XNOR U17884 ( .A(sreg[1718]), .B(n16992), .Z(n16973) );
  XOR U17885 ( .A(n16993), .B(n16973), .Z(c[1718]) );
  NANDN U17886 ( .A(n16975), .B(n16974), .Z(n16979) );
  NAND U17887 ( .A(n16977), .B(n16976), .Z(n16978) );
  NAND U17888 ( .A(n16979), .B(n16978), .Z(n16998) );
  AND U17889 ( .A(b[2]), .B(a[697]), .Z(n17004) );
  AND U17890 ( .A(a[698]), .B(b[1]), .Z(n17002) );
  AND U17891 ( .A(a[696]), .B(b[3]), .Z(n17001) );
  XOR U17892 ( .A(n17002), .B(n17001), .Z(n17003) );
  XOR U17893 ( .A(n17004), .B(n17003), .Z(n17007) );
  NAND U17894 ( .A(b[0]), .B(a[699]), .Z(n17008) );
  XOR U17895 ( .A(n17007), .B(n17008), .Z(n17010) );
  OR U17896 ( .A(n16981), .B(n16980), .Z(n16985) );
  NANDN U17897 ( .A(n16983), .B(n16982), .Z(n16984) );
  NAND U17898 ( .A(n16985), .B(n16984), .Z(n17009) );
  XNOR U17899 ( .A(n17010), .B(n17009), .Z(n16995) );
  NANDN U17900 ( .A(n16987), .B(n16986), .Z(n16991) );
  OR U17901 ( .A(n16989), .B(n16988), .Z(n16990) );
  NAND U17902 ( .A(n16991), .B(n16990), .Z(n16996) );
  XNOR U17903 ( .A(n16995), .B(n16996), .Z(n16997) );
  XNOR U17904 ( .A(n16998), .B(n16997), .Z(n17014) );
  XOR U17905 ( .A(n17013), .B(sreg[1719]), .Z(n16994) );
  XOR U17906 ( .A(n17014), .B(n16994), .Z(c[1719]) );
  NANDN U17907 ( .A(n16996), .B(n16995), .Z(n17000) );
  NAND U17908 ( .A(n16998), .B(n16997), .Z(n16999) );
  NAND U17909 ( .A(n17000), .B(n16999), .Z(n17021) );
  AND U17910 ( .A(b[2]), .B(a[698]), .Z(n17027) );
  AND U17911 ( .A(a[699]), .B(b[1]), .Z(n17025) );
  AND U17912 ( .A(a[697]), .B(b[3]), .Z(n17024) );
  XOR U17913 ( .A(n17025), .B(n17024), .Z(n17026) );
  XOR U17914 ( .A(n17027), .B(n17026), .Z(n17030) );
  NAND U17915 ( .A(b[0]), .B(a[700]), .Z(n17031) );
  XOR U17916 ( .A(n17030), .B(n17031), .Z(n17033) );
  OR U17917 ( .A(n17002), .B(n17001), .Z(n17006) );
  NANDN U17918 ( .A(n17004), .B(n17003), .Z(n17005) );
  NAND U17919 ( .A(n17006), .B(n17005), .Z(n17032) );
  XNOR U17920 ( .A(n17033), .B(n17032), .Z(n17018) );
  NANDN U17921 ( .A(n17008), .B(n17007), .Z(n17012) );
  OR U17922 ( .A(n17010), .B(n17009), .Z(n17011) );
  NAND U17923 ( .A(n17012), .B(n17011), .Z(n17019) );
  XNOR U17924 ( .A(n17018), .B(n17019), .Z(n17020) );
  XOR U17925 ( .A(n17021), .B(n17020), .Z(n17017) );
  XOR U17926 ( .A(sreg[1720]), .B(n17016), .Z(n17015) );
  XOR U17927 ( .A(n17017), .B(n17015), .Z(c[1720]) );
  NANDN U17928 ( .A(n17019), .B(n17018), .Z(n17023) );
  NAND U17929 ( .A(n17021), .B(n17020), .Z(n17022) );
  NAND U17930 ( .A(n17023), .B(n17022), .Z(n17039) );
  AND U17931 ( .A(b[2]), .B(a[699]), .Z(n17045) );
  AND U17932 ( .A(a[700]), .B(b[1]), .Z(n17043) );
  AND U17933 ( .A(a[698]), .B(b[3]), .Z(n17042) );
  XOR U17934 ( .A(n17043), .B(n17042), .Z(n17044) );
  XOR U17935 ( .A(n17045), .B(n17044), .Z(n17048) );
  NAND U17936 ( .A(b[0]), .B(a[701]), .Z(n17049) );
  XOR U17937 ( .A(n17048), .B(n17049), .Z(n17051) );
  OR U17938 ( .A(n17025), .B(n17024), .Z(n17029) );
  NANDN U17939 ( .A(n17027), .B(n17026), .Z(n17028) );
  NAND U17940 ( .A(n17029), .B(n17028), .Z(n17050) );
  XNOR U17941 ( .A(n17051), .B(n17050), .Z(n17036) );
  NANDN U17942 ( .A(n17031), .B(n17030), .Z(n17035) );
  OR U17943 ( .A(n17033), .B(n17032), .Z(n17034) );
  NAND U17944 ( .A(n17035), .B(n17034), .Z(n17037) );
  XNOR U17945 ( .A(n17036), .B(n17037), .Z(n17038) );
  XNOR U17946 ( .A(n17039), .B(n17038), .Z(n17054) );
  XNOR U17947 ( .A(n17054), .B(sreg[1721]), .Z(n17055) );
  XOR U17948 ( .A(n17056), .B(n17055), .Z(c[1721]) );
  NANDN U17949 ( .A(n17037), .B(n17036), .Z(n17041) );
  NAND U17950 ( .A(n17039), .B(n17038), .Z(n17040) );
  NAND U17951 ( .A(n17041), .B(n17040), .Z(n17063) );
  AND U17952 ( .A(b[2]), .B(a[700]), .Z(n17069) );
  AND U17953 ( .A(a[701]), .B(b[1]), .Z(n17067) );
  AND U17954 ( .A(a[699]), .B(b[3]), .Z(n17066) );
  XOR U17955 ( .A(n17067), .B(n17066), .Z(n17068) );
  XOR U17956 ( .A(n17069), .B(n17068), .Z(n17072) );
  NAND U17957 ( .A(b[0]), .B(a[702]), .Z(n17073) );
  XOR U17958 ( .A(n17072), .B(n17073), .Z(n17075) );
  OR U17959 ( .A(n17043), .B(n17042), .Z(n17047) );
  NANDN U17960 ( .A(n17045), .B(n17044), .Z(n17046) );
  NAND U17961 ( .A(n17047), .B(n17046), .Z(n17074) );
  XNOR U17962 ( .A(n17075), .B(n17074), .Z(n17060) );
  NANDN U17963 ( .A(n17049), .B(n17048), .Z(n17053) );
  OR U17964 ( .A(n17051), .B(n17050), .Z(n17052) );
  NAND U17965 ( .A(n17053), .B(n17052), .Z(n17061) );
  XNOR U17966 ( .A(n17060), .B(n17061), .Z(n17062) );
  XOR U17967 ( .A(n17063), .B(n17062), .Z(n17079) );
  NAND U17968 ( .A(n17054), .B(sreg[1721]), .Z(n17058) );
  OR U17969 ( .A(n17056), .B(n17055), .Z(n17057) );
  NAND U17970 ( .A(n17058), .B(n17057), .Z(n17078) );
  XNOR U17971 ( .A(sreg[1722]), .B(n17078), .Z(n17059) );
  XOR U17972 ( .A(n17079), .B(n17059), .Z(c[1722]) );
  NANDN U17973 ( .A(n17061), .B(n17060), .Z(n17065) );
  NAND U17974 ( .A(n17063), .B(n17062), .Z(n17064) );
  NAND U17975 ( .A(n17065), .B(n17064), .Z(n17086) );
  AND U17976 ( .A(b[2]), .B(a[701]), .Z(n17092) );
  AND U17977 ( .A(a[702]), .B(b[1]), .Z(n17090) );
  AND U17978 ( .A(a[700]), .B(b[3]), .Z(n17089) );
  XOR U17979 ( .A(n17090), .B(n17089), .Z(n17091) );
  XOR U17980 ( .A(n17092), .B(n17091), .Z(n17095) );
  NAND U17981 ( .A(b[0]), .B(a[703]), .Z(n17096) );
  XOR U17982 ( .A(n17095), .B(n17096), .Z(n17098) );
  OR U17983 ( .A(n17067), .B(n17066), .Z(n17071) );
  NANDN U17984 ( .A(n17069), .B(n17068), .Z(n17070) );
  NAND U17985 ( .A(n17071), .B(n17070), .Z(n17097) );
  XNOR U17986 ( .A(n17098), .B(n17097), .Z(n17083) );
  NANDN U17987 ( .A(n17073), .B(n17072), .Z(n17077) );
  OR U17988 ( .A(n17075), .B(n17074), .Z(n17076) );
  NAND U17989 ( .A(n17077), .B(n17076), .Z(n17084) );
  XNOR U17990 ( .A(n17083), .B(n17084), .Z(n17085) );
  XOR U17991 ( .A(n17086), .B(n17085), .Z(n17082) );
  XNOR U17992 ( .A(sreg[1723]), .B(n17081), .Z(n17080) );
  XOR U17993 ( .A(n17082), .B(n17080), .Z(c[1723]) );
  NANDN U17994 ( .A(n17084), .B(n17083), .Z(n17088) );
  NAND U17995 ( .A(n17086), .B(n17085), .Z(n17087) );
  NAND U17996 ( .A(n17088), .B(n17087), .Z(n17104) );
  AND U17997 ( .A(b[2]), .B(a[702]), .Z(n17110) );
  AND U17998 ( .A(a[703]), .B(b[1]), .Z(n17108) );
  AND U17999 ( .A(a[701]), .B(b[3]), .Z(n17107) );
  XOR U18000 ( .A(n17108), .B(n17107), .Z(n17109) );
  XOR U18001 ( .A(n17110), .B(n17109), .Z(n17113) );
  NAND U18002 ( .A(b[0]), .B(a[704]), .Z(n17114) );
  XOR U18003 ( .A(n17113), .B(n17114), .Z(n17116) );
  OR U18004 ( .A(n17090), .B(n17089), .Z(n17094) );
  NANDN U18005 ( .A(n17092), .B(n17091), .Z(n17093) );
  NAND U18006 ( .A(n17094), .B(n17093), .Z(n17115) );
  XNOR U18007 ( .A(n17116), .B(n17115), .Z(n17101) );
  NANDN U18008 ( .A(n17096), .B(n17095), .Z(n17100) );
  OR U18009 ( .A(n17098), .B(n17097), .Z(n17099) );
  NAND U18010 ( .A(n17100), .B(n17099), .Z(n17102) );
  XNOR U18011 ( .A(n17101), .B(n17102), .Z(n17103) );
  XNOR U18012 ( .A(n17104), .B(n17103), .Z(n17119) );
  XNOR U18013 ( .A(n17119), .B(sreg[1724]), .Z(n17120) );
  XOR U18014 ( .A(n17121), .B(n17120), .Z(c[1724]) );
  NANDN U18015 ( .A(n17102), .B(n17101), .Z(n17106) );
  NAND U18016 ( .A(n17104), .B(n17103), .Z(n17105) );
  NAND U18017 ( .A(n17106), .B(n17105), .Z(n17127) );
  AND U18018 ( .A(b[2]), .B(a[703]), .Z(n17133) );
  AND U18019 ( .A(a[704]), .B(b[1]), .Z(n17131) );
  AND U18020 ( .A(a[702]), .B(b[3]), .Z(n17130) );
  XOR U18021 ( .A(n17131), .B(n17130), .Z(n17132) );
  XOR U18022 ( .A(n17133), .B(n17132), .Z(n17136) );
  NAND U18023 ( .A(b[0]), .B(a[705]), .Z(n17137) );
  XOR U18024 ( .A(n17136), .B(n17137), .Z(n17139) );
  OR U18025 ( .A(n17108), .B(n17107), .Z(n17112) );
  NANDN U18026 ( .A(n17110), .B(n17109), .Z(n17111) );
  NAND U18027 ( .A(n17112), .B(n17111), .Z(n17138) );
  XNOR U18028 ( .A(n17139), .B(n17138), .Z(n17124) );
  NANDN U18029 ( .A(n17114), .B(n17113), .Z(n17118) );
  OR U18030 ( .A(n17116), .B(n17115), .Z(n17117) );
  NAND U18031 ( .A(n17118), .B(n17117), .Z(n17125) );
  XNOR U18032 ( .A(n17124), .B(n17125), .Z(n17126) );
  XNOR U18033 ( .A(n17127), .B(n17126), .Z(n17142) );
  XOR U18034 ( .A(sreg[1725]), .B(n17142), .Z(n17143) );
  NAND U18035 ( .A(n17119), .B(sreg[1724]), .Z(n17123) );
  OR U18036 ( .A(n17121), .B(n17120), .Z(n17122) );
  NAND U18037 ( .A(n17123), .B(n17122), .Z(n17144) );
  XOR U18038 ( .A(n17143), .B(n17144), .Z(c[1725]) );
  NANDN U18039 ( .A(n17125), .B(n17124), .Z(n17129) );
  NAND U18040 ( .A(n17127), .B(n17126), .Z(n17128) );
  NAND U18041 ( .A(n17129), .B(n17128), .Z(n17155) );
  AND U18042 ( .A(b[2]), .B(a[704]), .Z(n17161) );
  AND U18043 ( .A(a[705]), .B(b[1]), .Z(n17159) );
  AND U18044 ( .A(a[703]), .B(b[3]), .Z(n17158) );
  XOR U18045 ( .A(n17159), .B(n17158), .Z(n17160) );
  XOR U18046 ( .A(n17161), .B(n17160), .Z(n17164) );
  NAND U18047 ( .A(b[0]), .B(a[706]), .Z(n17165) );
  XOR U18048 ( .A(n17164), .B(n17165), .Z(n17167) );
  OR U18049 ( .A(n17131), .B(n17130), .Z(n17135) );
  NANDN U18050 ( .A(n17133), .B(n17132), .Z(n17134) );
  NAND U18051 ( .A(n17135), .B(n17134), .Z(n17166) );
  XNOR U18052 ( .A(n17167), .B(n17166), .Z(n17152) );
  NANDN U18053 ( .A(n17137), .B(n17136), .Z(n17141) );
  OR U18054 ( .A(n17139), .B(n17138), .Z(n17140) );
  NAND U18055 ( .A(n17141), .B(n17140), .Z(n17153) );
  XNOR U18056 ( .A(n17152), .B(n17153), .Z(n17154) );
  XNOR U18057 ( .A(n17155), .B(n17154), .Z(n17147) );
  XOR U18058 ( .A(sreg[1726]), .B(n17147), .Z(n17148) );
  OR U18059 ( .A(n17142), .B(sreg[1725]), .Z(n17146) );
  NANDN U18060 ( .A(n17144), .B(n17143), .Z(n17145) );
  AND U18061 ( .A(n17146), .B(n17145), .Z(n17149) );
  XOR U18062 ( .A(n17148), .B(n17149), .Z(c[1726]) );
  OR U18063 ( .A(n17147), .B(sreg[1726]), .Z(n17151) );
  NANDN U18064 ( .A(n17149), .B(n17148), .Z(n17150) );
  AND U18065 ( .A(n17151), .B(n17150), .Z(n17171) );
  NANDN U18066 ( .A(n17153), .B(n17152), .Z(n17157) );
  NAND U18067 ( .A(n17155), .B(n17154), .Z(n17156) );
  NAND U18068 ( .A(n17157), .B(n17156), .Z(n17176) );
  AND U18069 ( .A(b[2]), .B(a[705]), .Z(n17182) );
  AND U18070 ( .A(a[706]), .B(b[1]), .Z(n17180) );
  AND U18071 ( .A(a[704]), .B(b[3]), .Z(n17179) );
  XOR U18072 ( .A(n17180), .B(n17179), .Z(n17181) );
  XOR U18073 ( .A(n17182), .B(n17181), .Z(n17185) );
  NAND U18074 ( .A(b[0]), .B(a[707]), .Z(n17186) );
  XOR U18075 ( .A(n17185), .B(n17186), .Z(n17188) );
  OR U18076 ( .A(n17159), .B(n17158), .Z(n17163) );
  NANDN U18077 ( .A(n17161), .B(n17160), .Z(n17162) );
  NAND U18078 ( .A(n17163), .B(n17162), .Z(n17187) );
  XNOR U18079 ( .A(n17188), .B(n17187), .Z(n17173) );
  NANDN U18080 ( .A(n17165), .B(n17164), .Z(n17169) );
  OR U18081 ( .A(n17167), .B(n17166), .Z(n17168) );
  NAND U18082 ( .A(n17169), .B(n17168), .Z(n17174) );
  XNOR U18083 ( .A(n17173), .B(n17174), .Z(n17175) );
  XNOR U18084 ( .A(n17176), .B(n17175), .Z(n17172) );
  XOR U18085 ( .A(sreg[1727]), .B(n17172), .Z(n17170) );
  XOR U18086 ( .A(n17171), .B(n17170), .Z(c[1727]) );
  NANDN U18087 ( .A(n17174), .B(n17173), .Z(n17178) );
  NAND U18088 ( .A(n17176), .B(n17175), .Z(n17177) );
  NAND U18089 ( .A(n17178), .B(n17177), .Z(n17199) );
  AND U18090 ( .A(b[2]), .B(a[706]), .Z(n17205) );
  AND U18091 ( .A(a[707]), .B(b[1]), .Z(n17203) );
  AND U18092 ( .A(a[705]), .B(b[3]), .Z(n17202) );
  XOR U18093 ( .A(n17203), .B(n17202), .Z(n17204) );
  XOR U18094 ( .A(n17205), .B(n17204), .Z(n17208) );
  NAND U18095 ( .A(b[0]), .B(a[708]), .Z(n17209) );
  XOR U18096 ( .A(n17208), .B(n17209), .Z(n17211) );
  OR U18097 ( .A(n17180), .B(n17179), .Z(n17184) );
  NANDN U18098 ( .A(n17182), .B(n17181), .Z(n17183) );
  NAND U18099 ( .A(n17184), .B(n17183), .Z(n17210) );
  XNOR U18100 ( .A(n17211), .B(n17210), .Z(n17196) );
  NANDN U18101 ( .A(n17186), .B(n17185), .Z(n17190) );
  OR U18102 ( .A(n17188), .B(n17187), .Z(n17189) );
  NAND U18103 ( .A(n17190), .B(n17189), .Z(n17197) );
  XNOR U18104 ( .A(n17196), .B(n17197), .Z(n17198) );
  XNOR U18105 ( .A(n17199), .B(n17198), .Z(n17191) );
  XOR U18106 ( .A(sreg[1728]), .B(n17191), .Z(n17192) );
  XOR U18107 ( .A(n17193), .B(n17192), .Z(c[1728]) );
  OR U18108 ( .A(n17191), .B(sreg[1728]), .Z(n17195) );
  NANDN U18109 ( .A(n17193), .B(n17192), .Z(n17194) );
  AND U18110 ( .A(n17195), .B(n17194), .Z(n17233) );
  NANDN U18111 ( .A(n17197), .B(n17196), .Z(n17201) );
  NAND U18112 ( .A(n17199), .B(n17198), .Z(n17200) );
  NAND U18113 ( .A(n17201), .B(n17200), .Z(n17218) );
  AND U18114 ( .A(b[2]), .B(a[707]), .Z(n17224) );
  AND U18115 ( .A(a[708]), .B(b[1]), .Z(n17222) );
  AND U18116 ( .A(a[706]), .B(b[3]), .Z(n17221) );
  XOR U18117 ( .A(n17222), .B(n17221), .Z(n17223) );
  XOR U18118 ( .A(n17224), .B(n17223), .Z(n17227) );
  NAND U18119 ( .A(b[0]), .B(a[709]), .Z(n17228) );
  XOR U18120 ( .A(n17227), .B(n17228), .Z(n17230) );
  OR U18121 ( .A(n17203), .B(n17202), .Z(n17207) );
  NANDN U18122 ( .A(n17205), .B(n17204), .Z(n17206) );
  NAND U18123 ( .A(n17207), .B(n17206), .Z(n17229) );
  XNOR U18124 ( .A(n17230), .B(n17229), .Z(n17215) );
  NANDN U18125 ( .A(n17209), .B(n17208), .Z(n17213) );
  OR U18126 ( .A(n17211), .B(n17210), .Z(n17212) );
  NAND U18127 ( .A(n17213), .B(n17212), .Z(n17216) );
  XNOR U18128 ( .A(n17215), .B(n17216), .Z(n17217) );
  XNOR U18129 ( .A(n17218), .B(n17217), .Z(n17234) );
  XOR U18130 ( .A(sreg[1729]), .B(n17234), .Z(n17214) );
  XOR U18131 ( .A(n17233), .B(n17214), .Z(c[1729]) );
  NANDN U18132 ( .A(n17216), .B(n17215), .Z(n17220) );
  NAND U18133 ( .A(n17218), .B(n17217), .Z(n17219) );
  NAND U18134 ( .A(n17220), .B(n17219), .Z(n17239) );
  AND U18135 ( .A(b[2]), .B(a[708]), .Z(n17245) );
  AND U18136 ( .A(a[709]), .B(b[1]), .Z(n17243) );
  AND U18137 ( .A(a[707]), .B(b[3]), .Z(n17242) );
  XOR U18138 ( .A(n17243), .B(n17242), .Z(n17244) );
  XOR U18139 ( .A(n17245), .B(n17244), .Z(n17248) );
  NAND U18140 ( .A(b[0]), .B(a[710]), .Z(n17249) );
  XOR U18141 ( .A(n17248), .B(n17249), .Z(n17251) );
  OR U18142 ( .A(n17222), .B(n17221), .Z(n17226) );
  NANDN U18143 ( .A(n17224), .B(n17223), .Z(n17225) );
  NAND U18144 ( .A(n17226), .B(n17225), .Z(n17250) );
  XNOR U18145 ( .A(n17251), .B(n17250), .Z(n17236) );
  NANDN U18146 ( .A(n17228), .B(n17227), .Z(n17232) );
  OR U18147 ( .A(n17230), .B(n17229), .Z(n17231) );
  NAND U18148 ( .A(n17232), .B(n17231), .Z(n17237) );
  XNOR U18149 ( .A(n17236), .B(n17237), .Z(n17238) );
  XOR U18150 ( .A(n17239), .B(n17238), .Z(n17255) );
  XOR U18151 ( .A(sreg[1730]), .B(n17254), .Z(n17235) );
  XOR U18152 ( .A(n17255), .B(n17235), .Z(c[1730]) );
  NANDN U18153 ( .A(n17237), .B(n17236), .Z(n17241) );
  NAND U18154 ( .A(n17239), .B(n17238), .Z(n17240) );
  NAND U18155 ( .A(n17241), .B(n17240), .Z(n17260) );
  AND U18156 ( .A(b[2]), .B(a[709]), .Z(n17266) );
  AND U18157 ( .A(a[710]), .B(b[1]), .Z(n17264) );
  AND U18158 ( .A(a[708]), .B(b[3]), .Z(n17263) );
  XOR U18159 ( .A(n17264), .B(n17263), .Z(n17265) );
  XOR U18160 ( .A(n17266), .B(n17265), .Z(n17269) );
  NAND U18161 ( .A(b[0]), .B(a[711]), .Z(n17270) );
  XOR U18162 ( .A(n17269), .B(n17270), .Z(n17272) );
  OR U18163 ( .A(n17243), .B(n17242), .Z(n17247) );
  NANDN U18164 ( .A(n17245), .B(n17244), .Z(n17246) );
  NAND U18165 ( .A(n17247), .B(n17246), .Z(n17271) );
  XNOR U18166 ( .A(n17272), .B(n17271), .Z(n17257) );
  NANDN U18167 ( .A(n17249), .B(n17248), .Z(n17253) );
  OR U18168 ( .A(n17251), .B(n17250), .Z(n17252) );
  NAND U18169 ( .A(n17253), .B(n17252), .Z(n17258) );
  XNOR U18170 ( .A(n17257), .B(n17258), .Z(n17259) );
  XOR U18171 ( .A(n17260), .B(n17259), .Z(n17276) );
  XNOR U18172 ( .A(sreg[1731]), .B(n17275), .Z(n17256) );
  XOR U18173 ( .A(n17276), .B(n17256), .Z(c[1731]) );
  NANDN U18174 ( .A(n17258), .B(n17257), .Z(n17262) );
  NAND U18175 ( .A(n17260), .B(n17259), .Z(n17261) );
  NAND U18176 ( .A(n17262), .B(n17261), .Z(n17283) );
  AND U18177 ( .A(b[2]), .B(a[710]), .Z(n17289) );
  AND U18178 ( .A(a[711]), .B(b[1]), .Z(n17287) );
  AND U18179 ( .A(a[709]), .B(b[3]), .Z(n17286) );
  XOR U18180 ( .A(n17287), .B(n17286), .Z(n17288) );
  XOR U18181 ( .A(n17289), .B(n17288), .Z(n17292) );
  NAND U18182 ( .A(b[0]), .B(a[712]), .Z(n17293) );
  XOR U18183 ( .A(n17292), .B(n17293), .Z(n17295) );
  OR U18184 ( .A(n17264), .B(n17263), .Z(n17268) );
  NANDN U18185 ( .A(n17266), .B(n17265), .Z(n17267) );
  NAND U18186 ( .A(n17268), .B(n17267), .Z(n17294) );
  XNOR U18187 ( .A(n17295), .B(n17294), .Z(n17280) );
  NANDN U18188 ( .A(n17270), .B(n17269), .Z(n17274) );
  OR U18189 ( .A(n17272), .B(n17271), .Z(n17273) );
  NAND U18190 ( .A(n17274), .B(n17273), .Z(n17281) );
  XNOR U18191 ( .A(n17280), .B(n17281), .Z(n17282) );
  XOR U18192 ( .A(n17283), .B(n17282), .Z(n17279) );
  XNOR U18193 ( .A(sreg[1732]), .B(n17278), .Z(n17277) );
  XOR U18194 ( .A(n17279), .B(n17277), .Z(c[1732]) );
  NANDN U18195 ( .A(n17281), .B(n17280), .Z(n17285) );
  NAND U18196 ( .A(n17283), .B(n17282), .Z(n17284) );
  NAND U18197 ( .A(n17285), .B(n17284), .Z(n17301) );
  AND U18198 ( .A(b[2]), .B(a[711]), .Z(n17307) );
  AND U18199 ( .A(a[712]), .B(b[1]), .Z(n17305) );
  AND U18200 ( .A(a[710]), .B(b[3]), .Z(n17304) );
  XOR U18201 ( .A(n17305), .B(n17304), .Z(n17306) );
  XOR U18202 ( .A(n17307), .B(n17306), .Z(n17310) );
  NAND U18203 ( .A(b[0]), .B(a[713]), .Z(n17311) );
  XOR U18204 ( .A(n17310), .B(n17311), .Z(n17313) );
  OR U18205 ( .A(n17287), .B(n17286), .Z(n17291) );
  NANDN U18206 ( .A(n17289), .B(n17288), .Z(n17290) );
  NAND U18207 ( .A(n17291), .B(n17290), .Z(n17312) );
  XNOR U18208 ( .A(n17313), .B(n17312), .Z(n17298) );
  NANDN U18209 ( .A(n17293), .B(n17292), .Z(n17297) );
  OR U18210 ( .A(n17295), .B(n17294), .Z(n17296) );
  NAND U18211 ( .A(n17297), .B(n17296), .Z(n17299) );
  XNOR U18212 ( .A(n17298), .B(n17299), .Z(n17300) );
  XNOR U18213 ( .A(n17301), .B(n17300), .Z(n17316) );
  XNOR U18214 ( .A(n17316), .B(sreg[1733]), .Z(n17317) );
  XOR U18215 ( .A(n17318), .B(n17317), .Z(c[1733]) );
  NANDN U18216 ( .A(n17299), .B(n17298), .Z(n17303) );
  NAND U18217 ( .A(n17301), .B(n17300), .Z(n17302) );
  NAND U18218 ( .A(n17303), .B(n17302), .Z(n17325) );
  AND U18219 ( .A(b[2]), .B(a[712]), .Z(n17331) );
  AND U18220 ( .A(a[713]), .B(b[1]), .Z(n17329) );
  AND U18221 ( .A(a[711]), .B(b[3]), .Z(n17328) );
  XOR U18222 ( .A(n17329), .B(n17328), .Z(n17330) );
  XOR U18223 ( .A(n17331), .B(n17330), .Z(n17334) );
  NAND U18224 ( .A(b[0]), .B(a[714]), .Z(n17335) );
  XOR U18225 ( .A(n17334), .B(n17335), .Z(n17337) );
  OR U18226 ( .A(n17305), .B(n17304), .Z(n17309) );
  NANDN U18227 ( .A(n17307), .B(n17306), .Z(n17308) );
  NAND U18228 ( .A(n17309), .B(n17308), .Z(n17336) );
  XNOR U18229 ( .A(n17337), .B(n17336), .Z(n17322) );
  NANDN U18230 ( .A(n17311), .B(n17310), .Z(n17315) );
  OR U18231 ( .A(n17313), .B(n17312), .Z(n17314) );
  NAND U18232 ( .A(n17315), .B(n17314), .Z(n17323) );
  XNOR U18233 ( .A(n17322), .B(n17323), .Z(n17324) );
  XOR U18234 ( .A(n17325), .B(n17324), .Z(n17341) );
  NAND U18235 ( .A(n17316), .B(sreg[1733]), .Z(n17320) );
  OR U18236 ( .A(n17318), .B(n17317), .Z(n17319) );
  NAND U18237 ( .A(n17320), .B(n17319), .Z(n17340) );
  XNOR U18238 ( .A(sreg[1734]), .B(n17340), .Z(n17321) );
  XOR U18239 ( .A(n17341), .B(n17321), .Z(c[1734]) );
  NANDN U18240 ( .A(n17323), .B(n17322), .Z(n17327) );
  NAND U18241 ( .A(n17325), .B(n17324), .Z(n17326) );
  NAND U18242 ( .A(n17327), .B(n17326), .Z(n17346) );
  AND U18243 ( .A(b[2]), .B(a[713]), .Z(n17352) );
  AND U18244 ( .A(a[714]), .B(b[1]), .Z(n17350) );
  AND U18245 ( .A(a[712]), .B(b[3]), .Z(n17349) );
  XOR U18246 ( .A(n17350), .B(n17349), .Z(n17351) );
  XOR U18247 ( .A(n17352), .B(n17351), .Z(n17355) );
  NAND U18248 ( .A(b[0]), .B(a[715]), .Z(n17356) );
  XOR U18249 ( .A(n17355), .B(n17356), .Z(n17358) );
  OR U18250 ( .A(n17329), .B(n17328), .Z(n17333) );
  NANDN U18251 ( .A(n17331), .B(n17330), .Z(n17332) );
  NAND U18252 ( .A(n17333), .B(n17332), .Z(n17357) );
  XNOR U18253 ( .A(n17358), .B(n17357), .Z(n17343) );
  NANDN U18254 ( .A(n17335), .B(n17334), .Z(n17339) );
  OR U18255 ( .A(n17337), .B(n17336), .Z(n17338) );
  NAND U18256 ( .A(n17339), .B(n17338), .Z(n17344) );
  XNOR U18257 ( .A(n17343), .B(n17344), .Z(n17345) );
  XNOR U18258 ( .A(n17346), .B(n17345), .Z(n17362) );
  XOR U18259 ( .A(n17361), .B(sreg[1735]), .Z(n17342) );
  XOR U18260 ( .A(n17362), .B(n17342), .Z(c[1735]) );
  NANDN U18261 ( .A(n17344), .B(n17343), .Z(n17348) );
  NAND U18262 ( .A(n17346), .B(n17345), .Z(n17347) );
  NAND U18263 ( .A(n17348), .B(n17347), .Z(n17367) );
  AND U18264 ( .A(b[2]), .B(a[714]), .Z(n17373) );
  AND U18265 ( .A(a[715]), .B(b[1]), .Z(n17371) );
  AND U18266 ( .A(a[713]), .B(b[3]), .Z(n17370) );
  XOR U18267 ( .A(n17371), .B(n17370), .Z(n17372) );
  XOR U18268 ( .A(n17373), .B(n17372), .Z(n17376) );
  NAND U18269 ( .A(b[0]), .B(a[716]), .Z(n17377) );
  XOR U18270 ( .A(n17376), .B(n17377), .Z(n17379) );
  OR U18271 ( .A(n17350), .B(n17349), .Z(n17354) );
  NANDN U18272 ( .A(n17352), .B(n17351), .Z(n17353) );
  NAND U18273 ( .A(n17354), .B(n17353), .Z(n17378) );
  XNOR U18274 ( .A(n17379), .B(n17378), .Z(n17364) );
  NANDN U18275 ( .A(n17356), .B(n17355), .Z(n17360) );
  OR U18276 ( .A(n17358), .B(n17357), .Z(n17359) );
  NAND U18277 ( .A(n17360), .B(n17359), .Z(n17365) );
  XNOR U18278 ( .A(n17364), .B(n17365), .Z(n17366) );
  XOR U18279 ( .A(n17367), .B(n17366), .Z(n17383) );
  XOR U18280 ( .A(sreg[1736]), .B(n17382), .Z(n17363) );
  XOR U18281 ( .A(n17383), .B(n17363), .Z(c[1736]) );
  NANDN U18282 ( .A(n17365), .B(n17364), .Z(n17369) );
  NAND U18283 ( .A(n17367), .B(n17366), .Z(n17368) );
  NAND U18284 ( .A(n17369), .B(n17368), .Z(n17388) );
  AND U18285 ( .A(b[2]), .B(a[715]), .Z(n17394) );
  AND U18286 ( .A(a[716]), .B(b[1]), .Z(n17392) );
  AND U18287 ( .A(a[714]), .B(b[3]), .Z(n17391) );
  XOR U18288 ( .A(n17392), .B(n17391), .Z(n17393) );
  XOR U18289 ( .A(n17394), .B(n17393), .Z(n17397) );
  NAND U18290 ( .A(b[0]), .B(a[717]), .Z(n17398) );
  XOR U18291 ( .A(n17397), .B(n17398), .Z(n17400) );
  OR U18292 ( .A(n17371), .B(n17370), .Z(n17375) );
  NANDN U18293 ( .A(n17373), .B(n17372), .Z(n17374) );
  NAND U18294 ( .A(n17375), .B(n17374), .Z(n17399) );
  XNOR U18295 ( .A(n17400), .B(n17399), .Z(n17385) );
  NANDN U18296 ( .A(n17377), .B(n17376), .Z(n17381) );
  OR U18297 ( .A(n17379), .B(n17378), .Z(n17380) );
  NAND U18298 ( .A(n17381), .B(n17380), .Z(n17386) );
  XNOR U18299 ( .A(n17385), .B(n17386), .Z(n17387) );
  XOR U18300 ( .A(n17388), .B(n17387), .Z(n17404) );
  XNOR U18301 ( .A(sreg[1737]), .B(n17403), .Z(n17384) );
  XOR U18302 ( .A(n17404), .B(n17384), .Z(c[1737]) );
  NANDN U18303 ( .A(n17386), .B(n17385), .Z(n17390) );
  NAND U18304 ( .A(n17388), .B(n17387), .Z(n17389) );
  NAND U18305 ( .A(n17390), .B(n17389), .Z(n17411) );
  AND U18306 ( .A(b[2]), .B(a[716]), .Z(n17417) );
  AND U18307 ( .A(a[717]), .B(b[1]), .Z(n17415) );
  AND U18308 ( .A(a[715]), .B(b[3]), .Z(n17414) );
  XOR U18309 ( .A(n17415), .B(n17414), .Z(n17416) );
  XOR U18310 ( .A(n17417), .B(n17416), .Z(n17420) );
  NAND U18311 ( .A(b[0]), .B(a[718]), .Z(n17421) );
  XOR U18312 ( .A(n17420), .B(n17421), .Z(n17423) );
  OR U18313 ( .A(n17392), .B(n17391), .Z(n17396) );
  NANDN U18314 ( .A(n17394), .B(n17393), .Z(n17395) );
  NAND U18315 ( .A(n17396), .B(n17395), .Z(n17422) );
  XNOR U18316 ( .A(n17423), .B(n17422), .Z(n17408) );
  NANDN U18317 ( .A(n17398), .B(n17397), .Z(n17402) );
  OR U18318 ( .A(n17400), .B(n17399), .Z(n17401) );
  NAND U18319 ( .A(n17402), .B(n17401), .Z(n17409) );
  XNOR U18320 ( .A(n17408), .B(n17409), .Z(n17410) );
  XOR U18321 ( .A(n17411), .B(n17410), .Z(n17407) );
  XNOR U18322 ( .A(sreg[1738]), .B(n17406), .Z(n17405) );
  XOR U18323 ( .A(n17407), .B(n17405), .Z(c[1738]) );
  NANDN U18324 ( .A(n17409), .B(n17408), .Z(n17413) );
  NAND U18325 ( .A(n17411), .B(n17410), .Z(n17412) );
  NAND U18326 ( .A(n17413), .B(n17412), .Z(n17429) );
  AND U18327 ( .A(b[2]), .B(a[717]), .Z(n17435) );
  AND U18328 ( .A(a[718]), .B(b[1]), .Z(n17433) );
  AND U18329 ( .A(a[716]), .B(b[3]), .Z(n17432) );
  XOR U18330 ( .A(n17433), .B(n17432), .Z(n17434) );
  XOR U18331 ( .A(n17435), .B(n17434), .Z(n17438) );
  NAND U18332 ( .A(b[0]), .B(a[719]), .Z(n17439) );
  XOR U18333 ( .A(n17438), .B(n17439), .Z(n17441) );
  OR U18334 ( .A(n17415), .B(n17414), .Z(n17419) );
  NANDN U18335 ( .A(n17417), .B(n17416), .Z(n17418) );
  NAND U18336 ( .A(n17419), .B(n17418), .Z(n17440) );
  XNOR U18337 ( .A(n17441), .B(n17440), .Z(n17426) );
  NANDN U18338 ( .A(n17421), .B(n17420), .Z(n17425) );
  OR U18339 ( .A(n17423), .B(n17422), .Z(n17424) );
  NAND U18340 ( .A(n17425), .B(n17424), .Z(n17427) );
  XNOR U18341 ( .A(n17426), .B(n17427), .Z(n17428) );
  XNOR U18342 ( .A(n17429), .B(n17428), .Z(n17444) );
  XNOR U18343 ( .A(n17444), .B(sreg[1739]), .Z(n17445) );
  XOR U18344 ( .A(n17446), .B(n17445), .Z(c[1739]) );
  NANDN U18345 ( .A(n17427), .B(n17426), .Z(n17431) );
  NAND U18346 ( .A(n17429), .B(n17428), .Z(n17430) );
  NAND U18347 ( .A(n17431), .B(n17430), .Z(n17455) );
  AND U18348 ( .A(b[2]), .B(a[718]), .Z(n17461) );
  AND U18349 ( .A(a[719]), .B(b[1]), .Z(n17459) );
  AND U18350 ( .A(a[717]), .B(b[3]), .Z(n17458) );
  XOR U18351 ( .A(n17459), .B(n17458), .Z(n17460) );
  XOR U18352 ( .A(n17461), .B(n17460), .Z(n17464) );
  NAND U18353 ( .A(b[0]), .B(a[720]), .Z(n17465) );
  XOR U18354 ( .A(n17464), .B(n17465), .Z(n17467) );
  OR U18355 ( .A(n17433), .B(n17432), .Z(n17437) );
  NANDN U18356 ( .A(n17435), .B(n17434), .Z(n17436) );
  NAND U18357 ( .A(n17437), .B(n17436), .Z(n17466) );
  XNOR U18358 ( .A(n17467), .B(n17466), .Z(n17452) );
  NANDN U18359 ( .A(n17439), .B(n17438), .Z(n17443) );
  OR U18360 ( .A(n17441), .B(n17440), .Z(n17442) );
  NAND U18361 ( .A(n17443), .B(n17442), .Z(n17453) );
  XNOR U18362 ( .A(n17452), .B(n17453), .Z(n17454) );
  XOR U18363 ( .A(n17455), .B(n17454), .Z(n17451) );
  NAND U18364 ( .A(n17444), .B(sreg[1739]), .Z(n17448) );
  OR U18365 ( .A(n17446), .B(n17445), .Z(n17447) );
  NAND U18366 ( .A(n17448), .B(n17447), .Z(n17450) );
  XNOR U18367 ( .A(sreg[1740]), .B(n17450), .Z(n17449) );
  XOR U18368 ( .A(n17451), .B(n17449), .Z(c[1740]) );
  NANDN U18369 ( .A(n17453), .B(n17452), .Z(n17457) );
  NAND U18370 ( .A(n17455), .B(n17454), .Z(n17456) );
  NAND U18371 ( .A(n17457), .B(n17456), .Z(n17473) );
  AND U18372 ( .A(b[2]), .B(a[719]), .Z(n17485) );
  AND U18373 ( .A(a[720]), .B(b[1]), .Z(n17483) );
  AND U18374 ( .A(a[718]), .B(b[3]), .Z(n17482) );
  XOR U18375 ( .A(n17483), .B(n17482), .Z(n17484) );
  XOR U18376 ( .A(n17485), .B(n17484), .Z(n17476) );
  NAND U18377 ( .A(b[0]), .B(a[721]), .Z(n17477) );
  XOR U18378 ( .A(n17476), .B(n17477), .Z(n17479) );
  OR U18379 ( .A(n17459), .B(n17458), .Z(n17463) );
  NANDN U18380 ( .A(n17461), .B(n17460), .Z(n17462) );
  NAND U18381 ( .A(n17463), .B(n17462), .Z(n17478) );
  XNOR U18382 ( .A(n17479), .B(n17478), .Z(n17470) );
  NANDN U18383 ( .A(n17465), .B(n17464), .Z(n17469) );
  OR U18384 ( .A(n17467), .B(n17466), .Z(n17468) );
  NAND U18385 ( .A(n17469), .B(n17468), .Z(n17471) );
  XNOR U18386 ( .A(n17470), .B(n17471), .Z(n17472) );
  XNOR U18387 ( .A(n17473), .B(n17472), .Z(n17489) );
  XNOR U18388 ( .A(n17489), .B(sreg[1741]), .Z(n17490) );
  XOR U18389 ( .A(n17491), .B(n17490), .Z(c[1741]) );
  NANDN U18390 ( .A(n17471), .B(n17470), .Z(n17475) );
  NAND U18391 ( .A(n17473), .B(n17472), .Z(n17474) );
  NAND U18392 ( .A(n17475), .B(n17474), .Z(n17499) );
  NANDN U18393 ( .A(n17477), .B(n17476), .Z(n17481) );
  OR U18394 ( .A(n17479), .B(n17478), .Z(n17480) );
  AND U18395 ( .A(n17481), .B(n17480), .Z(n17498) );
  AND U18396 ( .A(b[2]), .B(a[720]), .Z(n17503) );
  AND U18397 ( .A(a[721]), .B(b[1]), .Z(n17501) );
  AND U18398 ( .A(a[719]), .B(b[3]), .Z(n17500) );
  XOR U18399 ( .A(n17501), .B(n17500), .Z(n17502) );
  XOR U18400 ( .A(n17503), .B(n17502), .Z(n17506) );
  NAND U18401 ( .A(b[0]), .B(a[722]), .Z(n17507) );
  XOR U18402 ( .A(n17506), .B(n17507), .Z(n17509) );
  OR U18403 ( .A(n17483), .B(n17482), .Z(n17487) );
  NANDN U18404 ( .A(n17485), .B(n17484), .Z(n17486) );
  NAND U18405 ( .A(n17487), .B(n17486), .Z(n17508) );
  XOR U18406 ( .A(n17509), .B(n17508), .Z(n17497) );
  XNOR U18407 ( .A(n17498), .B(n17497), .Z(n17488) );
  XNOR U18408 ( .A(n17499), .B(n17488), .Z(n17496) );
  NAND U18409 ( .A(n17489), .B(sreg[1741]), .Z(n17493) );
  OR U18410 ( .A(n17491), .B(n17490), .Z(n17492) );
  AND U18411 ( .A(n17493), .B(n17492), .Z(n17495) );
  XNOR U18412 ( .A(n17495), .B(sreg[1742]), .Z(n17494) );
  XOR U18413 ( .A(n17496), .B(n17494), .Z(c[1742]) );
  AND U18414 ( .A(b[2]), .B(a[721]), .Z(n17521) );
  AND U18415 ( .A(a[722]), .B(b[1]), .Z(n17519) );
  AND U18416 ( .A(a[720]), .B(b[3]), .Z(n17518) );
  XOR U18417 ( .A(n17519), .B(n17518), .Z(n17520) );
  XOR U18418 ( .A(n17521), .B(n17520), .Z(n17524) );
  NAND U18419 ( .A(b[0]), .B(a[723]), .Z(n17525) );
  XOR U18420 ( .A(n17524), .B(n17525), .Z(n17527) );
  OR U18421 ( .A(n17501), .B(n17500), .Z(n17505) );
  NANDN U18422 ( .A(n17503), .B(n17502), .Z(n17504) );
  NAND U18423 ( .A(n17505), .B(n17504), .Z(n17526) );
  XNOR U18424 ( .A(n17527), .B(n17526), .Z(n17512) );
  NANDN U18425 ( .A(n17507), .B(n17506), .Z(n17511) );
  OR U18426 ( .A(n17509), .B(n17508), .Z(n17510) );
  NAND U18427 ( .A(n17511), .B(n17510), .Z(n17513) );
  XNOR U18428 ( .A(n17512), .B(n17513), .Z(n17514) );
  XOR U18429 ( .A(n17515), .B(n17514), .Z(n17530) );
  XNOR U18430 ( .A(n17530), .B(sreg[1743]), .Z(n17532) );
  XNOR U18431 ( .A(n17531), .B(n17532), .Z(c[1743]) );
  NANDN U18432 ( .A(n17513), .B(n17512), .Z(n17517) );
  NANDN U18433 ( .A(n17515), .B(n17514), .Z(n17516) );
  NAND U18434 ( .A(n17517), .B(n17516), .Z(n17538) );
  AND U18435 ( .A(b[2]), .B(a[722]), .Z(n17544) );
  AND U18436 ( .A(a[723]), .B(b[1]), .Z(n17542) );
  AND U18437 ( .A(a[721]), .B(b[3]), .Z(n17541) );
  XOR U18438 ( .A(n17542), .B(n17541), .Z(n17543) );
  XOR U18439 ( .A(n17544), .B(n17543), .Z(n17547) );
  NAND U18440 ( .A(b[0]), .B(a[724]), .Z(n17548) );
  XOR U18441 ( .A(n17547), .B(n17548), .Z(n17550) );
  OR U18442 ( .A(n17519), .B(n17518), .Z(n17523) );
  NANDN U18443 ( .A(n17521), .B(n17520), .Z(n17522) );
  NAND U18444 ( .A(n17523), .B(n17522), .Z(n17549) );
  XNOR U18445 ( .A(n17550), .B(n17549), .Z(n17535) );
  NANDN U18446 ( .A(n17525), .B(n17524), .Z(n17529) );
  OR U18447 ( .A(n17527), .B(n17526), .Z(n17528) );
  NAND U18448 ( .A(n17529), .B(n17528), .Z(n17536) );
  XNOR U18449 ( .A(n17535), .B(n17536), .Z(n17537) );
  XNOR U18450 ( .A(n17538), .B(n17537), .Z(n17553) );
  XNOR U18451 ( .A(n17553), .B(sreg[1744]), .Z(n17555) );
  NAND U18452 ( .A(n17530), .B(sreg[1743]), .Z(n17534) );
  NANDN U18453 ( .A(n17532), .B(n17531), .Z(n17533) );
  AND U18454 ( .A(n17534), .B(n17533), .Z(n17554) );
  XOR U18455 ( .A(n17555), .B(n17554), .Z(c[1744]) );
  NANDN U18456 ( .A(n17536), .B(n17535), .Z(n17540) );
  NAND U18457 ( .A(n17538), .B(n17537), .Z(n17539) );
  NAND U18458 ( .A(n17540), .B(n17539), .Z(n17561) );
  AND U18459 ( .A(b[2]), .B(a[723]), .Z(n17567) );
  AND U18460 ( .A(a[724]), .B(b[1]), .Z(n17565) );
  AND U18461 ( .A(a[722]), .B(b[3]), .Z(n17564) );
  XOR U18462 ( .A(n17565), .B(n17564), .Z(n17566) );
  XOR U18463 ( .A(n17567), .B(n17566), .Z(n17570) );
  NAND U18464 ( .A(b[0]), .B(a[725]), .Z(n17571) );
  XOR U18465 ( .A(n17570), .B(n17571), .Z(n17573) );
  OR U18466 ( .A(n17542), .B(n17541), .Z(n17546) );
  NANDN U18467 ( .A(n17544), .B(n17543), .Z(n17545) );
  NAND U18468 ( .A(n17546), .B(n17545), .Z(n17572) );
  XNOR U18469 ( .A(n17573), .B(n17572), .Z(n17558) );
  NANDN U18470 ( .A(n17548), .B(n17547), .Z(n17552) );
  OR U18471 ( .A(n17550), .B(n17549), .Z(n17551) );
  NAND U18472 ( .A(n17552), .B(n17551), .Z(n17559) );
  XNOR U18473 ( .A(n17558), .B(n17559), .Z(n17560) );
  XNOR U18474 ( .A(n17561), .B(n17560), .Z(n17576) );
  XNOR U18475 ( .A(n17576), .B(sreg[1745]), .Z(n17578) );
  NAND U18476 ( .A(n17553), .B(sreg[1744]), .Z(n17557) );
  OR U18477 ( .A(n17555), .B(n17554), .Z(n17556) );
  AND U18478 ( .A(n17557), .B(n17556), .Z(n17577) );
  XOR U18479 ( .A(n17578), .B(n17577), .Z(c[1745]) );
  NANDN U18480 ( .A(n17559), .B(n17558), .Z(n17563) );
  NAND U18481 ( .A(n17561), .B(n17560), .Z(n17562) );
  NAND U18482 ( .A(n17563), .B(n17562), .Z(n17584) );
  AND U18483 ( .A(b[2]), .B(a[724]), .Z(n17590) );
  AND U18484 ( .A(a[725]), .B(b[1]), .Z(n17588) );
  AND U18485 ( .A(a[723]), .B(b[3]), .Z(n17587) );
  XOR U18486 ( .A(n17588), .B(n17587), .Z(n17589) );
  XOR U18487 ( .A(n17590), .B(n17589), .Z(n17593) );
  NAND U18488 ( .A(b[0]), .B(a[726]), .Z(n17594) );
  XOR U18489 ( .A(n17593), .B(n17594), .Z(n17596) );
  OR U18490 ( .A(n17565), .B(n17564), .Z(n17569) );
  NANDN U18491 ( .A(n17567), .B(n17566), .Z(n17568) );
  NAND U18492 ( .A(n17569), .B(n17568), .Z(n17595) );
  XNOR U18493 ( .A(n17596), .B(n17595), .Z(n17581) );
  NANDN U18494 ( .A(n17571), .B(n17570), .Z(n17575) );
  OR U18495 ( .A(n17573), .B(n17572), .Z(n17574) );
  NAND U18496 ( .A(n17575), .B(n17574), .Z(n17582) );
  XNOR U18497 ( .A(n17581), .B(n17582), .Z(n17583) );
  XNOR U18498 ( .A(n17584), .B(n17583), .Z(n17599) );
  XNOR U18499 ( .A(n17599), .B(sreg[1746]), .Z(n17601) );
  NAND U18500 ( .A(n17576), .B(sreg[1745]), .Z(n17580) );
  OR U18501 ( .A(n17578), .B(n17577), .Z(n17579) );
  AND U18502 ( .A(n17580), .B(n17579), .Z(n17600) );
  XOR U18503 ( .A(n17601), .B(n17600), .Z(c[1746]) );
  NANDN U18504 ( .A(n17582), .B(n17581), .Z(n17586) );
  NAND U18505 ( .A(n17584), .B(n17583), .Z(n17585) );
  NAND U18506 ( .A(n17586), .B(n17585), .Z(n17607) );
  AND U18507 ( .A(b[2]), .B(a[725]), .Z(n17613) );
  AND U18508 ( .A(a[726]), .B(b[1]), .Z(n17611) );
  AND U18509 ( .A(a[724]), .B(b[3]), .Z(n17610) );
  XOR U18510 ( .A(n17611), .B(n17610), .Z(n17612) );
  XOR U18511 ( .A(n17613), .B(n17612), .Z(n17616) );
  NAND U18512 ( .A(b[0]), .B(a[727]), .Z(n17617) );
  XOR U18513 ( .A(n17616), .B(n17617), .Z(n17619) );
  OR U18514 ( .A(n17588), .B(n17587), .Z(n17592) );
  NANDN U18515 ( .A(n17590), .B(n17589), .Z(n17591) );
  NAND U18516 ( .A(n17592), .B(n17591), .Z(n17618) );
  XNOR U18517 ( .A(n17619), .B(n17618), .Z(n17604) );
  NANDN U18518 ( .A(n17594), .B(n17593), .Z(n17598) );
  OR U18519 ( .A(n17596), .B(n17595), .Z(n17597) );
  NAND U18520 ( .A(n17598), .B(n17597), .Z(n17605) );
  XNOR U18521 ( .A(n17604), .B(n17605), .Z(n17606) );
  XNOR U18522 ( .A(n17607), .B(n17606), .Z(n17622) );
  XNOR U18523 ( .A(n17622), .B(sreg[1747]), .Z(n17624) );
  NAND U18524 ( .A(n17599), .B(sreg[1746]), .Z(n17603) );
  OR U18525 ( .A(n17601), .B(n17600), .Z(n17602) );
  AND U18526 ( .A(n17603), .B(n17602), .Z(n17623) );
  XOR U18527 ( .A(n17624), .B(n17623), .Z(c[1747]) );
  NANDN U18528 ( .A(n17605), .B(n17604), .Z(n17609) );
  NAND U18529 ( .A(n17607), .B(n17606), .Z(n17608) );
  NAND U18530 ( .A(n17609), .B(n17608), .Z(n17630) );
  AND U18531 ( .A(b[2]), .B(a[726]), .Z(n17636) );
  AND U18532 ( .A(a[727]), .B(b[1]), .Z(n17634) );
  AND U18533 ( .A(a[725]), .B(b[3]), .Z(n17633) );
  XOR U18534 ( .A(n17634), .B(n17633), .Z(n17635) );
  XOR U18535 ( .A(n17636), .B(n17635), .Z(n17639) );
  NAND U18536 ( .A(b[0]), .B(a[728]), .Z(n17640) );
  XOR U18537 ( .A(n17639), .B(n17640), .Z(n17642) );
  OR U18538 ( .A(n17611), .B(n17610), .Z(n17615) );
  NANDN U18539 ( .A(n17613), .B(n17612), .Z(n17614) );
  NAND U18540 ( .A(n17615), .B(n17614), .Z(n17641) );
  XNOR U18541 ( .A(n17642), .B(n17641), .Z(n17627) );
  NANDN U18542 ( .A(n17617), .B(n17616), .Z(n17621) );
  OR U18543 ( .A(n17619), .B(n17618), .Z(n17620) );
  NAND U18544 ( .A(n17621), .B(n17620), .Z(n17628) );
  XNOR U18545 ( .A(n17627), .B(n17628), .Z(n17629) );
  XNOR U18546 ( .A(n17630), .B(n17629), .Z(n17645) );
  XNOR U18547 ( .A(n17645), .B(sreg[1748]), .Z(n17647) );
  NAND U18548 ( .A(n17622), .B(sreg[1747]), .Z(n17626) );
  OR U18549 ( .A(n17624), .B(n17623), .Z(n17625) );
  AND U18550 ( .A(n17626), .B(n17625), .Z(n17646) );
  XOR U18551 ( .A(n17647), .B(n17646), .Z(c[1748]) );
  NANDN U18552 ( .A(n17628), .B(n17627), .Z(n17632) );
  NAND U18553 ( .A(n17630), .B(n17629), .Z(n17631) );
  NAND U18554 ( .A(n17632), .B(n17631), .Z(n17656) );
  AND U18555 ( .A(b[2]), .B(a[727]), .Z(n17662) );
  AND U18556 ( .A(a[728]), .B(b[1]), .Z(n17660) );
  AND U18557 ( .A(a[726]), .B(b[3]), .Z(n17659) );
  XOR U18558 ( .A(n17660), .B(n17659), .Z(n17661) );
  XOR U18559 ( .A(n17662), .B(n17661), .Z(n17665) );
  NAND U18560 ( .A(b[0]), .B(a[729]), .Z(n17666) );
  XOR U18561 ( .A(n17665), .B(n17666), .Z(n17668) );
  OR U18562 ( .A(n17634), .B(n17633), .Z(n17638) );
  NANDN U18563 ( .A(n17636), .B(n17635), .Z(n17637) );
  NAND U18564 ( .A(n17638), .B(n17637), .Z(n17667) );
  XNOR U18565 ( .A(n17668), .B(n17667), .Z(n17653) );
  NANDN U18566 ( .A(n17640), .B(n17639), .Z(n17644) );
  OR U18567 ( .A(n17642), .B(n17641), .Z(n17643) );
  NAND U18568 ( .A(n17644), .B(n17643), .Z(n17654) );
  XNOR U18569 ( .A(n17653), .B(n17654), .Z(n17655) );
  XOR U18570 ( .A(n17656), .B(n17655), .Z(n17652) );
  NAND U18571 ( .A(n17645), .B(sreg[1748]), .Z(n17649) );
  OR U18572 ( .A(n17647), .B(n17646), .Z(n17648) );
  NAND U18573 ( .A(n17649), .B(n17648), .Z(n17651) );
  XNOR U18574 ( .A(sreg[1749]), .B(n17651), .Z(n17650) );
  XOR U18575 ( .A(n17652), .B(n17650), .Z(c[1749]) );
  NANDN U18576 ( .A(n17654), .B(n17653), .Z(n17658) );
  NAND U18577 ( .A(n17656), .B(n17655), .Z(n17657) );
  NAND U18578 ( .A(n17658), .B(n17657), .Z(n17679) );
  AND U18579 ( .A(b[2]), .B(a[728]), .Z(n17685) );
  AND U18580 ( .A(a[729]), .B(b[1]), .Z(n17683) );
  AND U18581 ( .A(a[727]), .B(b[3]), .Z(n17682) );
  XOR U18582 ( .A(n17683), .B(n17682), .Z(n17684) );
  XOR U18583 ( .A(n17685), .B(n17684), .Z(n17688) );
  NAND U18584 ( .A(b[0]), .B(a[730]), .Z(n17689) );
  XOR U18585 ( .A(n17688), .B(n17689), .Z(n17691) );
  OR U18586 ( .A(n17660), .B(n17659), .Z(n17664) );
  NANDN U18587 ( .A(n17662), .B(n17661), .Z(n17663) );
  NAND U18588 ( .A(n17664), .B(n17663), .Z(n17690) );
  XNOR U18589 ( .A(n17691), .B(n17690), .Z(n17676) );
  NANDN U18590 ( .A(n17666), .B(n17665), .Z(n17670) );
  OR U18591 ( .A(n17668), .B(n17667), .Z(n17669) );
  NAND U18592 ( .A(n17670), .B(n17669), .Z(n17677) );
  XNOR U18593 ( .A(n17676), .B(n17677), .Z(n17678) );
  XNOR U18594 ( .A(n17679), .B(n17678), .Z(n17671) );
  XNOR U18595 ( .A(n17671), .B(sreg[1750]), .Z(n17672) );
  XOR U18596 ( .A(n17673), .B(n17672), .Z(c[1750]) );
  NAND U18597 ( .A(n17671), .B(sreg[1750]), .Z(n17675) );
  OR U18598 ( .A(n17673), .B(n17672), .Z(n17674) );
  NAND U18599 ( .A(n17675), .B(n17674), .Z(n17714) );
  NANDN U18600 ( .A(n17677), .B(n17676), .Z(n17681) );
  NAND U18601 ( .A(n17679), .B(n17678), .Z(n17680) );
  NAND U18602 ( .A(n17681), .B(n17680), .Z(n17697) );
  AND U18603 ( .A(b[2]), .B(a[729]), .Z(n17703) );
  AND U18604 ( .A(a[730]), .B(b[1]), .Z(n17701) );
  AND U18605 ( .A(a[728]), .B(b[3]), .Z(n17700) );
  XOR U18606 ( .A(n17701), .B(n17700), .Z(n17702) );
  XOR U18607 ( .A(n17703), .B(n17702), .Z(n17706) );
  NAND U18608 ( .A(b[0]), .B(a[731]), .Z(n17707) );
  XOR U18609 ( .A(n17706), .B(n17707), .Z(n17709) );
  OR U18610 ( .A(n17683), .B(n17682), .Z(n17687) );
  NANDN U18611 ( .A(n17685), .B(n17684), .Z(n17686) );
  NAND U18612 ( .A(n17687), .B(n17686), .Z(n17708) );
  XNOR U18613 ( .A(n17709), .B(n17708), .Z(n17694) );
  NANDN U18614 ( .A(n17689), .B(n17688), .Z(n17693) );
  OR U18615 ( .A(n17691), .B(n17690), .Z(n17692) );
  NAND U18616 ( .A(n17693), .B(n17692), .Z(n17695) );
  XNOR U18617 ( .A(n17694), .B(n17695), .Z(n17696) );
  XNOR U18618 ( .A(n17697), .B(n17696), .Z(n17712) );
  XOR U18619 ( .A(sreg[1751]), .B(n17712), .Z(n17713) );
  XOR U18620 ( .A(n17714), .B(n17713), .Z(c[1751]) );
  NANDN U18621 ( .A(n17695), .B(n17694), .Z(n17699) );
  NAND U18622 ( .A(n17697), .B(n17696), .Z(n17698) );
  NAND U18623 ( .A(n17699), .B(n17698), .Z(n17723) );
  AND U18624 ( .A(b[2]), .B(a[730]), .Z(n17729) );
  AND U18625 ( .A(a[731]), .B(b[1]), .Z(n17727) );
  AND U18626 ( .A(a[729]), .B(b[3]), .Z(n17726) );
  XOR U18627 ( .A(n17727), .B(n17726), .Z(n17728) );
  XOR U18628 ( .A(n17729), .B(n17728), .Z(n17732) );
  NAND U18629 ( .A(b[0]), .B(a[732]), .Z(n17733) );
  XOR U18630 ( .A(n17732), .B(n17733), .Z(n17735) );
  OR U18631 ( .A(n17701), .B(n17700), .Z(n17705) );
  NANDN U18632 ( .A(n17703), .B(n17702), .Z(n17704) );
  NAND U18633 ( .A(n17705), .B(n17704), .Z(n17734) );
  XNOR U18634 ( .A(n17735), .B(n17734), .Z(n17720) );
  NANDN U18635 ( .A(n17707), .B(n17706), .Z(n17711) );
  OR U18636 ( .A(n17709), .B(n17708), .Z(n17710) );
  NAND U18637 ( .A(n17711), .B(n17710), .Z(n17721) );
  XNOR U18638 ( .A(n17720), .B(n17721), .Z(n17722) );
  XOR U18639 ( .A(n17723), .B(n17722), .Z(n17719) );
  OR U18640 ( .A(n17712), .B(sreg[1751]), .Z(n17716) );
  NANDN U18641 ( .A(n17714), .B(n17713), .Z(n17715) );
  AND U18642 ( .A(n17716), .B(n17715), .Z(n17718) );
  XNOR U18643 ( .A(sreg[1752]), .B(n17718), .Z(n17717) );
  XOR U18644 ( .A(n17719), .B(n17717), .Z(c[1752]) );
  NANDN U18645 ( .A(n17721), .B(n17720), .Z(n17725) );
  NAND U18646 ( .A(n17723), .B(n17722), .Z(n17724) );
  NAND U18647 ( .A(n17725), .B(n17724), .Z(n17741) );
  AND U18648 ( .A(b[2]), .B(a[731]), .Z(n17747) );
  AND U18649 ( .A(a[732]), .B(b[1]), .Z(n17745) );
  AND U18650 ( .A(a[730]), .B(b[3]), .Z(n17744) );
  XOR U18651 ( .A(n17745), .B(n17744), .Z(n17746) );
  XOR U18652 ( .A(n17747), .B(n17746), .Z(n17750) );
  NAND U18653 ( .A(b[0]), .B(a[733]), .Z(n17751) );
  XOR U18654 ( .A(n17750), .B(n17751), .Z(n17753) );
  OR U18655 ( .A(n17727), .B(n17726), .Z(n17731) );
  NANDN U18656 ( .A(n17729), .B(n17728), .Z(n17730) );
  NAND U18657 ( .A(n17731), .B(n17730), .Z(n17752) );
  XNOR U18658 ( .A(n17753), .B(n17752), .Z(n17738) );
  NANDN U18659 ( .A(n17733), .B(n17732), .Z(n17737) );
  OR U18660 ( .A(n17735), .B(n17734), .Z(n17736) );
  NAND U18661 ( .A(n17737), .B(n17736), .Z(n17739) );
  XNOR U18662 ( .A(n17738), .B(n17739), .Z(n17740) );
  XNOR U18663 ( .A(n17741), .B(n17740), .Z(n17756) );
  XNOR U18664 ( .A(n17756), .B(sreg[1753]), .Z(n17757) );
  XOR U18665 ( .A(n17758), .B(n17757), .Z(c[1753]) );
  NANDN U18666 ( .A(n17739), .B(n17738), .Z(n17743) );
  NAND U18667 ( .A(n17741), .B(n17740), .Z(n17742) );
  NAND U18668 ( .A(n17743), .B(n17742), .Z(n17764) );
  AND U18669 ( .A(b[2]), .B(a[732]), .Z(n17770) );
  AND U18670 ( .A(a[733]), .B(b[1]), .Z(n17768) );
  AND U18671 ( .A(a[731]), .B(b[3]), .Z(n17767) );
  XOR U18672 ( .A(n17768), .B(n17767), .Z(n17769) );
  XOR U18673 ( .A(n17770), .B(n17769), .Z(n17773) );
  NAND U18674 ( .A(b[0]), .B(a[734]), .Z(n17774) );
  XOR U18675 ( .A(n17773), .B(n17774), .Z(n17776) );
  OR U18676 ( .A(n17745), .B(n17744), .Z(n17749) );
  NANDN U18677 ( .A(n17747), .B(n17746), .Z(n17748) );
  NAND U18678 ( .A(n17749), .B(n17748), .Z(n17775) );
  XNOR U18679 ( .A(n17776), .B(n17775), .Z(n17761) );
  NANDN U18680 ( .A(n17751), .B(n17750), .Z(n17755) );
  OR U18681 ( .A(n17753), .B(n17752), .Z(n17754) );
  NAND U18682 ( .A(n17755), .B(n17754), .Z(n17762) );
  XNOR U18683 ( .A(n17761), .B(n17762), .Z(n17763) );
  XNOR U18684 ( .A(n17764), .B(n17763), .Z(n17779) );
  XOR U18685 ( .A(sreg[1754]), .B(n17779), .Z(n17780) );
  NAND U18686 ( .A(n17756), .B(sreg[1753]), .Z(n17760) );
  OR U18687 ( .A(n17758), .B(n17757), .Z(n17759) );
  NAND U18688 ( .A(n17760), .B(n17759), .Z(n17781) );
  XOR U18689 ( .A(n17780), .B(n17781), .Z(c[1754]) );
  NANDN U18690 ( .A(n17762), .B(n17761), .Z(n17766) );
  NAND U18691 ( .A(n17764), .B(n17763), .Z(n17765) );
  NAND U18692 ( .A(n17766), .B(n17765), .Z(n17790) );
  AND U18693 ( .A(b[2]), .B(a[733]), .Z(n17796) );
  AND U18694 ( .A(a[734]), .B(b[1]), .Z(n17794) );
  AND U18695 ( .A(a[732]), .B(b[3]), .Z(n17793) );
  XOR U18696 ( .A(n17794), .B(n17793), .Z(n17795) );
  XOR U18697 ( .A(n17796), .B(n17795), .Z(n17799) );
  NAND U18698 ( .A(b[0]), .B(a[735]), .Z(n17800) );
  XOR U18699 ( .A(n17799), .B(n17800), .Z(n17802) );
  OR U18700 ( .A(n17768), .B(n17767), .Z(n17772) );
  NANDN U18701 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18702 ( .A(n17772), .B(n17771), .Z(n17801) );
  XNOR U18703 ( .A(n17802), .B(n17801), .Z(n17787) );
  NANDN U18704 ( .A(n17774), .B(n17773), .Z(n17778) );
  OR U18705 ( .A(n17776), .B(n17775), .Z(n17777) );
  NAND U18706 ( .A(n17778), .B(n17777), .Z(n17788) );
  XNOR U18707 ( .A(n17787), .B(n17788), .Z(n17789) );
  XOR U18708 ( .A(n17790), .B(n17789), .Z(n17786) );
  OR U18709 ( .A(n17779), .B(sreg[1754]), .Z(n17783) );
  NANDN U18710 ( .A(n17781), .B(n17780), .Z(n17782) );
  AND U18711 ( .A(n17783), .B(n17782), .Z(n17785) );
  XNOR U18712 ( .A(sreg[1755]), .B(n17785), .Z(n17784) );
  XOR U18713 ( .A(n17786), .B(n17784), .Z(c[1755]) );
  NANDN U18714 ( .A(n17788), .B(n17787), .Z(n17792) );
  NAND U18715 ( .A(n17790), .B(n17789), .Z(n17791) );
  NAND U18716 ( .A(n17792), .B(n17791), .Z(n17808) );
  AND U18717 ( .A(b[2]), .B(a[734]), .Z(n17814) );
  AND U18718 ( .A(a[735]), .B(b[1]), .Z(n17812) );
  AND U18719 ( .A(a[733]), .B(b[3]), .Z(n17811) );
  XOR U18720 ( .A(n17812), .B(n17811), .Z(n17813) );
  XOR U18721 ( .A(n17814), .B(n17813), .Z(n17817) );
  NAND U18722 ( .A(b[0]), .B(a[736]), .Z(n17818) );
  XOR U18723 ( .A(n17817), .B(n17818), .Z(n17820) );
  OR U18724 ( .A(n17794), .B(n17793), .Z(n17798) );
  NANDN U18725 ( .A(n17796), .B(n17795), .Z(n17797) );
  NAND U18726 ( .A(n17798), .B(n17797), .Z(n17819) );
  XNOR U18727 ( .A(n17820), .B(n17819), .Z(n17805) );
  NANDN U18728 ( .A(n17800), .B(n17799), .Z(n17804) );
  OR U18729 ( .A(n17802), .B(n17801), .Z(n17803) );
  NAND U18730 ( .A(n17804), .B(n17803), .Z(n17806) );
  XNOR U18731 ( .A(n17805), .B(n17806), .Z(n17807) );
  XNOR U18732 ( .A(n17808), .B(n17807), .Z(n17823) );
  XNOR U18733 ( .A(n17823), .B(sreg[1756]), .Z(n17824) );
  XOR U18734 ( .A(n17825), .B(n17824), .Z(c[1756]) );
  NANDN U18735 ( .A(n17806), .B(n17805), .Z(n17810) );
  NAND U18736 ( .A(n17808), .B(n17807), .Z(n17809) );
  NAND U18737 ( .A(n17810), .B(n17809), .Z(n17836) );
  AND U18738 ( .A(b[2]), .B(a[735]), .Z(n17842) );
  AND U18739 ( .A(a[736]), .B(b[1]), .Z(n17840) );
  AND U18740 ( .A(a[734]), .B(b[3]), .Z(n17839) );
  XOR U18741 ( .A(n17840), .B(n17839), .Z(n17841) );
  XOR U18742 ( .A(n17842), .B(n17841), .Z(n17845) );
  NAND U18743 ( .A(b[0]), .B(a[737]), .Z(n17846) );
  XOR U18744 ( .A(n17845), .B(n17846), .Z(n17848) );
  OR U18745 ( .A(n17812), .B(n17811), .Z(n17816) );
  NANDN U18746 ( .A(n17814), .B(n17813), .Z(n17815) );
  NAND U18747 ( .A(n17816), .B(n17815), .Z(n17847) );
  XNOR U18748 ( .A(n17848), .B(n17847), .Z(n17833) );
  NANDN U18749 ( .A(n17818), .B(n17817), .Z(n17822) );
  OR U18750 ( .A(n17820), .B(n17819), .Z(n17821) );
  NAND U18751 ( .A(n17822), .B(n17821), .Z(n17834) );
  XNOR U18752 ( .A(n17833), .B(n17834), .Z(n17835) );
  XNOR U18753 ( .A(n17836), .B(n17835), .Z(n17828) );
  XOR U18754 ( .A(sreg[1757]), .B(n17828), .Z(n17829) );
  NAND U18755 ( .A(n17823), .B(sreg[1756]), .Z(n17827) );
  OR U18756 ( .A(n17825), .B(n17824), .Z(n17826) );
  NAND U18757 ( .A(n17827), .B(n17826), .Z(n17830) );
  XOR U18758 ( .A(n17829), .B(n17830), .Z(c[1757]) );
  OR U18759 ( .A(n17828), .B(sreg[1757]), .Z(n17832) );
  NANDN U18760 ( .A(n17830), .B(n17829), .Z(n17831) );
  NAND U18761 ( .A(n17832), .B(n17831), .Z(n17871) );
  NANDN U18762 ( .A(n17834), .B(n17833), .Z(n17838) );
  NAND U18763 ( .A(n17836), .B(n17835), .Z(n17837) );
  NAND U18764 ( .A(n17838), .B(n17837), .Z(n17854) );
  AND U18765 ( .A(b[2]), .B(a[736]), .Z(n17860) );
  AND U18766 ( .A(a[737]), .B(b[1]), .Z(n17858) );
  AND U18767 ( .A(a[735]), .B(b[3]), .Z(n17857) );
  XOR U18768 ( .A(n17858), .B(n17857), .Z(n17859) );
  XOR U18769 ( .A(n17860), .B(n17859), .Z(n17863) );
  NAND U18770 ( .A(b[0]), .B(a[738]), .Z(n17864) );
  XOR U18771 ( .A(n17863), .B(n17864), .Z(n17866) );
  OR U18772 ( .A(n17840), .B(n17839), .Z(n17844) );
  NANDN U18773 ( .A(n17842), .B(n17841), .Z(n17843) );
  NAND U18774 ( .A(n17844), .B(n17843), .Z(n17865) );
  XNOR U18775 ( .A(n17866), .B(n17865), .Z(n17851) );
  NANDN U18776 ( .A(n17846), .B(n17845), .Z(n17850) );
  OR U18777 ( .A(n17848), .B(n17847), .Z(n17849) );
  NAND U18778 ( .A(n17850), .B(n17849), .Z(n17852) );
  XNOR U18779 ( .A(n17851), .B(n17852), .Z(n17853) );
  XNOR U18780 ( .A(n17854), .B(n17853), .Z(n17869) );
  XNOR U18781 ( .A(n17869), .B(sreg[1758]), .Z(n17870) );
  XOR U18782 ( .A(n17871), .B(n17870), .Z(c[1758]) );
  NANDN U18783 ( .A(n17852), .B(n17851), .Z(n17856) );
  NAND U18784 ( .A(n17854), .B(n17853), .Z(n17855) );
  NAND U18785 ( .A(n17856), .B(n17855), .Z(n17877) );
  AND U18786 ( .A(b[2]), .B(a[737]), .Z(n17883) );
  AND U18787 ( .A(a[738]), .B(b[1]), .Z(n17881) );
  AND U18788 ( .A(a[736]), .B(b[3]), .Z(n17880) );
  XOR U18789 ( .A(n17881), .B(n17880), .Z(n17882) );
  XOR U18790 ( .A(n17883), .B(n17882), .Z(n17886) );
  NAND U18791 ( .A(b[0]), .B(a[739]), .Z(n17887) );
  XOR U18792 ( .A(n17886), .B(n17887), .Z(n17889) );
  OR U18793 ( .A(n17858), .B(n17857), .Z(n17862) );
  NANDN U18794 ( .A(n17860), .B(n17859), .Z(n17861) );
  NAND U18795 ( .A(n17862), .B(n17861), .Z(n17888) );
  XNOR U18796 ( .A(n17889), .B(n17888), .Z(n17874) );
  NANDN U18797 ( .A(n17864), .B(n17863), .Z(n17868) );
  OR U18798 ( .A(n17866), .B(n17865), .Z(n17867) );
  NAND U18799 ( .A(n17868), .B(n17867), .Z(n17875) );
  XNOR U18800 ( .A(n17874), .B(n17875), .Z(n17876) );
  XNOR U18801 ( .A(n17877), .B(n17876), .Z(n17892) );
  XNOR U18802 ( .A(n17892), .B(sreg[1759]), .Z(n17894) );
  NAND U18803 ( .A(n17869), .B(sreg[1758]), .Z(n17873) );
  OR U18804 ( .A(n17871), .B(n17870), .Z(n17872) );
  AND U18805 ( .A(n17873), .B(n17872), .Z(n17893) );
  XOR U18806 ( .A(n17894), .B(n17893), .Z(c[1759]) );
  NANDN U18807 ( .A(n17875), .B(n17874), .Z(n17879) );
  NAND U18808 ( .A(n17877), .B(n17876), .Z(n17878) );
  NAND U18809 ( .A(n17879), .B(n17878), .Z(n17903) );
  AND U18810 ( .A(b[2]), .B(a[738]), .Z(n17915) );
  AND U18811 ( .A(a[739]), .B(b[1]), .Z(n17913) );
  AND U18812 ( .A(a[737]), .B(b[3]), .Z(n17912) );
  XOR U18813 ( .A(n17913), .B(n17912), .Z(n17914) );
  XOR U18814 ( .A(n17915), .B(n17914), .Z(n17906) );
  NAND U18815 ( .A(b[0]), .B(a[740]), .Z(n17907) );
  XOR U18816 ( .A(n17906), .B(n17907), .Z(n17909) );
  OR U18817 ( .A(n17881), .B(n17880), .Z(n17885) );
  NANDN U18818 ( .A(n17883), .B(n17882), .Z(n17884) );
  NAND U18819 ( .A(n17885), .B(n17884), .Z(n17908) );
  XNOR U18820 ( .A(n17909), .B(n17908), .Z(n17900) );
  NANDN U18821 ( .A(n17887), .B(n17886), .Z(n17891) );
  OR U18822 ( .A(n17889), .B(n17888), .Z(n17890) );
  NAND U18823 ( .A(n17891), .B(n17890), .Z(n17901) );
  XNOR U18824 ( .A(n17900), .B(n17901), .Z(n17902) );
  XOR U18825 ( .A(n17903), .B(n17902), .Z(n17899) );
  NAND U18826 ( .A(n17892), .B(sreg[1759]), .Z(n17896) );
  OR U18827 ( .A(n17894), .B(n17893), .Z(n17895) );
  NAND U18828 ( .A(n17896), .B(n17895), .Z(n17898) );
  XNOR U18829 ( .A(sreg[1760]), .B(n17898), .Z(n17897) );
  XOR U18830 ( .A(n17899), .B(n17897), .Z(c[1760]) );
  NANDN U18831 ( .A(n17901), .B(n17900), .Z(n17905) );
  NAND U18832 ( .A(n17903), .B(n17902), .Z(n17904) );
  NAND U18833 ( .A(n17905), .B(n17904), .Z(n17933) );
  NANDN U18834 ( .A(n17907), .B(n17906), .Z(n17911) );
  OR U18835 ( .A(n17909), .B(n17908), .Z(n17910) );
  NAND U18836 ( .A(n17911), .B(n17910), .Z(n17930) );
  AND U18837 ( .A(b[2]), .B(a[739]), .Z(n17921) );
  AND U18838 ( .A(a[740]), .B(b[1]), .Z(n17919) );
  AND U18839 ( .A(a[738]), .B(b[3]), .Z(n17918) );
  XOR U18840 ( .A(n17919), .B(n17918), .Z(n17920) );
  XOR U18841 ( .A(n17921), .B(n17920), .Z(n17924) );
  NAND U18842 ( .A(b[0]), .B(a[741]), .Z(n17925) );
  XNOR U18843 ( .A(n17924), .B(n17925), .Z(n17926) );
  OR U18844 ( .A(n17913), .B(n17912), .Z(n17917) );
  NANDN U18845 ( .A(n17915), .B(n17914), .Z(n17916) );
  AND U18846 ( .A(n17917), .B(n17916), .Z(n17927) );
  XNOR U18847 ( .A(n17926), .B(n17927), .Z(n17931) );
  XNOR U18848 ( .A(n17930), .B(n17931), .Z(n17932) );
  XNOR U18849 ( .A(n17933), .B(n17932), .Z(n17936) );
  XNOR U18850 ( .A(sreg[1761]), .B(n17936), .Z(n17937) );
  XOR U18851 ( .A(n17938), .B(n17937), .Z(c[1761]) );
  AND U18852 ( .A(b[2]), .B(a[740]), .Z(n17950) );
  AND U18853 ( .A(a[741]), .B(b[1]), .Z(n17948) );
  AND U18854 ( .A(a[739]), .B(b[3]), .Z(n17947) );
  XOR U18855 ( .A(n17948), .B(n17947), .Z(n17949) );
  XOR U18856 ( .A(n17950), .B(n17949), .Z(n17953) );
  NAND U18857 ( .A(b[0]), .B(a[742]), .Z(n17954) );
  XOR U18858 ( .A(n17953), .B(n17954), .Z(n17956) );
  OR U18859 ( .A(n17919), .B(n17918), .Z(n17923) );
  NANDN U18860 ( .A(n17921), .B(n17920), .Z(n17922) );
  NAND U18861 ( .A(n17923), .B(n17922), .Z(n17955) );
  XNOR U18862 ( .A(n17956), .B(n17955), .Z(n17941) );
  NANDN U18863 ( .A(n17925), .B(n17924), .Z(n17929) );
  NAND U18864 ( .A(n17927), .B(n17926), .Z(n17928) );
  NAND U18865 ( .A(n17929), .B(n17928), .Z(n17942) );
  XNOR U18866 ( .A(n17941), .B(n17942), .Z(n17943) );
  NANDN U18867 ( .A(n17931), .B(n17930), .Z(n17935) );
  NANDN U18868 ( .A(n17933), .B(n17932), .Z(n17934) );
  NAND U18869 ( .A(n17935), .B(n17934), .Z(n17944) );
  XOR U18870 ( .A(n17943), .B(n17944), .Z(n17959) );
  XNOR U18871 ( .A(n17959), .B(sreg[1762]), .Z(n17961) );
  NAND U18872 ( .A(sreg[1761]), .B(n17936), .Z(n17940) );
  OR U18873 ( .A(n17938), .B(n17937), .Z(n17939) );
  AND U18874 ( .A(n17940), .B(n17939), .Z(n17960) );
  XOR U18875 ( .A(n17961), .B(n17960), .Z(c[1762]) );
  NANDN U18876 ( .A(n17942), .B(n17941), .Z(n17946) );
  NANDN U18877 ( .A(n17944), .B(n17943), .Z(n17945) );
  NAND U18878 ( .A(n17946), .B(n17945), .Z(n17982) );
  AND U18879 ( .A(b[2]), .B(a[741]), .Z(n17976) );
  AND U18880 ( .A(a[742]), .B(b[1]), .Z(n17974) );
  AND U18881 ( .A(a[740]), .B(b[3]), .Z(n17973) );
  XOR U18882 ( .A(n17974), .B(n17973), .Z(n17975) );
  XOR U18883 ( .A(n17976), .B(n17975), .Z(n17967) );
  NAND U18884 ( .A(b[0]), .B(a[743]), .Z(n17968) );
  XOR U18885 ( .A(n17967), .B(n17968), .Z(n17970) );
  OR U18886 ( .A(n17948), .B(n17947), .Z(n17952) );
  NANDN U18887 ( .A(n17950), .B(n17949), .Z(n17951) );
  NAND U18888 ( .A(n17952), .B(n17951), .Z(n17969) );
  XNOR U18889 ( .A(n17970), .B(n17969), .Z(n17979) );
  NANDN U18890 ( .A(n17954), .B(n17953), .Z(n17958) );
  OR U18891 ( .A(n17956), .B(n17955), .Z(n17957) );
  NAND U18892 ( .A(n17958), .B(n17957), .Z(n17980) );
  XNOR U18893 ( .A(n17979), .B(n17980), .Z(n17981) );
  XNOR U18894 ( .A(n17982), .B(n17981), .Z(n17966) );
  NAND U18895 ( .A(n17959), .B(sreg[1762]), .Z(n17963) );
  OR U18896 ( .A(n17961), .B(n17960), .Z(n17962) );
  AND U18897 ( .A(n17963), .B(n17962), .Z(n17965) );
  XNOR U18898 ( .A(n17965), .B(sreg[1763]), .Z(n17964) );
  XOR U18899 ( .A(n17966), .B(n17964), .Z(c[1763]) );
  NANDN U18900 ( .A(n17968), .B(n17967), .Z(n17972) );
  OR U18901 ( .A(n17970), .B(n17969), .Z(n17971) );
  NAND U18902 ( .A(n17972), .B(n17971), .Z(n17985) );
  AND U18903 ( .A(b[2]), .B(a[742]), .Z(n17994) );
  AND U18904 ( .A(a[743]), .B(b[1]), .Z(n17992) );
  AND U18905 ( .A(a[741]), .B(b[3]), .Z(n17991) );
  XOR U18906 ( .A(n17992), .B(n17991), .Z(n17993) );
  XOR U18907 ( .A(n17994), .B(n17993), .Z(n17997) );
  NAND U18908 ( .A(b[0]), .B(a[744]), .Z(n17998) );
  XNOR U18909 ( .A(n17997), .B(n17998), .Z(n17999) );
  OR U18910 ( .A(n17974), .B(n17973), .Z(n17978) );
  NANDN U18911 ( .A(n17976), .B(n17975), .Z(n17977) );
  AND U18912 ( .A(n17978), .B(n17977), .Z(n18000) );
  XNOR U18913 ( .A(n17999), .B(n18000), .Z(n17986) );
  XNOR U18914 ( .A(n17985), .B(n17986), .Z(n17987) );
  NANDN U18915 ( .A(n17980), .B(n17979), .Z(n17984) );
  NAND U18916 ( .A(n17982), .B(n17981), .Z(n17983) );
  AND U18917 ( .A(n17984), .B(n17983), .Z(n17988) );
  XNOR U18918 ( .A(n17987), .B(n17988), .Z(n18003) );
  XOR U18919 ( .A(n18003), .B(sreg[1764]), .Z(n18005) );
  XNOR U18920 ( .A(n18004), .B(n18005), .Z(c[1764]) );
  NANDN U18921 ( .A(n17986), .B(n17985), .Z(n17990) );
  NAND U18922 ( .A(n17988), .B(n17987), .Z(n17989) );
  NAND U18923 ( .A(n17990), .B(n17989), .Z(n18012) );
  AND U18924 ( .A(b[2]), .B(a[743]), .Z(n18018) );
  AND U18925 ( .A(a[744]), .B(b[1]), .Z(n18016) );
  AND U18926 ( .A(a[742]), .B(b[3]), .Z(n18015) );
  XOR U18927 ( .A(n18016), .B(n18015), .Z(n18017) );
  XOR U18928 ( .A(n18018), .B(n18017), .Z(n18021) );
  NAND U18929 ( .A(b[0]), .B(a[745]), .Z(n18022) );
  XOR U18930 ( .A(n18021), .B(n18022), .Z(n18024) );
  OR U18931 ( .A(n17992), .B(n17991), .Z(n17996) );
  NANDN U18932 ( .A(n17994), .B(n17993), .Z(n17995) );
  NAND U18933 ( .A(n17996), .B(n17995), .Z(n18023) );
  XNOR U18934 ( .A(n18024), .B(n18023), .Z(n18009) );
  NANDN U18935 ( .A(n17998), .B(n17997), .Z(n18002) );
  NAND U18936 ( .A(n18000), .B(n17999), .Z(n18001) );
  NAND U18937 ( .A(n18002), .B(n18001), .Z(n18010) );
  XNOR U18938 ( .A(n18009), .B(n18010), .Z(n18011) );
  XNOR U18939 ( .A(n18012), .B(n18011), .Z(n18028) );
  NANDN U18940 ( .A(n18003), .B(sreg[1764]), .Z(n18007) );
  NANDN U18941 ( .A(n18005), .B(n18004), .Z(n18006) );
  AND U18942 ( .A(n18007), .B(n18006), .Z(n18027) );
  XNOR U18943 ( .A(n18027), .B(sreg[1765]), .Z(n18008) );
  XNOR U18944 ( .A(n18028), .B(n18008), .Z(c[1765]) );
  NANDN U18945 ( .A(n18010), .B(n18009), .Z(n18014) );
  NANDN U18946 ( .A(n18012), .B(n18011), .Z(n18013) );
  NAND U18947 ( .A(n18014), .B(n18013), .Z(n18035) );
  AND U18948 ( .A(b[2]), .B(a[744]), .Z(n18041) );
  AND U18949 ( .A(a[745]), .B(b[1]), .Z(n18039) );
  AND U18950 ( .A(a[743]), .B(b[3]), .Z(n18038) );
  XOR U18951 ( .A(n18039), .B(n18038), .Z(n18040) );
  XOR U18952 ( .A(n18041), .B(n18040), .Z(n18044) );
  NAND U18953 ( .A(b[0]), .B(a[746]), .Z(n18045) );
  XOR U18954 ( .A(n18044), .B(n18045), .Z(n18047) );
  OR U18955 ( .A(n18016), .B(n18015), .Z(n18020) );
  NANDN U18956 ( .A(n18018), .B(n18017), .Z(n18019) );
  NAND U18957 ( .A(n18020), .B(n18019), .Z(n18046) );
  XNOR U18958 ( .A(n18047), .B(n18046), .Z(n18032) );
  NANDN U18959 ( .A(n18022), .B(n18021), .Z(n18026) );
  OR U18960 ( .A(n18024), .B(n18023), .Z(n18025) );
  NAND U18961 ( .A(n18026), .B(n18025), .Z(n18033) );
  XNOR U18962 ( .A(n18032), .B(n18033), .Z(n18034) );
  XNOR U18963 ( .A(n18035), .B(n18034), .Z(n18030) );
  XNOR U18964 ( .A(sreg[1766]), .B(n18031), .Z(n18029) );
  XNOR U18965 ( .A(n18030), .B(n18029), .Z(c[1766]) );
  NANDN U18966 ( .A(n18033), .B(n18032), .Z(n18037) );
  NAND U18967 ( .A(n18035), .B(n18034), .Z(n18036) );
  NAND U18968 ( .A(n18037), .B(n18036), .Z(n18058) );
  AND U18969 ( .A(b[2]), .B(a[745]), .Z(n18064) );
  AND U18970 ( .A(a[746]), .B(b[1]), .Z(n18062) );
  AND U18971 ( .A(a[744]), .B(b[3]), .Z(n18061) );
  XOR U18972 ( .A(n18062), .B(n18061), .Z(n18063) );
  XOR U18973 ( .A(n18064), .B(n18063), .Z(n18067) );
  NAND U18974 ( .A(b[0]), .B(a[747]), .Z(n18068) );
  XOR U18975 ( .A(n18067), .B(n18068), .Z(n18070) );
  OR U18976 ( .A(n18039), .B(n18038), .Z(n18043) );
  NANDN U18977 ( .A(n18041), .B(n18040), .Z(n18042) );
  NAND U18978 ( .A(n18043), .B(n18042), .Z(n18069) );
  XNOR U18979 ( .A(n18070), .B(n18069), .Z(n18055) );
  NANDN U18980 ( .A(n18045), .B(n18044), .Z(n18049) );
  OR U18981 ( .A(n18047), .B(n18046), .Z(n18048) );
  NAND U18982 ( .A(n18049), .B(n18048), .Z(n18056) );
  XNOR U18983 ( .A(n18055), .B(n18056), .Z(n18057) );
  XNOR U18984 ( .A(n18058), .B(n18057), .Z(n18050) );
  XNOR U18985 ( .A(n18050), .B(sreg[1767]), .Z(n18051) );
  XOR U18986 ( .A(n18052), .B(n18051), .Z(c[1767]) );
  NAND U18987 ( .A(n18050), .B(sreg[1767]), .Z(n18054) );
  OR U18988 ( .A(n18052), .B(n18051), .Z(n18053) );
  AND U18989 ( .A(n18054), .B(n18053), .Z(n18093) );
  NANDN U18990 ( .A(n18056), .B(n18055), .Z(n18060) );
  NAND U18991 ( .A(n18058), .B(n18057), .Z(n18059) );
  NAND U18992 ( .A(n18060), .B(n18059), .Z(n18077) );
  AND U18993 ( .A(b[2]), .B(a[746]), .Z(n18083) );
  AND U18994 ( .A(a[747]), .B(b[1]), .Z(n18081) );
  AND U18995 ( .A(a[745]), .B(b[3]), .Z(n18080) );
  XOR U18996 ( .A(n18081), .B(n18080), .Z(n18082) );
  XOR U18997 ( .A(n18083), .B(n18082), .Z(n18086) );
  NAND U18998 ( .A(b[0]), .B(a[748]), .Z(n18087) );
  XOR U18999 ( .A(n18086), .B(n18087), .Z(n18089) );
  OR U19000 ( .A(n18062), .B(n18061), .Z(n18066) );
  NANDN U19001 ( .A(n18064), .B(n18063), .Z(n18065) );
  NAND U19002 ( .A(n18066), .B(n18065), .Z(n18088) );
  XNOR U19003 ( .A(n18089), .B(n18088), .Z(n18074) );
  NANDN U19004 ( .A(n18068), .B(n18067), .Z(n18072) );
  OR U19005 ( .A(n18070), .B(n18069), .Z(n18071) );
  NAND U19006 ( .A(n18072), .B(n18071), .Z(n18075) );
  XNOR U19007 ( .A(n18074), .B(n18075), .Z(n18076) );
  XNOR U19008 ( .A(n18077), .B(n18076), .Z(n18092) );
  XNOR U19009 ( .A(sreg[1768]), .B(n18092), .Z(n18073) );
  XOR U19010 ( .A(n18093), .B(n18073), .Z(c[1768]) );
  NANDN U19011 ( .A(n18075), .B(n18074), .Z(n18079) );
  NAND U19012 ( .A(n18077), .B(n18076), .Z(n18078) );
  NAND U19013 ( .A(n18079), .B(n18078), .Z(n18100) );
  AND U19014 ( .A(b[2]), .B(a[747]), .Z(n18106) );
  AND U19015 ( .A(a[748]), .B(b[1]), .Z(n18104) );
  AND U19016 ( .A(a[746]), .B(b[3]), .Z(n18103) );
  XOR U19017 ( .A(n18104), .B(n18103), .Z(n18105) );
  XOR U19018 ( .A(n18106), .B(n18105), .Z(n18109) );
  NAND U19019 ( .A(b[0]), .B(a[749]), .Z(n18110) );
  XOR U19020 ( .A(n18109), .B(n18110), .Z(n18112) );
  OR U19021 ( .A(n18081), .B(n18080), .Z(n18085) );
  NANDN U19022 ( .A(n18083), .B(n18082), .Z(n18084) );
  NAND U19023 ( .A(n18085), .B(n18084), .Z(n18111) );
  XNOR U19024 ( .A(n18112), .B(n18111), .Z(n18097) );
  NANDN U19025 ( .A(n18087), .B(n18086), .Z(n18091) );
  OR U19026 ( .A(n18089), .B(n18088), .Z(n18090) );
  NAND U19027 ( .A(n18091), .B(n18090), .Z(n18098) );
  XNOR U19028 ( .A(n18097), .B(n18098), .Z(n18099) );
  XOR U19029 ( .A(n18100), .B(n18099), .Z(n18096) );
  XNOR U19030 ( .A(sreg[1769]), .B(n18095), .Z(n18094) );
  XOR U19031 ( .A(n18096), .B(n18094), .Z(c[1769]) );
  NANDN U19032 ( .A(n18098), .B(n18097), .Z(n18102) );
  NAND U19033 ( .A(n18100), .B(n18099), .Z(n18101) );
  NAND U19034 ( .A(n18102), .B(n18101), .Z(n18118) );
  AND U19035 ( .A(b[2]), .B(a[748]), .Z(n18124) );
  AND U19036 ( .A(a[749]), .B(b[1]), .Z(n18122) );
  AND U19037 ( .A(a[747]), .B(b[3]), .Z(n18121) );
  XOR U19038 ( .A(n18122), .B(n18121), .Z(n18123) );
  XOR U19039 ( .A(n18124), .B(n18123), .Z(n18127) );
  NAND U19040 ( .A(b[0]), .B(a[750]), .Z(n18128) );
  XOR U19041 ( .A(n18127), .B(n18128), .Z(n18130) );
  OR U19042 ( .A(n18104), .B(n18103), .Z(n18108) );
  NANDN U19043 ( .A(n18106), .B(n18105), .Z(n18107) );
  NAND U19044 ( .A(n18108), .B(n18107), .Z(n18129) );
  XNOR U19045 ( .A(n18130), .B(n18129), .Z(n18115) );
  NANDN U19046 ( .A(n18110), .B(n18109), .Z(n18114) );
  OR U19047 ( .A(n18112), .B(n18111), .Z(n18113) );
  NAND U19048 ( .A(n18114), .B(n18113), .Z(n18116) );
  XNOR U19049 ( .A(n18115), .B(n18116), .Z(n18117) );
  XNOR U19050 ( .A(n18118), .B(n18117), .Z(n18133) );
  XNOR U19051 ( .A(n18133), .B(sreg[1770]), .Z(n18134) );
  XOR U19052 ( .A(n18135), .B(n18134), .Z(c[1770]) );
  NANDN U19053 ( .A(n18116), .B(n18115), .Z(n18120) );
  NAND U19054 ( .A(n18118), .B(n18117), .Z(n18119) );
  NAND U19055 ( .A(n18120), .B(n18119), .Z(n18141) );
  AND U19056 ( .A(b[2]), .B(a[749]), .Z(n18147) );
  AND U19057 ( .A(a[750]), .B(b[1]), .Z(n18145) );
  AND U19058 ( .A(a[748]), .B(b[3]), .Z(n18144) );
  XOR U19059 ( .A(n18145), .B(n18144), .Z(n18146) );
  XOR U19060 ( .A(n18147), .B(n18146), .Z(n18150) );
  NAND U19061 ( .A(b[0]), .B(a[751]), .Z(n18151) );
  XOR U19062 ( .A(n18150), .B(n18151), .Z(n18153) );
  OR U19063 ( .A(n18122), .B(n18121), .Z(n18126) );
  NANDN U19064 ( .A(n18124), .B(n18123), .Z(n18125) );
  NAND U19065 ( .A(n18126), .B(n18125), .Z(n18152) );
  XNOR U19066 ( .A(n18153), .B(n18152), .Z(n18138) );
  NANDN U19067 ( .A(n18128), .B(n18127), .Z(n18132) );
  OR U19068 ( .A(n18130), .B(n18129), .Z(n18131) );
  NAND U19069 ( .A(n18132), .B(n18131), .Z(n18139) );
  XNOR U19070 ( .A(n18138), .B(n18139), .Z(n18140) );
  XNOR U19071 ( .A(n18141), .B(n18140), .Z(n18156) );
  XOR U19072 ( .A(sreg[1771]), .B(n18156), .Z(n18157) );
  NAND U19073 ( .A(n18133), .B(sreg[1770]), .Z(n18137) );
  OR U19074 ( .A(n18135), .B(n18134), .Z(n18136) );
  NAND U19075 ( .A(n18137), .B(n18136), .Z(n18158) );
  XOR U19076 ( .A(n18157), .B(n18158), .Z(c[1771]) );
  NANDN U19077 ( .A(n18139), .B(n18138), .Z(n18143) );
  NAND U19078 ( .A(n18141), .B(n18140), .Z(n18142) );
  NAND U19079 ( .A(n18143), .B(n18142), .Z(n18167) );
  AND U19080 ( .A(b[2]), .B(a[750]), .Z(n18173) );
  AND U19081 ( .A(a[751]), .B(b[1]), .Z(n18171) );
  AND U19082 ( .A(a[749]), .B(b[3]), .Z(n18170) );
  XOR U19083 ( .A(n18171), .B(n18170), .Z(n18172) );
  XOR U19084 ( .A(n18173), .B(n18172), .Z(n18176) );
  NAND U19085 ( .A(b[0]), .B(a[752]), .Z(n18177) );
  XOR U19086 ( .A(n18176), .B(n18177), .Z(n18179) );
  OR U19087 ( .A(n18145), .B(n18144), .Z(n18149) );
  NANDN U19088 ( .A(n18147), .B(n18146), .Z(n18148) );
  NAND U19089 ( .A(n18149), .B(n18148), .Z(n18178) );
  XNOR U19090 ( .A(n18179), .B(n18178), .Z(n18164) );
  NANDN U19091 ( .A(n18151), .B(n18150), .Z(n18155) );
  OR U19092 ( .A(n18153), .B(n18152), .Z(n18154) );
  NAND U19093 ( .A(n18155), .B(n18154), .Z(n18165) );
  XNOR U19094 ( .A(n18164), .B(n18165), .Z(n18166) );
  XOR U19095 ( .A(n18167), .B(n18166), .Z(n18163) );
  OR U19096 ( .A(n18156), .B(sreg[1771]), .Z(n18160) );
  NANDN U19097 ( .A(n18158), .B(n18157), .Z(n18159) );
  AND U19098 ( .A(n18160), .B(n18159), .Z(n18162) );
  XNOR U19099 ( .A(sreg[1772]), .B(n18162), .Z(n18161) );
  XOR U19100 ( .A(n18163), .B(n18161), .Z(c[1772]) );
  NANDN U19101 ( .A(n18165), .B(n18164), .Z(n18169) );
  NAND U19102 ( .A(n18167), .B(n18166), .Z(n18168) );
  NAND U19103 ( .A(n18169), .B(n18168), .Z(n18185) );
  AND U19104 ( .A(b[2]), .B(a[751]), .Z(n18191) );
  AND U19105 ( .A(a[752]), .B(b[1]), .Z(n18189) );
  AND U19106 ( .A(a[750]), .B(b[3]), .Z(n18188) );
  XOR U19107 ( .A(n18189), .B(n18188), .Z(n18190) );
  XOR U19108 ( .A(n18191), .B(n18190), .Z(n18194) );
  NAND U19109 ( .A(b[0]), .B(a[753]), .Z(n18195) );
  XOR U19110 ( .A(n18194), .B(n18195), .Z(n18197) );
  OR U19111 ( .A(n18171), .B(n18170), .Z(n18175) );
  NANDN U19112 ( .A(n18173), .B(n18172), .Z(n18174) );
  NAND U19113 ( .A(n18175), .B(n18174), .Z(n18196) );
  XNOR U19114 ( .A(n18197), .B(n18196), .Z(n18182) );
  NANDN U19115 ( .A(n18177), .B(n18176), .Z(n18181) );
  OR U19116 ( .A(n18179), .B(n18178), .Z(n18180) );
  NAND U19117 ( .A(n18181), .B(n18180), .Z(n18183) );
  XNOR U19118 ( .A(n18182), .B(n18183), .Z(n18184) );
  XNOR U19119 ( .A(n18185), .B(n18184), .Z(n18200) );
  XNOR U19120 ( .A(n18200), .B(sreg[1773]), .Z(n18201) );
  XOR U19121 ( .A(n18202), .B(n18201), .Z(c[1773]) );
  NANDN U19122 ( .A(n18183), .B(n18182), .Z(n18187) );
  NAND U19123 ( .A(n18185), .B(n18184), .Z(n18186) );
  NAND U19124 ( .A(n18187), .B(n18186), .Z(n18211) );
  AND U19125 ( .A(b[2]), .B(a[752]), .Z(n18217) );
  AND U19126 ( .A(a[753]), .B(b[1]), .Z(n18215) );
  AND U19127 ( .A(a[751]), .B(b[3]), .Z(n18214) );
  XOR U19128 ( .A(n18215), .B(n18214), .Z(n18216) );
  XOR U19129 ( .A(n18217), .B(n18216), .Z(n18220) );
  NAND U19130 ( .A(b[0]), .B(a[754]), .Z(n18221) );
  XOR U19131 ( .A(n18220), .B(n18221), .Z(n18223) );
  OR U19132 ( .A(n18189), .B(n18188), .Z(n18193) );
  NANDN U19133 ( .A(n18191), .B(n18190), .Z(n18192) );
  NAND U19134 ( .A(n18193), .B(n18192), .Z(n18222) );
  XNOR U19135 ( .A(n18223), .B(n18222), .Z(n18208) );
  NANDN U19136 ( .A(n18195), .B(n18194), .Z(n18199) );
  OR U19137 ( .A(n18197), .B(n18196), .Z(n18198) );
  NAND U19138 ( .A(n18199), .B(n18198), .Z(n18209) );
  XNOR U19139 ( .A(n18208), .B(n18209), .Z(n18210) );
  XNOR U19140 ( .A(n18211), .B(n18210), .Z(n18207) );
  NAND U19141 ( .A(n18200), .B(sreg[1773]), .Z(n18204) );
  OR U19142 ( .A(n18202), .B(n18201), .Z(n18203) );
  AND U19143 ( .A(n18204), .B(n18203), .Z(n18206) );
  XNOR U19144 ( .A(n18206), .B(sreg[1774]), .Z(n18205) );
  XOR U19145 ( .A(n18207), .B(n18205), .Z(c[1774]) );
  NANDN U19146 ( .A(n18209), .B(n18208), .Z(n18213) );
  NAND U19147 ( .A(n18211), .B(n18210), .Z(n18212) );
  NAND U19148 ( .A(n18213), .B(n18212), .Z(n18229) );
  AND U19149 ( .A(b[2]), .B(a[753]), .Z(n18235) );
  AND U19150 ( .A(a[754]), .B(b[1]), .Z(n18233) );
  AND U19151 ( .A(a[752]), .B(b[3]), .Z(n18232) );
  XOR U19152 ( .A(n18233), .B(n18232), .Z(n18234) );
  XOR U19153 ( .A(n18235), .B(n18234), .Z(n18238) );
  NAND U19154 ( .A(b[0]), .B(a[755]), .Z(n18239) );
  XOR U19155 ( .A(n18238), .B(n18239), .Z(n18241) );
  OR U19156 ( .A(n18215), .B(n18214), .Z(n18219) );
  NANDN U19157 ( .A(n18217), .B(n18216), .Z(n18218) );
  NAND U19158 ( .A(n18219), .B(n18218), .Z(n18240) );
  XNOR U19159 ( .A(n18241), .B(n18240), .Z(n18226) );
  NANDN U19160 ( .A(n18221), .B(n18220), .Z(n18225) );
  OR U19161 ( .A(n18223), .B(n18222), .Z(n18224) );
  NAND U19162 ( .A(n18225), .B(n18224), .Z(n18227) );
  XNOR U19163 ( .A(n18226), .B(n18227), .Z(n18228) );
  XNOR U19164 ( .A(n18229), .B(n18228), .Z(n18244) );
  XNOR U19165 ( .A(n18244), .B(sreg[1775]), .Z(n18246) );
  XNOR U19166 ( .A(n18245), .B(n18246), .Z(c[1775]) );
  NANDN U19167 ( .A(n18227), .B(n18226), .Z(n18231) );
  NAND U19168 ( .A(n18229), .B(n18228), .Z(n18230) );
  NAND U19169 ( .A(n18231), .B(n18230), .Z(n18255) );
  AND U19170 ( .A(b[2]), .B(a[754]), .Z(n18267) );
  AND U19171 ( .A(a[755]), .B(b[1]), .Z(n18265) );
  AND U19172 ( .A(a[753]), .B(b[3]), .Z(n18264) );
  XOR U19173 ( .A(n18265), .B(n18264), .Z(n18266) );
  XOR U19174 ( .A(n18267), .B(n18266), .Z(n18258) );
  NAND U19175 ( .A(b[0]), .B(a[756]), .Z(n18259) );
  XOR U19176 ( .A(n18258), .B(n18259), .Z(n18261) );
  OR U19177 ( .A(n18233), .B(n18232), .Z(n18237) );
  NANDN U19178 ( .A(n18235), .B(n18234), .Z(n18236) );
  NAND U19179 ( .A(n18237), .B(n18236), .Z(n18260) );
  XNOR U19180 ( .A(n18261), .B(n18260), .Z(n18252) );
  NANDN U19181 ( .A(n18239), .B(n18238), .Z(n18243) );
  OR U19182 ( .A(n18241), .B(n18240), .Z(n18242) );
  NAND U19183 ( .A(n18243), .B(n18242), .Z(n18253) );
  XNOR U19184 ( .A(n18252), .B(n18253), .Z(n18254) );
  XOR U19185 ( .A(n18255), .B(n18254), .Z(n18251) );
  NAND U19186 ( .A(n18244), .B(sreg[1775]), .Z(n18248) );
  NANDN U19187 ( .A(n18246), .B(n18245), .Z(n18247) );
  NAND U19188 ( .A(n18248), .B(n18247), .Z(n18250) );
  XNOR U19189 ( .A(sreg[1776]), .B(n18250), .Z(n18249) );
  XOR U19190 ( .A(n18251), .B(n18249), .Z(c[1776]) );
  NANDN U19191 ( .A(n18253), .B(n18252), .Z(n18257) );
  NAND U19192 ( .A(n18255), .B(n18254), .Z(n18256) );
  NAND U19193 ( .A(n18257), .B(n18256), .Z(n18285) );
  NANDN U19194 ( .A(n18259), .B(n18258), .Z(n18263) );
  OR U19195 ( .A(n18261), .B(n18260), .Z(n18262) );
  NAND U19196 ( .A(n18263), .B(n18262), .Z(n18282) );
  AND U19197 ( .A(b[2]), .B(a[755]), .Z(n18273) );
  AND U19198 ( .A(a[756]), .B(b[1]), .Z(n18271) );
  AND U19199 ( .A(a[754]), .B(b[3]), .Z(n18270) );
  XOR U19200 ( .A(n18271), .B(n18270), .Z(n18272) );
  XOR U19201 ( .A(n18273), .B(n18272), .Z(n18276) );
  NAND U19202 ( .A(b[0]), .B(a[757]), .Z(n18277) );
  XNOR U19203 ( .A(n18276), .B(n18277), .Z(n18278) );
  OR U19204 ( .A(n18265), .B(n18264), .Z(n18269) );
  NANDN U19205 ( .A(n18267), .B(n18266), .Z(n18268) );
  AND U19206 ( .A(n18269), .B(n18268), .Z(n18279) );
  XNOR U19207 ( .A(n18278), .B(n18279), .Z(n18283) );
  XNOR U19208 ( .A(n18282), .B(n18283), .Z(n18284) );
  XNOR U19209 ( .A(n18285), .B(n18284), .Z(n18288) );
  XNOR U19210 ( .A(sreg[1777]), .B(n18288), .Z(n18289) );
  XOR U19211 ( .A(n18290), .B(n18289), .Z(c[1777]) );
  AND U19212 ( .A(b[2]), .B(a[756]), .Z(n18305) );
  AND U19213 ( .A(a[757]), .B(b[1]), .Z(n18303) );
  AND U19214 ( .A(a[755]), .B(b[3]), .Z(n18302) );
  XOR U19215 ( .A(n18303), .B(n18302), .Z(n18304) );
  XOR U19216 ( .A(n18305), .B(n18304), .Z(n18308) );
  NAND U19217 ( .A(b[0]), .B(a[758]), .Z(n18309) );
  XOR U19218 ( .A(n18308), .B(n18309), .Z(n18311) );
  OR U19219 ( .A(n18271), .B(n18270), .Z(n18275) );
  NANDN U19220 ( .A(n18273), .B(n18272), .Z(n18274) );
  NAND U19221 ( .A(n18275), .B(n18274), .Z(n18310) );
  XNOR U19222 ( .A(n18311), .B(n18310), .Z(n18296) );
  NANDN U19223 ( .A(n18277), .B(n18276), .Z(n18281) );
  NAND U19224 ( .A(n18279), .B(n18278), .Z(n18280) );
  NAND U19225 ( .A(n18281), .B(n18280), .Z(n18297) );
  XNOR U19226 ( .A(n18296), .B(n18297), .Z(n18298) );
  NANDN U19227 ( .A(n18283), .B(n18282), .Z(n18287) );
  NANDN U19228 ( .A(n18285), .B(n18284), .Z(n18286) );
  NAND U19229 ( .A(n18287), .B(n18286), .Z(n18299) );
  XOR U19230 ( .A(n18298), .B(n18299), .Z(n18295) );
  NAND U19231 ( .A(sreg[1777]), .B(n18288), .Z(n18292) );
  OR U19232 ( .A(n18290), .B(n18289), .Z(n18291) );
  NAND U19233 ( .A(n18292), .B(n18291), .Z(n18294) );
  XNOR U19234 ( .A(sreg[1778]), .B(n18294), .Z(n18293) );
  XNOR U19235 ( .A(n18295), .B(n18293), .Z(c[1778]) );
  NANDN U19236 ( .A(n18297), .B(n18296), .Z(n18301) );
  NANDN U19237 ( .A(n18299), .B(n18298), .Z(n18300) );
  NAND U19238 ( .A(n18301), .B(n18300), .Z(n18329) );
  AND U19239 ( .A(b[2]), .B(a[757]), .Z(n18323) );
  AND U19240 ( .A(a[758]), .B(b[1]), .Z(n18321) );
  AND U19241 ( .A(a[756]), .B(b[3]), .Z(n18320) );
  XOR U19242 ( .A(n18321), .B(n18320), .Z(n18322) );
  XOR U19243 ( .A(n18323), .B(n18322), .Z(n18314) );
  NAND U19244 ( .A(b[0]), .B(a[759]), .Z(n18315) );
  XOR U19245 ( .A(n18314), .B(n18315), .Z(n18317) );
  OR U19246 ( .A(n18303), .B(n18302), .Z(n18307) );
  NANDN U19247 ( .A(n18305), .B(n18304), .Z(n18306) );
  NAND U19248 ( .A(n18307), .B(n18306), .Z(n18316) );
  XNOR U19249 ( .A(n18317), .B(n18316), .Z(n18326) );
  NANDN U19250 ( .A(n18309), .B(n18308), .Z(n18313) );
  OR U19251 ( .A(n18311), .B(n18310), .Z(n18312) );
  NAND U19252 ( .A(n18313), .B(n18312), .Z(n18327) );
  XNOR U19253 ( .A(n18326), .B(n18327), .Z(n18328) );
  XNOR U19254 ( .A(n18329), .B(n18328), .Z(n18332) );
  XNOR U19255 ( .A(n18332), .B(sreg[1779]), .Z(n18333) );
  XOR U19256 ( .A(n18334), .B(n18333), .Z(c[1779]) );
  NANDN U19257 ( .A(n18315), .B(n18314), .Z(n18319) );
  OR U19258 ( .A(n18317), .B(n18316), .Z(n18318) );
  NAND U19259 ( .A(n18319), .B(n18318), .Z(n18349) );
  AND U19260 ( .A(b[2]), .B(a[758]), .Z(n18340) );
  AND U19261 ( .A(a[759]), .B(b[1]), .Z(n18338) );
  AND U19262 ( .A(a[757]), .B(b[3]), .Z(n18337) );
  XOR U19263 ( .A(n18338), .B(n18337), .Z(n18339) );
  XOR U19264 ( .A(n18340), .B(n18339), .Z(n18343) );
  NAND U19265 ( .A(b[0]), .B(a[760]), .Z(n18344) );
  XNOR U19266 ( .A(n18343), .B(n18344), .Z(n18345) );
  OR U19267 ( .A(n18321), .B(n18320), .Z(n18325) );
  NANDN U19268 ( .A(n18323), .B(n18322), .Z(n18324) );
  AND U19269 ( .A(n18325), .B(n18324), .Z(n18346) );
  XNOR U19270 ( .A(n18345), .B(n18346), .Z(n18350) );
  XNOR U19271 ( .A(n18349), .B(n18350), .Z(n18351) );
  NANDN U19272 ( .A(n18327), .B(n18326), .Z(n18331) );
  NAND U19273 ( .A(n18329), .B(n18328), .Z(n18330) );
  AND U19274 ( .A(n18331), .B(n18330), .Z(n18352) );
  XOR U19275 ( .A(n18351), .B(n18352), .Z(n18355) );
  XNOR U19276 ( .A(sreg[1780]), .B(n18355), .Z(n18357) );
  NAND U19277 ( .A(n18332), .B(sreg[1779]), .Z(n18336) );
  OR U19278 ( .A(n18334), .B(n18333), .Z(n18335) );
  AND U19279 ( .A(n18336), .B(n18335), .Z(n18356) );
  XOR U19280 ( .A(n18357), .B(n18356), .Z(c[1780]) );
  AND U19281 ( .A(b[2]), .B(a[759]), .Z(n18369) );
  AND U19282 ( .A(a[760]), .B(b[1]), .Z(n18367) );
  AND U19283 ( .A(a[758]), .B(b[3]), .Z(n18366) );
  XOR U19284 ( .A(n18367), .B(n18366), .Z(n18368) );
  XOR U19285 ( .A(n18369), .B(n18368), .Z(n18372) );
  NAND U19286 ( .A(b[0]), .B(a[761]), .Z(n18373) );
  XOR U19287 ( .A(n18372), .B(n18373), .Z(n18375) );
  OR U19288 ( .A(n18338), .B(n18337), .Z(n18342) );
  NANDN U19289 ( .A(n18340), .B(n18339), .Z(n18341) );
  NAND U19290 ( .A(n18342), .B(n18341), .Z(n18374) );
  XNOR U19291 ( .A(n18375), .B(n18374), .Z(n18360) );
  NANDN U19292 ( .A(n18344), .B(n18343), .Z(n18348) );
  NAND U19293 ( .A(n18346), .B(n18345), .Z(n18347) );
  NAND U19294 ( .A(n18348), .B(n18347), .Z(n18361) );
  XNOR U19295 ( .A(n18360), .B(n18361), .Z(n18362) );
  NANDN U19296 ( .A(n18350), .B(n18349), .Z(n18354) );
  NAND U19297 ( .A(n18352), .B(n18351), .Z(n18353) );
  NAND U19298 ( .A(n18354), .B(n18353), .Z(n18363) );
  XOR U19299 ( .A(n18362), .B(n18363), .Z(n18378) );
  XNOR U19300 ( .A(n18378), .B(sreg[1781]), .Z(n18380) );
  NAND U19301 ( .A(sreg[1780]), .B(n18355), .Z(n18359) );
  OR U19302 ( .A(n18357), .B(n18356), .Z(n18358) );
  AND U19303 ( .A(n18359), .B(n18358), .Z(n18379) );
  XOR U19304 ( .A(n18380), .B(n18379), .Z(c[1781]) );
  NANDN U19305 ( .A(n18361), .B(n18360), .Z(n18365) );
  NANDN U19306 ( .A(n18363), .B(n18362), .Z(n18364) );
  NAND U19307 ( .A(n18365), .B(n18364), .Z(n18399) );
  AND U19308 ( .A(b[2]), .B(a[760]), .Z(n18393) );
  AND U19309 ( .A(a[761]), .B(b[1]), .Z(n18391) );
  AND U19310 ( .A(a[759]), .B(b[3]), .Z(n18390) );
  XOR U19311 ( .A(n18391), .B(n18390), .Z(n18392) );
  XOR U19312 ( .A(n18393), .B(n18392), .Z(n18384) );
  NAND U19313 ( .A(b[0]), .B(a[762]), .Z(n18385) );
  XOR U19314 ( .A(n18384), .B(n18385), .Z(n18387) );
  OR U19315 ( .A(n18367), .B(n18366), .Z(n18371) );
  NANDN U19316 ( .A(n18369), .B(n18368), .Z(n18370) );
  NAND U19317 ( .A(n18371), .B(n18370), .Z(n18386) );
  XNOR U19318 ( .A(n18387), .B(n18386), .Z(n18396) );
  NANDN U19319 ( .A(n18373), .B(n18372), .Z(n18377) );
  OR U19320 ( .A(n18375), .B(n18374), .Z(n18376) );
  NAND U19321 ( .A(n18377), .B(n18376), .Z(n18397) );
  XNOR U19322 ( .A(n18396), .B(n18397), .Z(n18398) );
  XOR U19323 ( .A(n18399), .B(n18398), .Z(n18403) );
  NAND U19324 ( .A(n18378), .B(sreg[1781]), .Z(n18382) );
  OR U19325 ( .A(n18380), .B(n18379), .Z(n18381) );
  NAND U19326 ( .A(n18382), .B(n18381), .Z(n18402) );
  XNOR U19327 ( .A(sreg[1782]), .B(n18402), .Z(n18383) );
  XOR U19328 ( .A(n18403), .B(n18383), .Z(c[1782]) );
  NANDN U19329 ( .A(n18385), .B(n18384), .Z(n18389) );
  OR U19330 ( .A(n18387), .B(n18386), .Z(n18388) );
  NAND U19331 ( .A(n18389), .B(n18388), .Z(n18405) );
  AND U19332 ( .A(b[2]), .B(a[761]), .Z(n18414) );
  AND U19333 ( .A(a[762]), .B(b[1]), .Z(n18412) );
  AND U19334 ( .A(a[760]), .B(b[3]), .Z(n18411) );
  XOR U19335 ( .A(n18412), .B(n18411), .Z(n18413) );
  XOR U19336 ( .A(n18414), .B(n18413), .Z(n18417) );
  NAND U19337 ( .A(b[0]), .B(a[763]), .Z(n18418) );
  XNOR U19338 ( .A(n18417), .B(n18418), .Z(n18419) );
  OR U19339 ( .A(n18391), .B(n18390), .Z(n18395) );
  NANDN U19340 ( .A(n18393), .B(n18392), .Z(n18394) );
  AND U19341 ( .A(n18395), .B(n18394), .Z(n18420) );
  XNOR U19342 ( .A(n18419), .B(n18420), .Z(n18406) );
  XNOR U19343 ( .A(n18405), .B(n18406), .Z(n18407) );
  NANDN U19344 ( .A(n18397), .B(n18396), .Z(n18401) );
  NAND U19345 ( .A(n18399), .B(n18398), .Z(n18400) );
  AND U19346 ( .A(n18401), .B(n18400), .Z(n18408) );
  XNOR U19347 ( .A(n18407), .B(n18408), .Z(n18424) );
  XNOR U19348 ( .A(sreg[1783]), .B(n18423), .Z(n18404) );
  XOR U19349 ( .A(n18424), .B(n18404), .Z(c[1783]) );
  NANDN U19350 ( .A(n18406), .B(n18405), .Z(n18410) );
  NAND U19351 ( .A(n18408), .B(n18407), .Z(n18409) );
  NAND U19352 ( .A(n18410), .B(n18409), .Z(n18429) );
  AND U19353 ( .A(b[2]), .B(a[762]), .Z(n18435) );
  AND U19354 ( .A(a[763]), .B(b[1]), .Z(n18433) );
  AND U19355 ( .A(a[761]), .B(b[3]), .Z(n18432) );
  XOR U19356 ( .A(n18433), .B(n18432), .Z(n18434) );
  XOR U19357 ( .A(n18435), .B(n18434), .Z(n18438) );
  NAND U19358 ( .A(b[0]), .B(a[764]), .Z(n18439) );
  XOR U19359 ( .A(n18438), .B(n18439), .Z(n18441) );
  OR U19360 ( .A(n18412), .B(n18411), .Z(n18416) );
  NANDN U19361 ( .A(n18414), .B(n18413), .Z(n18415) );
  NAND U19362 ( .A(n18416), .B(n18415), .Z(n18440) );
  XNOR U19363 ( .A(n18441), .B(n18440), .Z(n18426) );
  NANDN U19364 ( .A(n18418), .B(n18417), .Z(n18422) );
  NAND U19365 ( .A(n18420), .B(n18419), .Z(n18421) );
  NAND U19366 ( .A(n18422), .B(n18421), .Z(n18427) );
  XNOR U19367 ( .A(n18426), .B(n18427), .Z(n18428) );
  XOR U19368 ( .A(n18429), .B(n18428), .Z(n18445) );
  XNOR U19369 ( .A(sreg[1784]), .B(n18444), .Z(n18425) );
  XNOR U19370 ( .A(n18445), .B(n18425), .Z(c[1784]) );
  NANDN U19371 ( .A(n18427), .B(n18426), .Z(n18431) );
  NANDN U19372 ( .A(n18429), .B(n18428), .Z(n18430) );
  NAND U19373 ( .A(n18431), .B(n18430), .Z(n18464) );
  AND U19374 ( .A(b[2]), .B(a[763]), .Z(n18458) );
  AND U19375 ( .A(a[764]), .B(b[1]), .Z(n18456) );
  AND U19376 ( .A(a[762]), .B(b[3]), .Z(n18455) );
  XOR U19377 ( .A(n18456), .B(n18455), .Z(n18457) );
  XOR U19378 ( .A(n18458), .B(n18457), .Z(n18449) );
  NAND U19379 ( .A(b[0]), .B(a[765]), .Z(n18450) );
  XOR U19380 ( .A(n18449), .B(n18450), .Z(n18452) );
  OR U19381 ( .A(n18433), .B(n18432), .Z(n18437) );
  NANDN U19382 ( .A(n18435), .B(n18434), .Z(n18436) );
  NAND U19383 ( .A(n18437), .B(n18436), .Z(n18451) );
  XNOR U19384 ( .A(n18452), .B(n18451), .Z(n18461) );
  NANDN U19385 ( .A(n18439), .B(n18438), .Z(n18443) );
  OR U19386 ( .A(n18441), .B(n18440), .Z(n18442) );
  NAND U19387 ( .A(n18443), .B(n18442), .Z(n18462) );
  XNOR U19388 ( .A(n18461), .B(n18462), .Z(n18463) );
  XNOR U19389 ( .A(n18464), .B(n18463), .Z(n18448) );
  XOR U19390 ( .A(n18447), .B(sreg[1785]), .Z(n18446) );
  XOR U19391 ( .A(n18448), .B(n18446), .Z(c[1785]) );
  NANDN U19392 ( .A(n18450), .B(n18449), .Z(n18454) );
  OR U19393 ( .A(n18452), .B(n18451), .Z(n18453) );
  NAND U19394 ( .A(n18454), .B(n18453), .Z(n18467) );
  AND U19395 ( .A(b[2]), .B(a[764]), .Z(n18476) );
  AND U19396 ( .A(a[765]), .B(b[1]), .Z(n18474) );
  AND U19397 ( .A(a[763]), .B(b[3]), .Z(n18473) );
  XOR U19398 ( .A(n18474), .B(n18473), .Z(n18475) );
  XOR U19399 ( .A(n18476), .B(n18475), .Z(n18479) );
  NAND U19400 ( .A(b[0]), .B(a[766]), .Z(n18480) );
  XNOR U19401 ( .A(n18479), .B(n18480), .Z(n18481) );
  OR U19402 ( .A(n18456), .B(n18455), .Z(n18460) );
  NANDN U19403 ( .A(n18458), .B(n18457), .Z(n18459) );
  AND U19404 ( .A(n18460), .B(n18459), .Z(n18482) );
  XNOR U19405 ( .A(n18481), .B(n18482), .Z(n18468) );
  XNOR U19406 ( .A(n18467), .B(n18468), .Z(n18469) );
  NANDN U19407 ( .A(n18462), .B(n18461), .Z(n18466) );
  NAND U19408 ( .A(n18464), .B(n18463), .Z(n18465) );
  AND U19409 ( .A(n18466), .B(n18465), .Z(n18470) );
  XOR U19410 ( .A(n18469), .B(n18470), .Z(n18485) );
  XNOR U19411 ( .A(sreg[1786]), .B(n18485), .Z(n18487) );
  XNOR U19412 ( .A(n18486), .B(n18487), .Z(c[1786]) );
  NANDN U19413 ( .A(n18468), .B(n18467), .Z(n18472) );
  NAND U19414 ( .A(n18470), .B(n18469), .Z(n18471) );
  NAND U19415 ( .A(n18472), .B(n18471), .Z(n18496) );
  AND U19416 ( .A(b[2]), .B(a[765]), .Z(n18502) );
  AND U19417 ( .A(a[766]), .B(b[1]), .Z(n18500) );
  AND U19418 ( .A(a[764]), .B(b[3]), .Z(n18499) );
  XOR U19419 ( .A(n18500), .B(n18499), .Z(n18501) );
  XOR U19420 ( .A(n18502), .B(n18501), .Z(n18505) );
  NAND U19421 ( .A(b[0]), .B(a[767]), .Z(n18506) );
  XOR U19422 ( .A(n18505), .B(n18506), .Z(n18508) );
  OR U19423 ( .A(n18474), .B(n18473), .Z(n18478) );
  NANDN U19424 ( .A(n18476), .B(n18475), .Z(n18477) );
  NAND U19425 ( .A(n18478), .B(n18477), .Z(n18507) );
  XNOR U19426 ( .A(n18508), .B(n18507), .Z(n18493) );
  NANDN U19427 ( .A(n18480), .B(n18479), .Z(n18484) );
  NAND U19428 ( .A(n18482), .B(n18481), .Z(n18483) );
  NAND U19429 ( .A(n18484), .B(n18483), .Z(n18494) );
  XNOR U19430 ( .A(n18493), .B(n18494), .Z(n18495) );
  XNOR U19431 ( .A(n18496), .B(n18495), .Z(n18492) );
  NAND U19432 ( .A(sreg[1786]), .B(n18485), .Z(n18489) );
  NANDN U19433 ( .A(n18487), .B(n18486), .Z(n18488) );
  AND U19434 ( .A(n18489), .B(n18488), .Z(n18491) );
  XNOR U19435 ( .A(n18491), .B(sreg[1787]), .Z(n18490) );
  XNOR U19436 ( .A(n18492), .B(n18490), .Z(c[1787]) );
  NANDN U19437 ( .A(n18494), .B(n18493), .Z(n18498) );
  NANDN U19438 ( .A(n18496), .B(n18495), .Z(n18497) );
  NAND U19439 ( .A(n18498), .B(n18497), .Z(n18526) );
  AND U19440 ( .A(b[2]), .B(a[766]), .Z(n18520) );
  AND U19441 ( .A(a[767]), .B(b[1]), .Z(n18518) );
  AND U19442 ( .A(a[765]), .B(b[3]), .Z(n18517) );
  XOR U19443 ( .A(n18518), .B(n18517), .Z(n18519) );
  XOR U19444 ( .A(n18520), .B(n18519), .Z(n18511) );
  NAND U19445 ( .A(b[0]), .B(a[768]), .Z(n18512) );
  XOR U19446 ( .A(n18511), .B(n18512), .Z(n18514) );
  OR U19447 ( .A(n18500), .B(n18499), .Z(n18504) );
  NANDN U19448 ( .A(n18502), .B(n18501), .Z(n18503) );
  NAND U19449 ( .A(n18504), .B(n18503), .Z(n18513) );
  XNOR U19450 ( .A(n18514), .B(n18513), .Z(n18523) );
  NANDN U19451 ( .A(n18506), .B(n18505), .Z(n18510) );
  OR U19452 ( .A(n18508), .B(n18507), .Z(n18509) );
  NAND U19453 ( .A(n18510), .B(n18509), .Z(n18524) );
  XNOR U19454 ( .A(n18523), .B(n18524), .Z(n18525) );
  XNOR U19455 ( .A(n18526), .B(n18525), .Z(n18529) );
  XOR U19456 ( .A(sreg[1788]), .B(n18529), .Z(n18530) );
  XOR U19457 ( .A(n18531), .B(n18530), .Z(c[1788]) );
  NANDN U19458 ( .A(n18512), .B(n18511), .Z(n18516) );
  OR U19459 ( .A(n18514), .B(n18513), .Z(n18515) );
  NAND U19460 ( .A(n18516), .B(n18515), .Z(n18535) );
  AND U19461 ( .A(b[2]), .B(a[767]), .Z(n18544) );
  AND U19462 ( .A(a[768]), .B(b[1]), .Z(n18542) );
  AND U19463 ( .A(a[766]), .B(b[3]), .Z(n18541) );
  XOR U19464 ( .A(n18542), .B(n18541), .Z(n18543) );
  XOR U19465 ( .A(n18544), .B(n18543), .Z(n18547) );
  NAND U19466 ( .A(b[0]), .B(a[769]), .Z(n18548) );
  XNOR U19467 ( .A(n18547), .B(n18548), .Z(n18549) );
  OR U19468 ( .A(n18518), .B(n18517), .Z(n18522) );
  NANDN U19469 ( .A(n18520), .B(n18519), .Z(n18521) );
  AND U19470 ( .A(n18522), .B(n18521), .Z(n18550) );
  XNOR U19471 ( .A(n18549), .B(n18550), .Z(n18536) );
  XNOR U19472 ( .A(n18535), .B(n18536), .Z(n18537) );
  NANDN U19473 ( .A(n18524), .B(n18523), .Z(n18528) );
  NAND U19474 ( .A(n18526), .B(n18525), .Z(n18527) );
  AND U19475 ( .A(n18528), .B(n18527), .Z(n18538) );
  XNOR U19476 ( .A(n18537), .B(n18538), .Z(n18554) );
  OR U19477 ( .A(n18529), .B(sreg[1788]), .Z(n18533) );
  NANDN U19478 ( .A(n18531), .B(n18530), .Z(n18532) );
  AND U19479 ( .A(n18533), .B(n18532), .Z(n18553) );
  XNOR U19480 ( .A(sreg[1789]), .B(n18553), .Z(n18534) );
  XOR U19481 ( .A(n18554), .B(n18534), .Z(c[1789]) );
  NANDN U19482 ( .A(n18536), .B(n18535), .Z(n18540) );
  NAND U19483 ( .A(n18538), .B(n18537), .Z(n18539) );
  NAND U19484 ( .A(n18540), .B(n18539), .Z(n18559) );
  AND U19485 ( .A(b[2]), .B(a[768]), .Z(n18565) );
  AND U19486 ( .A(a[769]), .B(b[1]), .Z(n18563) );
  AND U19487 ( .A(a[767]), .B(b[3]), .Z(n18562) );
  XOR U19488 ( .A(n18563), .B(n18562), .Z(n18564) );
  XOR U19489 ( .A(n18565), .B(n18564), .Z(n18568) );
  NAND U19490 ( .A(b[0]), .B(a[770]), .Z(n18569) );
  XOR U19491 ( .A(n18568), .B(n18569), .Z(n18571) );
  OR U19492 ( .A(n18542), .B(n18541), .Z(n18546) );
  NANDN U19493 ( .A(n18544), .B(n18543), .Z(n18545) );
  NAND U19494 ( .A(n18546), .B(n18545), .Z(n18570) );
  XNOR U19495 ( .A(n18571), .B(n18570), .Z(n18556) );
  NANDN U19496 ( .A(n18548), .B(n18547), .Z(n18552) );
  NAND U19497 ( .A(n18550), .B(n18549), .Z(n18551) );
  NAND U19498 ( .A(n18552), .B(n18551), .Z(n18557) );
  XNOR U19499 ( .A(n18556), .B(n18557), .Z(n18558) );
  XNOR U19500 ( .A(n18559), .B(n18558), .Z(n18575) );
  XOR U19501 ( .A(n18574), .B(sreg[1790]), .Z(n18555) );
  XNOR U19502 ( .A(n18575), .B(n18555), .Z(c[1790]) );
  NANDN U19503 ( .A(n18557), .B(n18556), .Z(n18561) );
  NANDN U19504 ( .A(n18559), .B(n18558), .Z(n18560) );
  NAND U19505 ( .A(n18561), .B(n18560), .Z(n18580) );
  AND U19506 ( .A(b[2]), .B(a[769]), .Z(n18586) );
  AND U19507 ( .A(a[770]), .B(b[1]), .Z(n18584) );
  AND U19508 ( .A(a[768]), .B(b[3]), .Z(n18583) );
  XOR U19509 ( .A(n18584), .B(n18583), .Z(n18585) );
  XOR U19510 ( .A(n18586), .B(n18585), .Z(n18589) );
  NAND U19511 ( .A(b[0]), .B(a[771]), .Z(n18590) );
  XOR U19512 ( .A(n18589), .B(n18590), .Z(n18592) );
  OR U19513 ( .A(n18563), .B(n18562), .Z(n18567) );
  NANDN U19514 ( .A(n18565), .B(n18564), .Z(n18566) );
  NAND U19515 ( .A(n18567), .B(n18566), .Z(n18591) );
  XNOR U19516 ( .A(n18592), .B(n18591), .Z(n18577) );
  NANDN U19517 ( .A(n18569), .B(n18568), .Z(n18573) );
  OR U19518 ( .A(n18571), .B(n18570), .Z(n18572) );
  NAND U19519 ( .A(n18573), .B(n18572), .Z(n18578) );
  XNOR U19520 ( .A(n18577), .B(n18578), .Z(n18579) );
  XNOR U19521 ( .A(n18580), .B(n18579), .Z(n18596) );
  XNOR U19522 ( .A(sreg[1791]), .B(n18597), .Z(n18576) );
  XNOR U19523 ( .A(n18596), .B(n18576), .Z(c[1791]) );
  NANDN U19524 ( .A(n18578), .B(n18577), .Z(n18582) );
  NAND U19525 ( .A(n18580), .B(n18579), .Z(n18581) );
  AND U19526 ( .A(n18582), .B(n18581), .Z(n18603) );
  AND U19527 ( .A(b[2]), .B(a[770]), .Z(n18611) );
  AND U19528 ( .A(a[771]), .B(b[1]), .Z(n18609) );
  AND U19529 ( .A(a[769]), .B(b[3]), .Z(n18608) );
  XOR U19530 ( .A(n18609), .B(n18608), .Z(n18610) );
  XOR U19531 ( .A(n18611), .B(n18610), .Z(n18604) );
  NAND U19532 ( .A(b[0]), .B(a[772]), .Z(n18605) );
  XOR U19533 ( .A(n18604), .B(n18605), .Z(n18606) );
  OR U19534 ( .A(n18584), .B(n18583), .Z(n18588) );
  NANDN U19535 ( .A(n18586), .B(n18585), .Z(n18587) );
  AND U19536 ( .A(n18588), .B(n18587), .Z(n18607) );
  XOR U19537 ( .A(n18606), .B(n18607), .Z(n18601) );
  NANDN U19538 ( .A(n18590), .B(n18589), .Z(n18594) );
  OR U19539 ( .A(n18592), .B(n18591), .Z(n18593) );
  AND U19540 ( .A(n18594), .B(n18593), .Z(n18602) );
  XOR U19541 ( .A(n18601), .B(n18602), .Z(n18595) );
  XNOR U19542 ( .A(n18603), .B(n18595), .Z(n18600) );
  XNOR U19543 ( .A(sreg[1792]), .B(n18599), .Z(n18598) );
  XOR U19544 ( .A(n18600), .B(n18598), .Z(c[1792]) );
  AND U19545 ( .A(b[2]), .B(a[771]), .Z(n18622) );
  AND U19546 ( .A(a[772]), .B(b[1]), .Z(n18620) );
  AND U19547 ( .A(a[770]), .B(b[3]), .Z(n18619) );
  XOR U19548 ( .A(n18620), .B(n18619), .Z(n18621) );
  XOR U19549 ( .A(n18622), .B(n18621), .Z(n18625) );
  NAND U19550 ( .A(b[0]), .B(a[773]), .Z(n18626) );
  XNOR U19551 ( .A(n18625), .B(n18626), .Z(n18627) );
  OR U19552 ( .A(n18609), .B(n18608), .Z(n18613) );
  NANDN U19553 ( .A(n18611), .B(n18610), .Z(n18612) );
  AND U19554 ( .A(n18613), .B(n18612), .Z(n18628) );
  XNOR U19555 ( .A(n18627), .B(n18628), .Z(n18632) );
  XNOR U19556 ( .A(n18631), .B(n18632), .Z(n18633) );
  XNOR U19557 ( .A(n18634), .B(n18633), .Z(n18614) );
  XNOR U19558 ( .A(sreg[1793]), .B(n18614), .Z(n18615) );
  XOR U19559 ( .A(n18616), .B(n18615), .Z(c[1793]) );
  NAND U19560 ( .A(sreg[1793]), .B(n18614), .Z(n18618) );
  OR U19561 ( .A(n18616), .B(n18615), .Z(n18617) );
  NAND U19562 ( .A(n18618), .B(n18617), .Z(n18657) );
  AND U19563 ( .A(b[2]), .B(a[772]), .Z(n18646) );
  AND U19564 ( .A(a[773]), .B(b[1]), .Z(n18644) );
  AND U19565 ( .A(a[771]), .B(b[3]), .Z(n18643) );
  XOR U19566 ( .A(n18644), .B(n18643), .Z(n18645) );
  XOR U19567 ( .A(n18646), .B(n18645), .Z(n18649) );
  NAND U19568 ( .A(b[0]), .B(a[774]), .Z(n18650) );
  XOR U19569 ( .A(n18649), .B(n18650), .Z(n18652) );
  OR U19570 ( .A(n18620), .B(n18619), .Z(n18624) );
  NANDN U19571 ( .A(n18622), .B(n18621), .Z(n18623) );
  NAND U19572 ( .A(n18624), .B(n18623), .Z(n18651) );
  XNOR U19573 ( .A(n18652), .B(n18651), .Z(n18637) );
  NANDN U19574 ( .A(n18626), .B(n18625), .Z(n18630) );
  NAND U19575 ( .A(n18628), .B(n18627), .Z(n18629) );
  NAND U19576 ( .A(n18630), .B(n18629), .Z(n18638) );
  XNOR U19577 ( .A(n18637), .B(n18638), .Z(n18639) );
  NANDN U19578 ( .A(n18632), .B(n18631), .Z(n18636) );
  NANDN U19579 ( .A(n18634), .B(n18633), .Z(n18635) );
  AND U19580 ( .A(n18636), .B(n18635), .Z(n18640) );
  XNOR U19581 ( .A(n18639), .B(n18640), .Z(n18655) );
  XOR U19582 ( .A(sreg[1794]), .B(n18655), .Z(n18656) );
  XOR U19583 ( .A(n18657), .B(n18656), .Z(c[1794]) );
  NANDN U19584 ( .A(n18638), .B(n18637), .Z(n18642) );
  NAND U19585 ( .A(n18640), .B(n18639), .Z(n18641) );
  NAND U19586 ( .A(n18642), .B(n18641), .Z(n18678) );
  AND U19587 ( .A(b[2]), .B(a[773]), .Z(n18672) );
  AND U19588 ( .A(a[774]), .B(b[1]), .Z(n18670) );
  AND U19589 ( .A(a[772]), .B(b[3]), .Z(n18669) );
  XOR U19590 ( .A(n18670), .B(n18669), .Z(n18671) );
  XOR U19591 ( .A(n18672), .B(n18671), .Z(n18663) );
  NAND U19592 ( .A(b[0]), .B(a[775]), .Z(n18664) );
  XOR U19593 ( .A(n18663), .B(n18664), .Z(n18666) );
  OR U19594 ( .A(n18644), .B(n18643), .Z(n18648) );
  NANDN U19595 ( .A(n18646), .B(n18645), .Z(n18647) );
  NAND U19596 ( .A(n18648), .B(n18647), .Z(n18665) );
  XNOR U19597 ( .A(n18666), .B(n18665), .Z(n18675) );
  NANDN U19598 ( .A(n18650), .B(n18649), .Z(n18654) );
  OR U19599 ( .A(n18652), .B(n18651), .Z(n18653) );
  NAND U19600 ( .A(n18654), .B(n18653), .Z(n18676) );
  XNOR U19601 ( .A(n18675), .B(n18676), .Z(n18677) );
  XOR U19602 ( .A(n18678), .B(n18677), .Z(n18662) );
  OR U19603 ( .A(n18655), .B(sreg[1794]), .Z(n18659) );
  NANDN U19604 ( .A(n18657), .B(n18656), .Z(n18658) );
  AND U19605 ( .A(n18659), .B(n18658), .Z(n18661) );
  XNOR U19606 ( .A(sreg[1795]), .B(n18661), .Z(n18660) );
  XOR U19607 ( .A(n18662), .B(n18660), .Z(c[1795]) );
  NANDN U19608 ( .A(n18664), .B(n18663), .Z(n18668) );
  OR U19609 ( .A(n18666), .B(n18665), .Z(n18667) );
  NAND U19610 ( .A(n18668), .B(n18667), .Z(n18693) );
  AND U19611 ( .A(b[2]), .B(a[774]), .Z(n18684) );
  AND U19612 ( .A(a[775]), .B(b[1]), .Z(n18682) );
  AND U19613 ( .A(a[773]), .B(b[3]), .Z(n18681) );
  XOR U19614 ( .A(n18682), .B(n18681), .Z(n18683) );
  XOR U19615 ( .A(n18684), .B(n18683), .Z(n18687) );
  NAND U19616 ( .A(b[0]), .B(a[776]), .Z(n18688) );
  XNOR U19617 ( .A(n18687), .B(n18688), .Z(n18689) );
  OR U19618 ( .A(n18670), .B(n18669), .Z(n18674) );
  NANDN U19619 ( .A(n18672), .B(n18671), .Z(n18673) );
  AND U19620 ( .A(n18674), .B(n18673), .Z(n18690) );
  XNOR U19621 ( .A(n18689), .B(n18690), .Z(n18694) );
  XNOR U19622 ( .A(n18693), .B(n18694), .Z(n18695) );
  NANDN U19623 ( .A(n18676), .B(n18675), .Z(n18680) );
  NAND U19624 ( .A(n18678), .B(n18677), .Z(n18679) );
  AND U19625 ( .A(n18680), .B(n18679), .Z(n18696) );
  XOR U19626 ( .A(n18695), .B(n18696), .Z(n18699) );
  XNOR U19627 ( .A(sreg[1796]), .B(n18699), .Z(n18700) );
  XOR U19628 ( .A(n18701), .B(n18700), .Z(c[1796]) );
  AND U19629 ( .A(b[2]), .B(a[775]), .Z(n18713) );
  AND U19630 ( .A(a[776]), .B(b[1]), .Z(n18711) );
  AND U19631 ( .A(a[774]), .B(b[3]), .Z(n18710) );
  XOR U19632 ( .A(n18711), .B(n18710), .Z(n18712) );
  XOR U19633 ( .A(n18713), .B(n18712), .Z(n18716) );
  NAND U19634 ( .A(b[0]), .B(a[777]), .Z(n18717) );
  XOR U19635 ( .A(n18716), .B(n18717), .Z(n18719) );
  OR U19636 ( .A(n18682), .B(n18681), .Z(n18686) );
  NANDN U19637 ( .A(n18684), .B(n18683), .Z(n18685) );
  NAND U19638 ( .A(n18686), .B(n18685), .Z(n18718) );
  XNOR U19639 ( .A(n18719), .B(n18718), .Z(n18704) );
  NANDN U19640 ( .A(n18688), .B(n18687), .Z(n18692) );
  NAND U19641 ( .A(n18690), .B(n18689), .Z(n18691) );
  NAND U19642 ( .A(n18692), .B(n18691), .Z(n18705) );
  XNOR U19643 ( .A(n18704), .B(n18705), .Z(n18706) );
  NANDN U19644 ( .A(n18694), .B(n18693), .Z(n18698) );
  NAND U19645 ( .A(n18696), .B(n18695), .Z(n18697) );
  AND U19646 ( .A(n18698), .B(n18697), .Z(n18707) );
  XNOR U19647 ( .A(n18706), .B(n18707), .Z(n18722) );
  XOR U19648 ( .A(sreg[1797]), .B(n18722), .Z(n18723) );
  NAND U19649 ( .A(sreg[1796]), .B(n18699), .Z(n18703) );
  OR U19650 ( .A(n18701), .B(n18700), .Z(n18702) );
  NAND U19651 ( .A(n18703), .B(n18702), .Z(n18724) );
  XOR U19652 ( .A(n18723), .B(n18724), .Z(c[1797]) );
  NANDN U19653 ( .A(n18705), .B(n18704), .Z(n18709) );
  NAND U19654 ( .A(n18707), .B(n18706), .Z(n18708) );
  NAND U19655 ( .A(n18709), .B(n18708), .Z(n18731) );
  AND U19656 ( .A(b[2]), .B(a[776]), .Z(n18737) );
  AND U19657 ( .A(a[777]), .B(b[1]), .Z(n18735) );
  AND U19658 ( .A(a[775]), .B(b[3]), .Z(n18734) );
  XOR U19659 ( .A(n18735), .B(n18734), .Z(n18736) );
  XOR U19660 ( .A(n18737), .B(n18736), .Z(n18740) );
  NAND U19661 ( .A(b[0]), .B(a[778]), .Z(n18741) );
  XOR U19662 ( .A(n18740), .B(n18741), .Z(n18743) );
  OR U19663 ( .A(n18711), .B(n18710), .Z(n18715) );
  NANDN U19664 ( .A(n18713), .B(n18712), .Z(n18714) );
  NAND U19665 ( .A(n18715), .B(n18714), .Z(n18742) );
  XNOR U19666 ( .A(n18743), .B(n18742), .Z(n18728) );
  NANDN U19667 ( .A(n18717), .B(n18716), .Z(n18721) );
  OR U19668 ( .A(n18719), .B(n18718), .Z(n18720) );
  NAND U19669 ( .A(n18721), .B(n18720), .Z(n18729) );
  XNOR U19670 ( .A(n18728), .B(n18729), .Z(n18730) );
  XOR U19671 ( .A(n18731), .B(n18730), .Z(n18747) );
  OR U19672 ( .A(n18722), .B(sreg[1797]), .Z(n18726) );
  NANDN U19673 ( .A(n18724), .B(n18723), .Z(n18725) );
  AND U19674 ( .A(n18726), .B(n18725), .Z(n18746) );
  XNOR U19675 ( .A(sreg[1798]), .B(n18746), .Z(n18727) );
  XOR U19676 ( .A(n18747), .B(n18727), .Z(c[1798]) );
  NANDN U19677 ( .A(n18729), .B(n18728), .Z(n18733) );
  NAND U19678 ( .A(n18731), .B(n18730), .Z(n18732) );
  NAND U19679 ( .A(n18733), .B(n18732), .Z(n18754) );
  AND U19680 ( .A(b[2]), .B(a[777]), .Z(n18760) );
  AND U19681 ( .A(a[778]), .B(b[1]), .Z(n18758) );
  AND U19682 ( .A(a[776]), .B(b[3]), .Z(n18757) );
  XOR U19683 ( .A(n18758), .B(n18757), .Z(n18759) );
  XOR U19684 ( .A(n18760), .B(n18759), .Z(n18763) );
  NAND U19685 ( .A(b[0]), .B(a[779]), .Z(n18764) );
  XOR U19686 ( .A(n18763), .B(n18764), .Z(n18766) );
  OR U19687 ( .A(n18735), .B(n18734), .Z(n18739) );
  NANDN U19688 ( .A(n18737), .B(n18736), .Z(n18738) );
  NAND U19689 ( .A(n18739), .B(n18738), .Z(n18765) );
  XNOR U19690 ( .A(n18766), .B(n18765), .Z(n18751) );
  NANDN U19691 ( .A(n18741), .B(n18740), .Z(n18745) );
  OR U19692 ( .A(n18743), .B(n18742), .Z(n18744) );
  NAND U19693 ( .A(n18745), .B(n18744), .Z(n18752) );
  XNOR U19694 ( .A(n18751), .B(n18752), .Z(n18753) );
  XNOR U19695 ( .A(n18754), .B(n18753), .Z(n18750) );
  XOR U19696 ( .A(n18749), .B(sreg[1799]), .Z(n18748) );
  XOR U19697 ( .A(n18750), .B(n18748), .Z(c[1799]) );
  NANDN U19698 ( .A(n18752), .B(n18751), .Z(n18756) );
  NAND U19699 ( .A(n18754), .B(n18753), .Z(n18755) );
  NAND U19700 ( .A(n18756), .B(n18755), .Z(n18777) );
  AND U19701 ( .A(b[2]), .B(a[778]), .Z(n18783) );
  AND U19702 ( .A(a[779]), .B(b[1]), .Z(n18781) );
  AND U19703 ( .A(a[777]), .B(b[3]), .Z(n18780) );
  XOR U19704 ( .A(n18781), .B(n18780), .Z(n18782) );
  XOR U19705 ( .A(n18783), .B(n18782), .Z(n18786) );
  NAND U19706 ( .A(b[0]), .B(a[780]), .Z(n18787) );
  XOR U19707 ( .A(n18786), .B(n18787), .Z(n18789) );
  OR U19708 ( .A(n18758), .B(n18757), .Z(n18762) );
  NANDN U19709 ( .A(n18760), .B(n18759), .Z(n18761) );
  NAND U19710 ( .A(n18762), .B(n18761), .Z(n18788) );
  XNOR U19711 ( .A(n18789), .B(n18788), .Z(n18774) );
  NANDN U19712 ( .A(n18764), .B(n18763), .Z(n18768) );
  OR U19713 ( .A(n18766), .B(n18765), .Z(n18767) );
  NAND U19714 ( .A(n18768), .B(n18767), .Z(n18775) );
  XNOR U19715 ( .A(n18774), .B(n18775), .Z(n18776) );
  XNOR U19716 ( .A(n18777), .B(n18776), .Z(n18769) );
  XOR U19717 ( .A(sreg[1800]), .B(n18769), .Z(n18770) );
  XOR U19718 ( .A(n18771), .B(n18770), .Z(c[1800]) );
  OR U19719 ( .A(n18769), .B(sreg[1800]), .Z(n18773) );
  NANDN U19720 ( .A(n18771), .B(n18770), .Z(n18772) );
  AND U19721 ( .A(n18773), .B(n18772), .Z(n18793) );
  NANDN U19722 ( .A(n18775), .B(n18774), .Z(n18779) );
  NAND U19723 ( .A(n18777), .B(n18776), .Z(n18778) );
  NAND U19724 ( .A(n18779), .B(n18778), .Z(n18798) );
  AND U19725 ( .A(b[2]), .B(a[779]), .Z(n18804) );
  AND U19726 ( .A(a[780]), .B(b[1]), .Z(n18802) );
  AND U19727 ( .A(a[778]), .B(b[3]), .Z(n18801) );
  XOR U19728 ( .A(n18802), .B(n18801), .Z(n18803) );
  XOR U19729 ( .A(n18804), .B(n18803), .Z(n18807) );
  NAND U19730 ( .A(b[0]), .B(a[781]), .Z(n18808) );
  XOR U19731 ( .A(n18807), .B(n18808), .Z(n18810) );
  OR U19732 ( .A(n18781), .B(n18780), .Z(n18785) );
  NANDN U19733 ( .A(n18783), .B(n18782), .Z(n18784) );
  NAND U19734 ( .A(n18785), .B(n18784), .Z(n18809) );
  XNOR U19735 ( .A(n18810), .B(n18809), .Z(n18795) );
  NANDN U19736 ( .A(n18787), .B(n18786), .Z(n18791) );
  OR U19737 ( .A(n18789), .B(n18788), .Z(n18790) );
  NAND U19738 ( .A(n18791), .B(n18790), .Z(n18796) );
  XNOR U19739 ( .A(n18795), .B(n18796), .Z(n18797) );
  XNOR U19740 ( .A(n18798), .B(n18797), .Z(n18794) );
  XOR U19741 ( .A(sreg[1801]), .B(n18794), .Z(n18792) );
  XOR U19742 ( .A(n18793), .B(n18792), .Z(c[1801]) );
  NANDN U19743 ( .A(n18796), .B(n18795), .Z(n18800) );
  NAND U19744 ( .A(n18798), .B(n18797), .Z(n18799) );
  NAND U19745 ( .A(n18800), .B(n18799), .Z(n18816) );
  AND U19746 ( .A(b[2]), .B(a[780]), .Z(n18822) );
  AND U19747 ( .A(a[781]), .B(b[1]), .Z(n18820) );
  AND U19748 ( .A(a[779]), .B(b[3]), .Z(n18819) );
  XOR U19749 ( .A(n18820), .B(n18819), .Z(n18821) );
  XOR U19750 ( .A(n18822), .B(n18821), .Z(n18825) );
  NAND U19751 ( .A(b[0]), .B(a[782]), .Z(n18826) );
  XOR U19752 ( .A(n18825), .B(n18826), .Z(n18828) );
  OR U19753 ( .A(n18802), .B(n18801), .Z(n18806) );
  NANDN U19754 ( .A(n18804), .B(n18803), .Z(n18805) );
  NAND U19755 ( .A(n18806), .B(n18805), .Z(n18827) );
  XNOR U19756 ( .A(n18828), .B(n18827), .Z(n18813) );
  NANDN U19757 ( .A(n18808), .B(n18807), .Z(n18812) );
  OR U19758 ( .A(n18810), .B(n18809), .Z(n18811) );
  NAND U19759 ( .A(n18812), .B(n18811), .Z(n18814) );
  XNOR U19760 ( .A(n18813), .B(n18814), .Z(n18815) );
  XNOR U19761 ( .A(n18816), .B(n18815), .Z(n18831) );
  XNOR U19762 ( .A(n18831), .B(sreg[1802]), .Z(n18833) );
  XNOR U19763 ( .A(n18832), .B(n18833), .Z(c[1802]) );
  NANDN U19764 ( .A(n18814), .B(n18813), .Z(n18818) );
  NAND U19765 ( .A(n18816), .B(n18815), .Z(n18817) );
  NAND U19766 ( .A(n18818), .B(n18817), .Z(n18842) );
  AND U19767 ( .A(b[2]), .B(a[781]), .Z(n18848) );
  AND U19768 ( .A(a[782]), .B(b[1]), .Z(n18846) );
  AND U19769 ( .A(a[780]), .B(b[3]), .Z(n18845) );
  XOR U19770 ( .A(n18846), .B(n18845), .Z(n18847) );
  XOR U19771 ( .A(n18848), .B(n18847), .Z(n18851) );
  NAND U19772 ( .A(b[0]), .B(a[783]), .Z(n18852) );
  XOR U19773 ( .A(n18851), .B(n18852), .Z(n18854) );
  OR U19774 ( .A(n18820), .B(n18819), .Z(n18824) );
  NANDN U19775 ( .A(n18822), .B(n18821), .Z(n18823) );
  NAND U19776 ( .A(n18824), .B(n18823), .Z(n18853) );
  XNOR U19777 ( .A(n18854), .B(n18853), .Z(n18839) );
  NANDN U19778 ( .A(n18826), .B(n18825), .Z(n18830) );
  OR U19779 ( .A(n18828), .B(n18827), .Z(n18829) );
  NAND U19780 ( .A(n18830), .B(n18829), .Z(n18840) );
  XNOR U19781 ( .A(n18839), .B(n18840), .Z(n18841) );
  XNOR U19782 ( .A(n18842), .B(n18841), .Z(n18838) );
  NAND U19783 ( .A(n18831), .B(sreg[1802]), .Z(n18835) );
  NANDN U19784 ( .A(n18833), .B(n18832), .Z(n18834) );
  AND U19785 ( .A(n18835), .B(n18834), .Z(n18837) );
  XNOR U19786 ( .A(n18837), .B(sreg[1803]), .Z(n18836) );
  XOR U19787 ( .A(n18838), .B(n18836), .Z(c[1803]) );
  NANDN U19788 ( .A(n18840), .B(n18839), .Z(n18844) );
  NAND U19789 ( .A(n18842), .B(n18841), .Z(n18843) );
  NAND U19790 ( .A(n18844), .B(n18843), .Z(n18860) );
  AND U19791 ( .A(b[2]), .B(a[782]), .Z(n18866) );
  AND U19792 ( .A(a[783]), .B(b[1]), .Z(n18864) );
  AND U19793 ( .A(a[781]), .B(b[3]), .Z(n18863) );
  XOR U19794 ( .A(n18864), .B(n18863), .Z(n18865) );
  XOR U19795 ( .A(n18866), .B(n18865), .Z(n18869) );
  NAND U19796 ( .A(b[0]), .B(a[784]), .Z(n18870) );
  XOR U19797 ( .A(n18869), .B(n18870), .Z(n18872) );
  OR U19798 ( .A(n18846), .B(n18845), .Z(n18850) );
  NANDN U19799 ( .A(n18848), .B(n18847), .Z(n18849) );
  NAND U19800 ( .A(n18850), .B(n18849), .Z(n18871) );
  XNOR U19801 ( .A(n18872), .B(n18871), .Z(n18857) );
  NANDN U19802 ( .A(n18852), .B(n18851), .Z(n18856) );
  OR U19803 ( .A(n18854), .B(n18853), .Z(n18855) );
  NAND U19804 ( .A(n18856), .B(n18855), .Z(n18858) );
  XNOR U19805 ( .A(n18857), .B(n18858), .Z(n18859) );
  XNOR U19806 ( .A(n18860), .B(n18859), .Z(n18875) );
  XNOR U19807 ( .A(n18875), .B(sreg[1804]), .Z(n18877) );
  XNOR U19808 ( .A(n18876), .B(n18877), .Z(c[1804]) );
  NANDN U19809 ( .A(n18858), .B(n18857), .Z(n18862) );
  NAND U19810 ( .A(n18860), .B(n18859), .Z(n18861) );
  NAND U19811 ( .A(n18862), .B(n18861), .Z(n18883) );
  AND U19812 ( .A(b[2]), .B(a[783]), .Z(n18889) );
  AND U19813 ( .A(a[784]), .B(b[1]), .Z(n18887) );
  AND U19814 ( .A(a[782]), .B(b[3]), .Z(n18886) );
  XOR U19815 ( .A(n18887), .B(n18886), .Z(n18888) );
  XOR U19816 ( .A(n18889), .B(n18888), .Z(n18892) );
  NAND U19817 ( .A(b[0]), .B(a[785]), .Z(n18893) );
  XOR U19818 ( .A(n18892), .B(n18893), .Z(n18895) );
  OR U19819 ( .A(n18864), .B(n18863), .Z(n18868) );
  NANDN U19820 ( .A(n18866), .B(n18865), .Z(n18867) );
  NAND U19821 ( .A(n18868), .B(n18867), .Z(n18894) );
  XNOR U19822 ( .A(n18895), .B(n18894), .Z(n18880) );
  NANDN U19823 ( .A(n18870), .B(n18869), .Z(n18874) );
  OR U19824 ( .A(n18872), .B(n18871), .Z(n18873) );
  NAND U19825 ( .A(n18874), .B(n18873), .Z(n18881) );
  XNOR U19826 ( .A(n18880), .B(n18881), .Z(n18882) );
  XNOR U19827 ( .A(n18883), .B(n18882), .Z(n18898) );
  XNOR U19828 ( .A(n18898), .B(sreg[1805]), .Z(n18900) );
  NAND U19829 ( .A(n18875), .B(sreg[1804]), .Z(n18879) );
  NANDN U19830 ( .A(n18877), .B(n18876), .Z(n18878) );
  AND U19831 ( .A(n18879), .B(n18878), .Z(n18899) );
  XOR U19832 ( .A(n18900), .B(n18899), .Z(c[1805]) );
  NANDN U19833 ( .A(n18881), .B(n18880), .Z(n18885) );
  NAND U19834 ( .A(n18883), .B(n18882), .Z(n18884) );
  NAND U19835 ( .A(n18885), .B(n18884), .Z(n18909) );
  AND U19836 ( .A(b[2]), .B(a[784]), .Z(n18915) );
  AND U19837 ( .A(a[785]), .B(b[1]), .Z(n18913) );
  AND U19838 ( .A(a[783]), .B(b[3]), .Z(n18912) );
  XOR U19839 ( .A(n18913), .B(n18912), .Z(n18914) );
  XOR U19840 ( .A(n18915), .B(n18914), .Z(n18918) );
  NAND U19841 ( .A(b[0]), .B(a[786]), .Z(n18919) );
  XOR U19842 ( .A(n18918), .B(n18919), .Z(n18921) );
  OR U19843 ( .A(n18887), .B(n18886), .Z(n18891) );
  NANDN U19844 ( .A(n18889), .B(n18888), .Z(n18890) );
  NAND U19845 ( .A(n18891), .B(n18890), .Z(n18920) );
  XNOR U19846 ( .A(n18921), .B(n18920), .Z(n18906) );
  NANDN U19847 ( .A(n18893), .B(n18892), .Z(n18897) );
  OR U19848 ( .A(n18895), .B(n18894), .Z(n18896) );
  NAND U19849 ( .A(n18897), .B(n18896), .Z(n18907) );
  XNOR U19850 ( .A(n18906), .B(n18907), .Z(n18908) );
  XOR U19851 ( .A(n18909), .B(n18908), .Z(n18905) );
  NAND U19852 ( .A(n18898), .B(sreg[1805]), .Z(n18902) );
  OR U19853 ( .A(n18900), .B(n18899), .Z(n18901) );
  NAND U19854 ( .A(n18902), .B(n18901), .Z(n18904) );
  XNOR U19855 ( .A(sreg[1806]), .B(n18904), .Z(n18903) );
  XOR U19856 ( .A(n18905), .B(n18903), .Z(c[1806]) );
  NANDN U19857 ( .A(n18907), .B(n18906), .Z(n18911) );
  NAND U19858 ( .A(n18909), .B(n18908), .Z(n18910) );
  NAND U19859 ( .A(n18911), .B(n18910), .Z(n18927) );
  AND U19860 ( .A(b[2]), .B(a[785]), .Z(n18933) );
  AND U19861 ( .A(a[786]), .B(b[1]), .Z(n18931) );
  AND U19862 ( .A(a[784]), .B(b[3]), .Z(n18930) );
  XOR U19863 ( .A(n18931), .B(n18930), .Z(n18932) );
  XOR U19864 ( .A(n18933), .B(n18932), .Z(n18936) );
  NAND U19865 ( .A(b[0]), .B(a[787]), .Z(n18937) );
  XOR U19866 ( .A(n18936), .B(n18937), .Z(n18939) );
  OR U19867 ( .A(n18913), .B(n18912), .Z(n18917) );
  NANDN U19868 ( .A(n18915), .B(n18914), .Z(n18916) );
  NAND U19869 ( .A(n18917), .B(n18916), .Z(n18938) );
  XNOR U19870 ( .A(n18939), .B(n18938), .Z(n18924) );
  NANDN U19871 ( .A(n18919), .B(n18918), .Z(n18923) );
  OR U19872 ( .A(n18921), .B(n18920), .Z(n18922) );
  NAND U19873 ( .A(n18923), .B(n18922), .Z(n18925) );
  XNOR U19874 ( .A(n18924), .B(n18925), .Z(n18926) );
  XNOR U19875 ( .A(n18927), .B(n18926), .Z(n18942) );
  XNOR U19876 ( .A(n18942), .B(sreg[1807]), .Z(n18943) );
  XOR U19877 ( .A(n18944), .B(n18943), .Z(c[1807]) );
  NANDN U19878 ( .A(n18925), .B(n18924), .Z(n18929) );
  NAND U19879 ( .A(n18927), .B(n18926), .Z(n18928) );
  NAND U19880 ( .A(n18929), .B(n18928), .Z(n18950) );
  AND U19881 ( .A(b[2]), .B(a[786]), .Z(n18956) );
  AND U19882 ( .A(a[787]), .B(b[1]), .Z(n18954) );
  AND U19883 ( .A(a[785]), .B(b[3]), .Z(n18953) );
  XOR U19884 ( .A(n18954), .B(n18953), .Z(n18955) );
  XOR U19885 ( .A(n18956), .B(n18955), .Z(n18959) );
  NAND U19886 ( .A(b[0]), .B(a[788]), .Z(n18960) );
  XOR U19887 ( .A(n18959), .B(n18960), .Z(n18962) );
  OR U19888 ( .A(n18931), .B(n18930), .Z(n18935) );
  NANDN U19889 ( .A(n18933), .B(n18932), .Z(n18934) );
  NAND U19890 ( .A(n18935), .B(n18934), .Z(n18961) );
  XNOR U19891 ( .A(n18962), .B(n18961), .Z(n18947) );
  NANDN U19892 ( .A(n18937), .B(n18936), .Z(n18941) );
  OR U19893 ( .A(n18939), .B(n18938), .Z(n18940) );
  NAND U19894 ( .A(n18941), .B(n18940), .Z(n18948) );
  XNOR U19895 ( .A(n18947), .B(n18948), .Z(n18949) );
  XNOR U19896 ( .A(n18950), .B(n18949), .Z(n18965) );
  XOR U19897 ( .A(sreg[1808]), .B(n18965), .Z(n18966) );
  NAND U19898 ( .A(n18942), .B(sreg[1807]), .Z(n18946) );
  OR U19899 ( .A(n18944), .B(n18943), .Z(n18945) );
  NAND U19900 ( .A(n18946), .B(n18945), .Z(n18967) );
  XOR U19901 ( .A(n18966), .B(n18967), .Z(c[1808]) );
  NANDN U19902 ( .A(n18948), .B(n18947), .Z(n18952) );
  NAND U19903 ( .A(n18950), .B(n18949), .Z(n18951) );
  NAND U19904 ( .A(n18952), .B(n18951), .Z(n18974) );
  AND U19905 ( .A(b[2]), .B(a[787]), .Z(n18980) );
  AND U19906 ( .A(a[788]), .B(b[1]), .Z(n18978) );
  AND U19907 ( .A(a[786]), .B(b[3]), .Z(n18977) );
  XOR U19908 ( .A(n18978), .B(n18977), .Z(n18979) );
  XOR U19909 ( .A(n18980), .B(n18979), .Z(n18983) );
  NAND U19910 ( .A(b[0]), .B(a[789]), .Z(n18984) );
  XOR U19911 ( .A(n18983), .B(n18984), .Z(n18986) );
  OR U19912 ( .A(n18954), .B(n18953), .Z(n18958) );
  NANDN U19913 ( .A(n18956), .B(n18955), .Z(n18957) );
  NAND U19914 ( .A(n18958), .B(n18957), .Z(n18985) );
  XNOR U19915 ( .A(n18986), .B(n18985), .Z(n18971) );
  NANDN U19916 ( .A(n18960), .B(n18959), .Z(n18964) );
  OR U19917 ( .A(n18962), .B(n18961), .Z(n18963) );
  NAND U19918 ( .A(n18964), .B(n18963), .Z(n18972) );
  XNOR U19919 ( .A(n18971), .B(n18972), .Z(n18973) );
  XOR U19920 ( .A(n18974), .B(n18973), .Z(n18990) );
  OR U19921 ( .A(n18965), .B(sreg[1808]), .Z(n18969) );
  NANDN U19922 ( .A(n18967), .B(n18966), .Z(n18968) );
  AND U19923 ( .A(n18969), .B(n18968), .Z(n18989) );
  XNOR U19924 ( .A(sreg[1809]), .B(n18989), .Z(n18970) );
  XOR U19925 ( .A(n18990), .B(n18970), .Z(c[1809]) );
  NANDN U19926 ( .A(n18972), .B(n18971), .Z(n18976) );
  NAND U19927 ( .A(n18974), .B(n18973), .Z(n18975) );
  NAND U19928 ( .A(n18976), .B(n18975), .Z(n18995) );
  AND U19929 ( .A(b[2]), .B(a[788]), .Z(n19001) );
  AND U19930 ( .A(a[789]), .B(b[1]), .Z(n18999) );
  AND U19931 ( .A(a[787]), .B(b[3]), .Z(n18998) );
  XOR U19932 ( .A(n18999), .B(n18998), .Z(n19000) );
  XOR U19933 ( .A(n19001), .B(n19000), .Z(n19004) );
  NAND U19934 ( .A(b[0]), .B(a[790]), .Z(n19005) );
  XOR U19935 ( .A(n19004), .B(n19005), .Z(n19007) );
  OR U19936 ( .A(n18978), .B(n18977), .Z(n18982) );
  NANDN U19937 ( .A(n18980), .B(n18979), .Z(n18981) );
  NAND U19938 ( .A(n18982), .B(n18981), .Z(n19006) );
  XNOR U19939 ( .A(n19007), .B(n19006), .Z(n18992) );
  NANDN U19940 ( .A(n18984), .B(n18983), .Z(n18988) );
  OR U19941 ( .A(n18986), .B(n18985), .Z(n18987) );
  NAND U19942 ( .A(n18988), .B(n18987), .Z(n18993) );
  XNOR U19943 ( .A(n18992), .B(n18993), .Z(n18994) );
  XNOR U19944 ( .A(n18995), .B(n18994), .Z(n19011) );
  XOR U19945 ( .A(n19010), .B(sreg[1810]), .Z(n18991) );
  XOR U19946 ( .A(n19011), .B(n18991), .Z(c[1810]) );
  NANDN U19947 ( .A(n18993), .B(n18992), .Z(n18997) );
  NAND U19948 ( .A(n18995), .B(n18994), .Z(n18996) );
  NAND U19949 ( .A(n18997), .B(n18996), .Z(n19016) );
  AND U19950 ( .A(b[2]), .B(a[789]), .Z(n19022) );
  AND U19951 ( .A(a[790]), .B(b[1]), .Z(n19020) );
  AND U19952 ( .A(a[788]), .B(b[3]), .Z(n19019) );
  XOR U19953 ( .A(n19020), .B(n19019), .Z(n19021) );
  XOR U19954 ( .A(n19022), .B(n19021), .Z(n19025) );
  NAND U19955 ( .A(b[0]), .B(a[791]), .Z(n19026) );
  XOR U19956 ( .A(n19025), .B(n19026), .Z(n19028) );
  OR U19957 ( .A(n18999), .B(n18998), .Z(n19003) );
  NANDN U19958 ( .A(n19001), .B(n19000), .Z(n19002) );
  NAND U19959 ( .A(n19003), .B(n19002), .Z(n19027) );
  XNOR U19960 ( .A(n19028), .B(n19027), .Z(n19013) );
  NANDN U19961 ( .A(n19005), .B(n19004), .Z(n19009) );
  OR U19962 ( .A(n19007), .B(n19006), .Z(n19008) );
  NAND U19963 ( .A(n19009), .B(n19008), .Z(n19014) );
  XNOR U19964 ( .A(n19013), .B(n19014), .Z(n19015) );
  XOR U19965 ( .A(n19016), .B(n19015), .Z(n19032) );
  XOR U19966 ( .A(sreg[1811]), .B(n19031), .Z(n19012) );
  XOR U19967 ( .A(n19032), .B(n19012), .Z(c[1811]) );
  NANDN U19968 ( .A(n19014), .B(n19013), .Z(n19018) );
  NAND U19969 ( .A(n19016), .B(n19015), .Z(n19017) );
  NAND U19970 ( .A(n19018), .B(n19017), .Z(n19039) );
  AND U19971 ( .A(b[2]), .B(a[790]), .Z(n19045) );
  AND U19972 ( .A(a[791]), .B(b[1]), .Z(n19043) );
  AND U19973 ( .A(a[789]), .B(b[3]), .Z(n19042) );
  XOR U19974 ( .A(n19043), .B(n19042), .Z(n19044) );
  XOR U19975 ( .A(n19045), .B(n19044), .Z(n19048) );
  NAND U19976 ( .A(b[0]), .B(a[792]), .Z(n19049) );
  XOR U19977 ( .A(n19048), .B(n19049), .Z(n19051) );
  OR U19978 ( .A(n19020), .B(n19019), .Z(n19024) );
  NANDN U19979 ( .A(n19022), .B(n19021), .Z(n19023) );
  NAND U19980 ( .A(n19024), .B(n19023), .Z(n19050) );
  XNOR U19981 ( .A(n19051), .B(n19050), .Z(n19036) );
  NANDN U19982 ( .A(n19026), .B(n19025), .Z(n19030) );
  OR U19983 ( .A(n19028), .B(n19027), .Z(n19029) );
  NAND U19984 ( .A(n19030), .B(n19029), .Z(n19037) );
  XNOR U19985 ( .A(n19036), .B(n19037), .Z(n19038) );
  XNOR U19986 ( .A(n19039), .B(n19038), .Z(n19035) );
  XOR U19987 ( .A(n19034), .B(sreg[1812]), .Z(n19033) );
  XOR U19988 ( .A(n19035), .B(n19033), .Z(c[1812]) );
  NANDN U19989 ( .A(n19037), .B(n19036), .Z(n19041) );
  NAND U19990 ( .A(n19039), .B(n19038), .Z(n19040) );
  NAND U19991 ( .A(n19041), .B(n19040), .Z(n19057) );
  AND U19992 ( .A(b[2]), .B(a[791]), .Z(n19063) );
  AND U19993 ( .A(a[792]), .B(b[1]), .Z(n19061) );
  AND U19994 ( .A(a[790]), .B(b[3]), .Z(n19060) );
  XOR U19995 ( .A(n19061), .B(n19060), .Z(n19062) );
  XOR U19996 ( .A(n19063), .B(n19062), .Z(n19066) );
  NAND U19997 ( .A(b[0]), .B(a[793]), .Z(n19067) );
  XOR U19998 ( .A(n19066), .B(n19067), .Z(n19069) );
  OR U19999 ( .A(n19043), .B(n19042), .Z(n19047) );
  NANDN U20000 ( .A(n19045), .B(n19044), .Z(n19046) );
  NAND U20001 ( .A(n19047), .B(n19046), .Z(n19068) );
  XNOR U20002 ( .A(n19069), .B(n19068), .Z(n19054) );
  NANDN U20003 ( .A(n19049), .B(n19048), .Z(n19053) );
  OR U20004 ( .A(n19051), .B(n19050), .Z(n19052) );
  NAND U20005 ( .A(n19053), .B(n19052), .Z(n19055) );
  XNOR U20006 ( .A(n19054), .B(n19055), .Z(n19056) );
  XNOR U20007 ( .A(n19057), .B(n19056), .Z(n19072) );
  XNOR U20008 ( .A(n19072), .B(sreg[1813]), .Z(n19074) );
  XNOR U20009 ( .A(n19073), .B(n19074), .Z(c[1813]) );
  NANDN U20010 ( .A(n19055), .B(n19054), .Z(n19059) );
  NAND U20011 ( .A(n19057), .B(n19056), .Z(n19058) );
  NAND U20012 ( .A(n19059), .B(n19058), .Z(n19080) );
  AND U20013 ( .A(b[2]), .B(a[792]), .Z(n19086) );
  AND U20014 ( .A(a[793]), .B(b[1]), .Z(n19084) );
  AND U20015 ( .A(a[791]), .B(b[3]), .Z(n19083) );
  XOR U20016 ( .A(n19084), .B(n19083), .Z(n19085) );
  XOR U20017 ( .A(n19086), .B(n19085), .Z(n19089) );
  NAND U20018 ( .A(b[0]), .B(a[794]), .Z(n19090) );
  XOR U20019 ( .A(n19089), .B(n19090), .Z(n19092) );
  OR U20020 ( .A(n19061), .B(n19060), .Z(n19065) );
  NANDN U20021 ( .A(n19063), .B(n19062), .Z(n19064) );
  NAND U20022 ( .A(n19065), .B(n19064), .Z(n19091) );
  XNOR U20023 ( .A(n19092), .B(n19091), .Z(n19077) );
  NANDN U20024 ( .A(n19067), .B(n19066), .Z(n19071) );
  OR U20025 ( .A(n19069), .B(n19068), .Z(n19070) );
  NAND U20026 ( .A(n19071), .B(n19070), .Z(n19078) );
  XNOR U20027 ( .A(n19077), .B(n19078), .Z(n19079) );
  XNOR U20028 ( .A(n19080), .B(n19079), .Z(n19095) );
  XOR U20029 ( .A(sreg[1814]), .B(n19095), .Z(n19096) );
  NAND U20030 ( .A(n19072), .B(sreg[1813]), .Z(n19076) );
  NANDN U20031 ( .A(n19074), .B(n19073), .Z(n19075) );
  NAND U20032 ( .A(n19076), .B(n19075), .Z(n19097) );
  XOR U20033 ( .A(n19096), .B(n19097), .Z(c[1814]) );
  NANDN U20034 ( .A(n19078), .B(n19077), .Z(n19082) );
  NAND U20035 ( .A(n19080), .B(n19079), .Z(n19081) );
  NAND U20036 ( .A(n19082), .B(n19081), .Z(n19104) );
  AND U20037 ( .A(b[2]), .B(a[793]), .Z(n19110) );
  AND U20038 ( .A(a[794]), .B(b[1]), .Z(n19108) );
  AND U20039 ( .A(a[792]), .B(b[3]), .Z(n19107) );
  XOR U20040 ( .A(n19108), .B(n19107), .Z(n19109) );
  XOR U20041 ( .A(n19110), .B(n19109), .Z(n19113) );
  NAND U20042 ( .A(b[0]), .B(a[795]), .Z(n19114) );
  XOR U20043 ( .A(n19113), .B(n19114), .Z(n19116) );
  OR U20044 ( .A(n19084), .B(n19083), .Z(n19088) );
  NANDN U20045 ( .A(n19086), .B(n19085), .Z(n19087) );
  NAND U20046 ( .A(n19088), .B(n19087), .Z(n19115) );
  XNOR U20047 ( .A(n19116), .B(n19115), .Z(n19101) );
  NANDN U20048 ( .A(n19090), .B(n19089), .Z(n19094) );
  OR U20049 ( .A(n19092), .B(n19091), .Z(n19093) );
  NAND U20050 ( .A(n19094), .B(n19093), .Z(n19102) );
  XNOR U20051 ( .A(n19101), .B(n19102), .Z(n19103) );
  XOR U20052 ( .A(n19104), .B(n19103), .Z(n19120) );
  OR U20053 ( .A(n19095), .B(sreg[1814]), .Z(n19099) );
  NANDN U20054 ( .A(n19097), .B(n19096), .Z(n19098) );
  AND U20055 ( .A(n19099), .B(n19098), .Z(n19119) );
  XNOR U20056 ( .A(sreg[1815]), .B(n19119), .Z(n19100) );
  XOR U20057 ( .A(n19120), .B(n19100), .Z(c[1815]) );
  NANDN U20058 ( .A(n19102), .B(n19101), .Z(n19106) );
  NAND U20059 ( .A(n19104), .B(n19103), .Z(n19105) );
  NAND U20060 ( .A(n19106), .B(n19105), .Z(n19127) );
  AND U20061 ( .A(b[2]), .B(a[794]), .Z(n19133) );
  AND U20062 ( .A(a[795]), .B(b[1]), .Z(n19131) );
  AND U20063 ( .A(a[793]), .B(b[3]), .Z(n19130) );
  XOR U20064 ( .A(n19131), .B(n19130), .Z(n19132) );
  XOR U20065 ( .A(n19133), .B(n19132), .Z(n19136) );
  NAND U20066 ( .A(b[0]), .B(a[796]), .Z(n19137) );
  XOR U20067 ( .A(n19136), .B(n19137), .Z(n19139) );
  OR U20068 ( .A(n19108), .B(n19107), .Z(n19112) );
  NANDN U20069 ( .A(n19110), .B(n19109), .Z(n19111) );
  NAND U20070 ( .A(n19112), .B(n19111), .Z(n19138) );
  XNOR U20071 ( .A(n19139), .B(n19138), .Z(n19124) );
  NANDN U20072 ( .A(n19114), .B(n19113), .Z(n19118) );
  OR U20073 ( .A(n19116), .B(n19115), .Z(n19117) );
  NAND U20074 ( .A(n19118), .B(n19117), .Z(n19125) );
  XNOR U20075 ( .A(n19124), .B(n19125), .Z(n19126) );
  XOR U20076 ( .A(n19127), .B(n19126), .Z(n19123) );
  XNOR U20077 ( .A(sreg[1816]), .B(n19122), .Z(n19121) );
  XOR U20078 ( .A(n19123), .B(n19121), .Z(c[1816]) );
  NANDN U20079 ( .A(n19125), .B(n19124), .Z(n19129) );
  NAND U20080 ( .A(n19127), .B(n19126), .Z(n19128) );
  NAND U20081 ( .A(n19129), .B(n19128), .Z(n19150) );
  AND U20082 ( .A(b[2]), .B(a[795]), .Z(n19156) );
  AND U20083 ( .A(a[796]), .B(b[1]), .Z(n19154) );
  AND U20084 ( .A(a[794]), .B(b[3]), .Z(n19153) );
  XOR U20085 ( .A(n19154), .B(n19153), .Z(n19155) );
  XOR U20086 ( .A(n19156), .B(n19155), .Z(n19159) );
  NAND U20087 ( .A(b[0]), .B(a[797]), .Z(n19160) );
  XOR U20088 ( .A(n19159), .B(n19160), .Z(n19162) );
  OR U20089 ( .A(n19131), .B(n19130), .Z(n19135) );
  NANDN U20090 ( .A(n19133), .B(n19132), .Z(n19134) );
  NAND U20091 ( .A(n19135), .B(n19134), .Z(n19161) );
  XNOR U20092 ( .A(n19162), .B(n19161), .Z(n19147) );
  NANDN U20093 ( .A(n19137), .B(n19136), .Z(n19141) );
  OR U20094 ( .A(n19139), .B(n19138), .Z(n19140) );
  NAND U20095 ( .A(n19141), .B(n19140), .Z(n19148) );
  XNOR U20096 ( .A(n19147), .B(n19148), .Z(n19149) );
  XNOR U20097 ( .A(n19150), .B(n19149), .Z(n19142) );
  XOR U20098 ( .A(sreg[1817]), .B(n19142), .Z(n19144) );
  XNOR U20099 ( .A(n19143), .B(n19144), .Z(c[1817]) );
  OR U20100 ( .A(n19142), .B(sreg[1817]), .Z(n19146) );
  NAND U20101 ( .A(n19144), .B(n19143), .Z(n19145) );
  AND U20102 ( .A(n19146), .B(n19145), .Z(n19166) );
  NANDN U20103 ( .A(n19148), .B(n19147), .Z(n19152) );
  NAND U20104 ( .A(n19150), .B(n19149), .Z(n19151) );
  NAND U20105 ( .A(n19152), .B(n19151), .Z(n19171) );
  AND U20106 ( .A(b[2]), .B(a[796]), .Z(n19177) );
  AND U20107 ( .A(a[797]), .B(b[1]), .Z(n19175) );
  AND U20108 ( .A(a[795]), .B(b[3]), .Z(n19174) );
  XOR U20109 ( .A(n19175), .B(n19174), .Z(n19176) );
  XOR U20110 ( .A(n19177), .B(n19176), .Z(n19180) );
  NAND U20111 ( .A(b[0]), .B(a[798]), .Z(n19181) );
  XOR U20112 ( .A(n19180), .B(n19181), .Z(n19183) );
  OR U20113 ( .A(n19154), .B(n19153), .Z(n19158) );
  NANDN U20114 ( .A(n19156), .B(n19155), .Z(n19157) );
  NAND U20115 ( .A(n19158), .B(n19157), .Z(n19182) );
  XNOR U20116 ( .A(n19183), .B(n19182), .Z(n19168) );
  NANDN U20117 ( .A(n19160), .B(n19159), .Z(n19164) );
  OR U20118 ( .A(n19162), .B(n19161), .Z(n19163) );
  NAND U20119 ( .A(n19164), .B(n19163), .Z(n19169) );
  XNOR U20120 ( .A(n19168), .B(n19169), .Z(n19170) );
  XNOR U20121 ( .A(n19171), .B(n19170), .Z(n19167) );
  XOR U20122 ( .A(sreg[1818]), .B(n19167), .Z(n19165) );
  XOR U20123 ( .A(n19166), .B(n19165), .Z(c[1818]) );
  NANDN U20124 ( .A(n19169), .B(n19168), .Z(n19173) );
  NAND U20125 ( .A(n19171), .B(n19170), .Z(n19172) );
  NAND U20126 ( .A(n19173), .B(n19172), .Z(n19189) );
  AND U20127 ( .A(b[2]), .B(a[797]), .Z(n19195) );
  AND U20128 ( .A(a[798]), .B(b[1]), .Z(n19193) );
  AND U20129 ( .A(a[796]), .B(b[3]), .Z(n19192) );
  XOR U20130 ( .A(n19193), .B(n19192), .Z(n19194) );
  XOR U20131 ( .A(n19195), .B(n19194), .Z(n19198) );
  NAND U20132 ( .A(b[0]), .B(a[799]), .Z(n19199) );
  XOR U20133 ( .A(n19198), .B(n19199), .Z(n19201) );
  OR U20134 ( .A(n19175), .B(n19174), .Z(n19179) );
  NANDN U20135 ( .A(n19177), .B(n19176), .Z(n19178) );
  NAND U20136 ( .A(n19179), .B(n19178), .Z(n19200) );
  XNOR U20137 ( .A(n19201), .B(n19200), .Z(n19186) );
  NANDN U20138 ( .A(n19181), .B(n19180), .Z(n19185) );
  OR U20139 ( .A(n19183), .B(n19182), .Z(n19184) );
  NAND U20140 ( .A(n19185), .B(n19184), .Z(n19187) );
  XNOR U20141 ( .A(n19186), .B(n19187), .Z(n19188) );
  XNOR U20142 ( .A(n19189), .B(n19188), .Z(n19204) );
  XNOR U20143 ( .A(n19204), .B(sreg[1819]), .Z(n19206) );
  XNOR U20144 ( .A(n19205), .B(n19206), .Z(c[1819]) );
  NANDN U20145 ( .A(n19187), .B(n19186), .Z(n19191) );
  NAND U20146 ( .A(n19189), .B(n19188), .Z(n19190) );
  NAND U20147 ( .A(n19191), .B(n19190), .Z(n19212) );
  AND U20148 ( .A(b[2]), .B(a[798]), .Z(n19224) );
  AND U20149 ( .A(a[799]), .B(b[1]), .Z(n19222) );
  AND U20150 ( .A(a[797]), .B(b[3]), .Z(n19221) );
  XOR U20151 ( .A(n19222), .B(n19221), .Z(n19223) );
  XOR U20152 ( .A(n19224), .B(n19223), .Z(n19215) );
  NAND U20153 ( .A(b[0]), .B(a[800]), .Z(n19216) );
  XOR U20154 ( .A(n19215), .B(n19216), .Z(n19218) );
  OR U20155 ( .A(n19193), .B(n19192), .Z(n19197) );
  NANDN U20156 ( .A(n19195), .B(n19194), .Z(n19196) );
  NAND U20157 ( .A(n19197), .B(n19196), .Z(n19217) );
  XNOR U20158 ( .A(n19218), .B(n19217), .Z(n19209) );
  NANDN U20159 ( .A(n19199), .B(n19198), .Z(n19203) );
  OR U20160 ( .A(n19201), .B(n19200), .Z(n19202) );
  NAND U20161 ( .A(n19203), .B(n19202), .Z(n19210) );
  XNOR U20162 ( .A(n19209), .B(n19210), .Z(n19211) );
  XNOR U20163 ( .A(n19212), .B(n19211), .Z(n19228) );
  XOR U20164 ( .A(sreg[1820]), .B(n19228), .Z(n19229) );
  NAND U20165 ( .A(n19204), .B(sreg[1819]), .Z(n19208) );
  NANDN U20166 ( .A(n19206), .B(n19205), .Z(n19207) );
  NAND U20167 ( .A(n19208), .B(n19207), .Z(n19230) );
  XOR U20168 ( .A(n19229), .B(n19230), .Z(c[1820]) );
  NANDN U20169 ( .A(n19210), .B(n19209), .Z(n19214) );
  NAND U20170 ( .A(n19212), .B(n19211), .Z(n19213) );
  NAND U20171 ( .A(n19214), .B(n19213), .Z(n19238) );
  NANDN U20172 ( .A(n19216), .B(n19215), .Z(n19220) );
  OR U20173 ( .A(n19218), .B(n19217), .Z(n19219) );
  AND U20174 ( .A(n19220), .B(n19219), .Z(n19237) );
  AND U20175 ( .A(b[2]), .B(a[799]), .Z(n19248) );
  AND U20176 ( .A(a[800]), .B(b[1]), .Z(n19246) );
  AND U20177 ( .A(a[798]), .B(b[3]), .Z(n19245) );
  XOR U20178 ( .A(n19246), .B(n19245), .Z(n19247) );
  XOR U20179 ( .A(n19248), .B(n19247), .Z(n19239) );
  NAND U20180 ( .A(b[0]), .B(a[801]), .Z(n19240) );
  XOR U20181 ( .A(n19239), .B(n19240), .Z(n19242) );
  OR U20182 ( .A(n19222), .B(n19221), .Z(n19226) );
  NANDN U20183 ( .A(n19224), .B(n19223), .Z(n19225) );
  NAND U20184 ( .A(n19226), .B(n19225), .Z(n19241) );
  XOR U20185 ( .A(n19242), .B(n19241), .Z(n19236) );
  XNOR U20186 ( .A(n19237), .B(n19236), .Z(n19227) );
  XNOR U20187 ( .A(n19238), .B(n19227), .Z(n19235) );
  OR U20188 ( .A(n19228), .B(sreg[1820]), .Z(n19232) );
  NANDN U20189 ( .A(n19230), .B(n19229), .Z(n19231) );
  AND U20190 ( .A(n19232), .B(n19231), .Z(n19234) );
  XOR U20191 ( .A(sreg[1821]), .B(n19234), .Z(n19233) );
  XOR U20192 ( .A(n19235), .B(n19233), .Z(c[1821]) );
  NANDN U20193 ( .A(n19240), .B(n19239), .Z(n19244) );
  OR U20194 ( .A(n19242), .B(n19241), .Z(n19243) );
  AND U20195 ( .A(n19244), .B(n19243), .Z(n19253) );
  AND U20196 ( .A(b[2]), .B(a[800]), .Z(n19258) );
  AND U20197 ( .A(a[801]), .B(b[1]), .Z(n19256) );
  AND U20198 ( .A(a[799]), .B(b[3]), .Z(n19255) );
  XOR U20199 ( .A(n19256), .B(n19255), .Z(n19257) );
  XOR U20200 ( .A(n19258), .B(n19257), .Z(n19261) );
  NAND U20201 ( .A(b[0]), .B(a[802]), .Z(n19262) );
  XOR U20202 ( .A(n19261), .B(n19262), .Z(n19264) );
  OR U20203 ( .A(n19246), .B(n19245), .Z(n19250) );
  NANDN U20204 ( .A(n19248), .B(n19247), .Z(n19249) );
  NAND U20205 ( .A(n19250), .B(n19249), .Z(n19263) );
  XOR U20206 ( .A(n19264), .B(n19263), .Z(n19252) );
  XNOR U20207 ( .A(n19253), .B(n19252), .Z(n19251) );
  XOR U20208 ( .A(n19254), .B(n19251), .Z(n19267) );
  XNOR U20209 ( .A(n19267), .B(sreg[1822]), .Z(n19269) );
  XNOR U20210 ( .A(n19268), .B(n19269), .Z(c[1822]) );
  AND U20211 ( .A(b[2]), .B(a[801]), .Z(n19284) );
  AND U20212 ( .A(a[802]), .B(b[1]), .Z(n19282) );
  AND U20213 ( .A(a[800]), .B(b[3]), .Z(n19281) );
  XOR U20214 ( .A(n19282), .B(n19281), .Z(n19283) );
  XOR U20215 ( .A(n19284), .B(n19283), .Z(n19287) );
  NAND U20216 ( .A(b[0]), .B(a[803]), .Z(n19288) );
  XOR U20217 ( .A(n19287), .B(n19288), .Z(n19290) );
  OR U20218 ( .A(n19256), .B(n19255), .Z(n19260) );
  NANDN U20219 ( .A(n19258), .B(n19257), .Z(n19259) );
  NAND U20220 ( .A(n19260), .B(n19259), .Z(n19289) );
  XNOR U20221 ( .A(n19290), .B(n19289), .Z(n19275) );
  NANDN U20222 ( .A(n19262), .B(n19261), .Z(n19266) );
  OR U20223 ( .A(n19264), .B(n19263), .Z(n19265) );
  NAND U20224 ( .A(n19266), .B(n19265), .Z(n19276) );
  XNOR U20225 ( .A(n19275), .B(n19276), .Z(n19277) );
  XOR U20226 ( .A(n19278), .B(n19277), .Z(n19274) );
  NAND U20227 ( .A(n19267), .B(sreg[1822]), .Z(n19271) );
  NANDN U20228 ( .A(n19269), .B(n19268), .Z(n19270) );
  NAND U20229 ( .A(n19271), .B(n19270), .Z(n19273) );
  XNOR U20230 ( .A(sreg[1823]), .B(n19273), .Z(n19272) );
  XNOR U20231 ( .A(n19274), .B(n19272), .Z(c[1823]) );
  NANDN U20232 ( .A(n19276), .B(n19275), .Z(n19280) );
  NANDN U20233 ( .A(n19278), .B(n19277), .Z(n19279) );
  AND U20234 ( .A(n19280), .B(n19279), .Z(n19296) );
  AND U20235 ( .A(b[2]), .B(a[802]), .Z(n19300) );
  AND U20236 ( .A(a[803]), .B(b[1]), .Z(n19298) );
  AND U20237 ( .A(a[801]), .B(b[3]), .Z(n19297) );
  XOR U20238 ( .A(n19298), .B(n19297), .Z(n19299) );
  XOR U20239 ( .A(n19300), .B(n19299), .Z(n19303) );
  NAND U20240 ( .A(b[0]), .B(a[804]), .Z(n19304) );
  XOR U20241 ( .A(n19303), .B(n19304), .Z(n19305) );
  OR U20242 ( .A(n19282), .B(n19281), .Z(n19286) );
  NANDN U20243 ( .A(n19284), .B(n19283), .Z(n19285) );
  AND U20244 ( .A(n19286), .B(n19285), .Z(n19306) );
  XOR U20245 ( .A(n19305), .B(n19306), .Z(n19294) );
  NANDN U20246 ( .A(n19288), .B(n19287), .Z(n19292) );
  OR U20247 ( .A(n19290), .B(n19289), .Z(n19291) );
  AND U20248 ( .A(n19292), .B(n19291), .Z(n19295) );
  XOR U20249 ( .A(n19294), .B(n19295), .Z(n19293) );
  XOR U20250 ( .A(n19296), .B(n19293), .Z(n19308) );
  XNOR U20251 ( .A(sreg[1824]), .B(n19308), .Z(n19309) );
  XOR U20252 ( .A(n19310), .B(n19309), .Z(c[1824]) );
  AND U20253 ( .A(b[2]), .B(a[803]), .Z(n19319) );
  AND U20254 ( .A(a[804]), .B(b[1]), .Z(n19317) );
  AND U20255 ( .A(a[802]), .B(b[3]), .Z(n19316) );
  XOR U20256 ( .A(n19317), .B(n19316), .Z(n19318) );
  XOR U20257 ( .A(n19319), .B(n19318), .Z(n19322) );
  NAND U20258 ( .A(b[0]), .B(a[805]), .Z(n19323) );
  XOR U20259 ( .A(n19322), .B(n19323), .Z(n19324) );
  OR U20260 ( .A(n19298), .B(n19297), .Z(n19302) );
  NANDN U20261 ( .A(n19300), .B(n19299), .Z(n19301) );
  AND U20262 ( .A(n19302), .B(n19301), .Z(n19325) );
  XOR U20263 ( .A(n19324), .B(n19325), .Z(n19313) );
  XOR U20264 ( .A(n19313), .B(n19314), .Z(n19307) );
  XOR U20265 ( .A(n19315), .B(n19307), .Z(n19326) );
  XOR U20266 ( .A(sreg[1825]), .B(n19326), .Z(n19328) );
  NAND U20267 ( .A(sreg[1824]), .B(n19308), .Z(n19312) );
  OR U20268 ( .A(n19310), .B(n19309), .Z(n19311) );
  NAND U20269 ( .A(n19312), .B(n19311), .Z(n19327) );
  XNOR U20270 ( .A(n19328), .B(n19327), .Z(c[1825]) );
  AND U20271 ( .A(b[2]), .B(a[804]), .Z(n19343) );
  AND U20272 ( .A(a[805]), .B(b[1]), .Z(n19341) );
  AND U20273 ( .A(a[803]), .B(b[3]), .Z(n19340) );
  XOR U20274 ( .A(n19341), .B(n19340), .Z(n19342) );
  XOR U20275 ( .A(n19343), .B(n19342), .Z(n19346) );
  NAND U20276 ( .A(b[0]), .B(a[806]), .Z(n19347) );
  XOR U20277 ( .A(n19346), .B(n19347), .Z(n19349) );
  OR U20278 ( .A(n19317), .B(n19316), .Z(n19321) );
  NANDN U20279 ( .A(n19319), .B(n19318), .Z(n19320) );
  NAND U20280 ( .A(n19321), .B(n19320), .Z(n19348) );
  XNOR U20281 ( .A(n19349), .B(n19348), .Z(n19334) );
  XNOR U20282 ( .A(n19334), .B(n19335), .Z(n19337) );
  XOR U20283 ( .A(n19336), .B(n19337), .Z(n19333) );
  NANDN U20284 ( .A(sreg[1825]), .B(n19326), .Z(n19330) );
  OR U20285 ( .A(n19328), .B(n19327), .Z(n19329) );
  AND U20286 ( .A(n19330), .B(n19329), .Z(n19332) );
  XNOR U20287 ( .A(sreg[1826]), .B(n19332), .Z(n19331) );
  XOR U20288 ( .A(n19333), .B(n19331), .Z(c[1826]) );
  NANDN U20289 ( .A(n19335), .B(n19334), .Z(n19339) );
  NAND U20290 ( .A(n19337), .B(n19336), .Z(n19338) );
  NAND U20291 ( .A(n19339), .B(n19338), .Z(n19360) );
  AND U20292 ( .A(b[2]), .B(a[805]), .Z(n19366) );
  AND U20293 ( .A(a[806]), .B(b[1]), .Z(n19364) );
  AND U20294 ( .A(a[804]), .B(b[3]), .Z(n19363) );
  XOR U20295 ( .A(n19364), .B(n19363), .Z(n19365) );
  XOR U20296 ( .A(n19366), .B(n19365), .Z(n19369) );
  NAND U20297 ( .A(b[0]), .B(a[807]), .Z(n19370) );
  XOR U20298 ( .A(n19369), .B(n19370), .Z(n19372) );
  OR U20299 ( .A(n19341), .B(n19340), .Z(n19345) );
  NANDN U20300 ( .A(n19343), .B(n19342), .Z(n19344) );
  NAND U20301 ( .A(n19345), .B(n19344), .Z(n19371) );
  XNOR U20302 ( .A(n19372), .B(n19371), .Z(n19357) );
  NANDN U20303 ( .A(n19347), .B(n19346), .Z(n19351) );
  OR U20304 ( .A(n19349), .B(n19348), .Z(n19350) );
  NAND U20305 ( .A(n19351), .B(n19350), .Z(n19358) );
  XNOR U20306 ( .A(n19357), .B(n19358), .Z(n19359) );
  XNOR U20307 ( .A(n19360), .B(n19359), .Z(n19352) );
  XNOR U20308 ( .A(n19352), .B(sreg[1827]), .Z(n19353) );
  XOR U20309 ( .A(n19354), .B(n19353), .Z(c[1827]) );
  NAND U20310 ( .A(n19352), .B(sreg[1827]), .Z(n19356) );
  OR U20311 ( .A(n19354), .B(n19353), .Z(n19355) );
  NAND U20312 ( .A(n19356), .B(n19355), .Z(n19377) );
  NANDN U20313 ( .A(n19358), .B(n19357), .Z(n19362) );
  NAND U20314 ( .A(n19360), .B(n19359), .Z(n19361) );
  NAND U20315 ( .A(n19362), .B(n19361), .Z(n19383) );
  AND U20316 ( .A(b[2]), .B(a[806]), .Z(n19389) );
  AND U20317 ( .A(a[807]), .B(b[1]), .Z(n19387) );
  AND U20318 ( .A(a[805]), .B(b[3]), .Z(n19386) );
  XOR U20319 ( .A(n19387), .B(n19386), .Z(n19388) );
  XOR U20320 ( .A(n19389), .B(n19388), .Z(n19392) );
  NAND U20321 ( .A(b[0]), .B(a[808]), .Z(n19393) );
  XOR U20322 ( .A(n19392), .B(n19393), .Z(n19395) );
  OR U20323 ( .A(n19364), .B(n19363), .Z(n19368) );
  NANDN U20324 ( .A(n19366), .B(n19365), .Z(n19367) );
  NAND U20325 ( .A(n19368), .B(n19367), .Z(n19394) );
  XNOR U20326 ( .A(n19395), .B(n19394), .Z(n19380) );
  NANDN U20327 ( .A(n19370), .B(n19369), .Z(n19374) );
  OR U20328 ( .A(n19372), .B(n19371), .Z(n19373) );
  NAND U20329 ( .A(n19374), .B(n19373), .Z(n19381) );
  XNOR U20330 ( .A(n19380), .B(n19381), .Z(n19382) );
  XNOR U20331 ( .A(n19383), .B(n19382), .Z(n19375) );
  XOR U20332 ( .A(sreg[1828]), .B(n19375), .Z(n19376) );
  XOR U20333 ( .A(n19377), .B(n19376), .Z(c[1828]) );
  OR U20334 ( .A(n19375), .B(sreg[1828]), .Z(n19379) );
  NANDN U20335 ( .A(n19377), .B(n19376), .Z(n19378) );
  AND U20336 ( .A(n19379), .B(n19378), .Z(n19418) );
  NANDN U20337 ( .A(n19381), .B(n19380), .Z(n19385) );
  NAND U20338 ( .A(n19383), .B(n19382), .Z(n19384) );
  NAND U20339 ( .A(n19385), .B(n19384), .Z(n19402) );
  AND U20340 ( .A(b[2]), .B(a[807]), .Z(n19408) );
  AND U20341 ( .A(a[808]), .B(b[1]), .Z(n19406) );
  AND U20342 ( .A(a[806]), .B(b[3]), .Z(n19405) );
  XOR U20343 ( .A(n19406), .B(n19405), .Z(n19407) );
  XOR U20344 ( .A(n19408), .B(n19407), .Z(n19411) );
  NAND U20345 ( .A(b[0]), .B(a[809]), .Z(n19412) );
  XOR U20346 ( .A(n19411), .B(n19412), .Z(n19414) );
  OR U20347 ( .A(n19387), .B(n19386), .Z(n19391) );
  NANDN U20348 ( .A(n19389), .B(n19388), .Z(n19390) );
  NAND U20349 ( .A(n19391), .B(n19390), .Z(n19413) );
  XNOR U20350 ( .A(n19414), .B(n19413), .Z(n19399) );
  NANDN U20351 ( .A(n19393), .B(n19392), .Z(n19397) );
  OR U20352 ( .A(n19395), .B(n19394), .Z(n19396) );
  NAND U20353 ( .A(n19397), .B(n19396), .Z(n19400) );
  XNOR U20354 ( .A(n19399), .B(n19400), .Z(n19401) );
  XNOR U20355 ( .A(n19402), .B(n19401), .Z(n19417) );
  XOR U20356 ( .A(n19417), .B(sreg[1829]), .Z(n19398) );
  XOR U20357 ( .A(n19418), .B(n19398), .Z(c[1829]) );
  NANDN U20358 ( .A(n19400), .B(n19399), .Z(n19404) );
  NAND U20359 ( .A(n19402), .B(n19401), .Z(n19403) );
  NAND U20360 ( .A(n19404), .B(n19403), .Z(n19425) );
  AND U20361 ( .A(b[2]), .B(a[808]), .Z(n19431) );
  AND U20362 ( .A(a[809]), .B(b[1]), .Z(n19429) );
  AND U20363 ( .A(a[807]), .B(b[3]), .Z(n19428) );
  XOR U20364 ( .A(n19429), .B(n19428), .Z(n19430) );
  XOR U20365 ( .A(n19431), .B(n19430), .Z(n19434) );
  NAND U20366 ( .A(b[0]), .B(a[810]), .Z(n19435) );
  XOR U20367 ( .A(n19434), .B(n19435), .Z(n19437) );
  OR U20368 ( .A(n19406), .B(n19405), .Z(n19410) );
  NANDN U20369 ( .A(n19408), .B(n19407), .Z(n19409) );
  NAND U20370 ( .A(n19410), .B(n19409), .Z(n19436) );
  XNOR U20371 ( .A(n19437), .B(n19436), .Z(n19422) );
  NANDN U20372 ( .A(n19412), .B(n19411), .Z(n19416) );
  OR U20373 ( .A(n19414), .B(n19413), .Z(n19415) );
  NAND U20374 ( .A(n19416), .B(n19415), .Z(n19423) );
  XNOR U20375 ( .A(n19422), .B(n19423), .Z(n19424) );
  XNOR U20376 ( .A(n19425), .B(n19424), .Z(n19421) );
  XOR U20377 ( .A(n19420), .B(sreg[1830]), .Z(n19419) );
  XOR U20378 ( .A(n19421), .B(n19419), .Z(c[1830]) );
  NANDN U20379 ( .A(n19423), .B(n19422), .Z(n19427) );
  NAND U20380 ( .A(n19425), .B(n19424), .Z(n19426) );
  NAND U20381 ( .A(n19427), .B(n19426), .Z(n19443) );
  AND U20382 ( .A(b[2]), .B(a[809]), .Z(n19449) );
  AND U20383 ( .A(a[810]), .B(b[1]), .Z(n19447) );
  AND U20384 ( .A(a[808]), .B(b[3]), .Z(n19446) );
  XOR U20385 ( .A(n19447), .B(n19446), .Z(n19448) );
  XOR U20386 ( .A(n19449), .B(n19448), .Z(n19452) );
  NAND U20387 ( .A(b[0]), .B(a[811]), .Z(n19453) );
  XOR U20388 ( .A(n19452), .B(n19453), .Z(n19455) );
  OR U20389 ( .A(n19429), .B(n19428), .Z(n19433) );
  NANDN U20390 ( .A(n19431), .B(n19430), .Z(n19432) );
  NAND U20391 ( .A(n19433), .B(n19432), .Z(n19454) );
  XNOR U20392 ( .A(n19455), .B(n19454), .Z(n19440) );
  NANDN U20393 ( .A(n19435), .B(n19434), .Z(n19439) );
  OR U20394 ( .A(n19437), .B(n19436), .Z(n19438) );
  NAND U20395 ( .A(n19439), .B(n19438), .Z(n19441) );
  XNOR U20396 ( .A(n19440), .B(n19441), .Z(n19442) );
  XNOR U20397 ( .A(n19443), .B(n19442), .Z(n19458) );
  XNOR U20398 ( .A(n19458), .B(sreg[1831]), .Z(n19460) );
  XNOR U20399 ( .A(n19459), .B(n19460), .Z(c[1831]) );
  NANDN U20400 ( .A(n19441), .B(n19440), .Z(n19445) );
  NAND U20401 ( .A(n19443), .B(n19442), .Z(n19444) );
  NAND U20402 ( .A(n19445), .B(n19444), .Z(n19467) );
  AND U20403 ( .A(b[2]), .B(a[810]), .Z(n19473) );
  AND U20404 ( .A(a[811]), .B(b[1]), .Z(n19471) );
  AND U20405 ( .A(a[809]), .B(b[3]), .Z(n19470) );
  XOR U20406 ( .A(n19471), .B(n19470), .Z(n19472) );
  XOR U20407 ( .A(n19473), .B(n19472), .Z(n19476) );
  NAND U20408 ( .A(b[0]), .B(a[812]), .Z(n19477) );
  XOR U20409 ( .A(n19476), .B(n19477), .Z(n19479) );
  OR U20410 ( .A(n19447), .B(n19446), .Z(n19451) );
  NANDN U20411 ( .A(n19449), .B(n19448), .Z(n19450) );
  NAND U20412 ( .A(n19451), .B(n19450), .Z(n19478) );
  XNOR U20413 ( .A(n19479), .B(n19478), .Z(n19464) );
  NANDN U20414 ( .A(n19453), .B(n19452), .Z(n19457) );
  OR U20415 ( .A(n19455), .B(n19454), .Z(n19456) );
  NAND U20416 ( .A(n19457), .B(n19456), .Z(n19465) );
  XNOR U20417 ( .A(n19464), .B(n19465), .Z(n19466) );
  XOR U20418 ( .A(n19467), .B(n19466), .Z(n19483) );
  NAND U20419 ( .A(n19458), .B(sreg[1831]), .Z(n19462) );
  NANDN U20420 ( .A(n19460), .B(n19459), .Z(n19461) );
  NAND U20421 ( .A(n19462), .B(n19461), .Z(n19482) );
  XNOR U20422 ( .A(sreg[1832]), .B(n19482), .Z(n19463) );
  XOR U20423 ( .A(n19483), .B(n19463), .Z(c[1832]) );
  NANDN U20424 ( .A(n19465), .B(n19464), .Z(n19469) );
  NAND U20425 ( .A(n19467), .B(n19466), .Z(n19468) );
  NAND U20426 ( .A(n19469), .B(n19468), .Z(n19488) );
  AND U20427 ( .A(b[2]), .B(a[811]), .Z(n19494) );
  AND U20428 ( .A(a[812]), .B(b[1]), .Z(n19492) );
  AND U20429 ( .A(a[810]), .B(b[3]), .Z(n19491) );
  XOR U20430 ( .A(n19492), .B(n19491), .Z(n19493) );
  XOR U20431 ( .A(n19494), .B(n19493), .Z(n19497) );
  NAND U20432 ( .A(b[0]), .B(a[813]), .Z(n19498) );
  XOR U20433 ( .A(n19497), .B(n19498), .Z(n19500) );
  OR U20434 ( .A(n19471), .B(n19470), .Z(n19475) );
  NANDN U20435 ( .A(n19473), .B(n19472), .Z(n19474) );
  NAND U20436 ( .A(n19475), .B(n19474), .Z(n19499) );
  XNOR U20437 ( .A(n19500), .B(n19499), .Z(n19485) );
  NANDN U20438 ( .A(n19477), .B(n19476), .Z(n19481) );
  OR U20439 ( .A(n19479), .B(n19478), .Z(n19480) );
  NAND U20440 ( .A(n19481), .B(n19480), .Z(n19486) );
  XNOR U20441 ( .A(n19485), .B(n19486), .Z(n19487) );
  XNOR U20442 ( .A(n19488), .B(n19487), .Z(n19504) );
  XOR U20443 ( .A(n19503), .B(sreg[1833]), .Z(n19484) );
  XOR U20444 ( .A(n19504), .B(n19484), .Z(c[1833]) );
  NANDN U20445 ( .A(n19486), .B(n19485), .Z(n19490) );
  NAND U20446 ( .A(n19488), .B(n19487), .Z(n19489) );
  NAND U20447 ( .A(n19490), .B(n19489), .Z(n19509) );
  AND U20448 ( .A(b[2]), .B(a[812]), .Z(n19515) );
  AND U20449 ( .A(a[813]), .B(b[1]), .Z(n19513) );
  AND U20450 ( .A(a[811]), .B(b[3]), .Z(n19512) );
  XOR U20451 ( .A(n19513), .B(n19512), .Z(n19514) );
  XOR U20452 ( .A(n19515), .B(n19514), .Z(n19518) );
  NAND U20453 ( .A(b[0]), .B(a[814]), .Z(n19519) );
  XOR U20454 ( .A(n19518), .B(n19519), .Z(n19521) );
  OR U20455 ( .A(n19492), .B(n19491), .Z(n19496) );
  NANDN U20456 ( .A(n19494), .B(n19493), .Z(n19495) );
  NAND U20457 ( .A(n19496), .B(n19495), .Z(n19520) );
  XNOR U20458 ( .A(n19521), .B(n19520), .Z(n19506) );
  NANDN U20459 ( .A(n19498), .B(n19497), .Z(n19502) );
  OR U20460 ( .A(n19500), .B(n19499), .Z(n19501) );
  NAND U20461 ( .A(n19502), .B(n19501), .Z(n19507) );
  XNOR U20462 ( .A(n19506), .B(n19507), .Z(n19508) );
  XOR U20463 ( .A(n19509), .B(n19508), .Z(n19525) );
  XOR U20464 ( .A(sreg[1834]), .B(n19524), .Z(n19505) );
  XOR U20465 ( .A(n19525), .B(n19505), .Z(c[1834]) );
  NANDN U20466 ( .A(n19507), .B(n19506), .Z(n19511) );
  NAND U20467 ( .A(n19509), .B(n19508), .Z(n19510) );
  NAND U20468 ( .A(n19511), .B(n19510), .Z(n19532) );
  AND U20469 ( .A(b[2]), .B(a[813]), .Z(n19538) );
  AND U20470 ( .A(a[814]), .B(b[1]), .Z(n19536) );
  AND U20471 ( .A(a[812]), .B(b[3]), .Z(n19535) );
  XOR U20472 ( .A(n19536), .B(n19535), .Z(n19537) );
  XOR U20473 ( .A(n19538), .B(n19537), .Z(n19541) );
  NAND U20474 ( .A(b[0]), .B(a[815]), .Z(n19542) );
  XOR U20475 ( .A(n19541), .B(n19542), .Z(n19544) );
  OR U20476 ( .A(n19513), .B(n19512), .Z(n19517) );
  NANDN U20477 ( .A(n19515), .B(n19514), .Z(n19516) );
  NAND U20478 ( .A(n19517), .B(n19516), .Z(n19543) );
  XNOR U20479 ( .A(n19544), .B(n19543), .Z(n19529) );
  NANDN U20480 ( .A(n19519), .B(n19518), .Z(n19523) );
  OR U20481 ( .A(n19521), .B(n19520), .Z(n19522) );
  NAND U20482 ( .A(n19523), .B(n19522), .Z(n19530) );
  XNOR U20483 ( .A(n19529), .B(n19530), .Z(n19531) );
  XOR U20484 ( .A(n19532), .B(n19531), .Z(n19528) );
  XNOR U20485 ( .A(sreg[1835]), .B(n19527), .Z(n19526) );
  XOR U20486 ( .A(n19528), .B(n19526), .Z(c[1835]) );
  NANDN U20487 ( .A(n19530), .B(n19529), .Z(n19534) );
  NAND U20488 ( .A(n19532), .B(n19531), .Z(n19533) );
  NAND U20489 ( .A(n19534), .B(n19533), .Z(n19550) );
  AND U20490 ( .A(b[2]), .B(a[814]), .Z(n19556) );
  AND U20491 ( .A(a[815]), .B(b[1]), .Z(n19554) );
  AND U20492 ( .A(a[813]), .B(b[3]), .Z(n19553) );
  XOR U20493 ( .A(n19554), .B(n19553), .Z(n19555) );
  XOR U20494 ( .A(n19556), .B(n19555), .Z(n19559) );
  NAND U20495 ( .A(b[0]), .B(a[816]), .Z(n19560) );
  XOR U20496 ( .A(n19559), .B(n19560), .Z(n19562) );
  OR U20497 ( .A(n19536), .B(n19535), .Z(n19540) );
  NANDN U20498 ( .A(n19538), .B(n19537), .Z(n19539) );
  NAND U20499 ( .A(n19540), .B(n19539), .Z(n19561) );
  XNOR U20500 ( .A(n19562), .B(n19561), .Z(n19547) );
  NANDN U20501 ( .A(n19542), .B(n19541), .Z(n19546) );
  OR U20502 ( .A(n19544), .B(n19543), .Z(n19545) );
  NAND U20503 ( .A(n19546), .B(n19545), .Z(n19548) );
  XNOR U20504 ( .A(n19547), .B(n19548), .Z(n19549) );
  XNOR U20505 ( .A(n19550), .B(n19549), .Z(n19565) );
  XNOR U20506 ( .A(n19565), .B(sreg[1836]), .Z(n19566) );
  XOR U20507 ( .A(n19567), .B(n19566), .Z(c[1836]) );
  NANDN U20508 ( .A(n19548), .B(n19547), .Z(n19552) );
  NAND U20509 ( .A(n19550), .B(n19549), .Z(n19551) );
  NAND U20510 ( .A(n19552), .B(n19551), .Z(n19574) );
  AND U20511 ( .A(b[2]), .B(a[815]), .Z(n19580) );
  AND U20512 ( .A(a[816]), .B(b[1]), .Z(n19578) );
  AND U20513 ( .A(a[814]), .B(b[3]), .Z(n19577) );
  XOR U20514 ( .A(n19578), .B(n19577), .Z(n19579) );
  XOR U20515 ( .A(n19580), .B(n19579), .Z(n19583) );
  NAND U20516 ( .A(b[0]), .B(a[817]), .Z(n19584) );
  XOR U20517 ( .A(n19583), .B(n19584), .Z(n19586) );
  OR U20518 ( .A(n19554), .B(n19553), .Z(n19558) );
  NANDN U20519 ( .A(n19556), .B(n19555), .Z(n19557) );
  NAND U20520 ( .A(n19558), .B(n19557), .Z(n19585) );
  XNOR U20521 ( .A(n19586), .B(n19585), .Z(n19571) );
  NANDN U20522 ( .A(n19560), .B(n19559), .Z(n19564) );
  OR U20523 ( .A(n19562), .B(n19561), .Z(n19563) );
  NAND U20524 ( .A(n19564), .B(n19563), .Z(n19572) );
  XNOR U20525 ( .A(n19571), .B(n19572), .Z(n19573) );
  XOR U20526 ( .A(n19574), .B(n19573), .Z(n19590) );
  NAND U20527 ( .A(n19565), .B(sreg[1836]), .Z(n19569) );
  OR U20528 ( .A(n19567), .B(n19566), .Z(n19568) );
  NAND U20529 ( .A(n19569), .B(n19568), .Z(n19589) );
  XNOR U20530 ( .A(sreg[1837]), .B(n19589), .Z(n19570) );
  XOR U20531 ( .A(n19590), .B(n19570), .Z(c[1837]) );
  NANDN U20532 ( .A(n19572), .B(n19571), .Z(n19576) );
  NAND U20533 ( .A(n19574), .B(n19573), .Z(n19575) );
  NAND U20534 ( .A(n19576), .B(n19575), .Z(n19597) );
  AND U20535 ( .A(b[2]), .B(a[816]), .Z(n19603) );
  AND U20536 ( .A(a[817]), .B(b[1]), .Z(n19601) );
  AND U20537 ( .A(a[815]), .B(b[3]), .Z(n19600) );
  XOR U20538 ( .A(n19601), .B(n19600), .Z(n19602) );
  XOR U20539 ( .A(n19603), .B(n19602), .Z(n19606) );
  NAND U20540 ( .A(b[0]), .B(a[818]), .Z(n19607) );
  XOR U20541 ( .A(n19606), .B(n19607), .Z(n19609) );
  OR U20542 ( .A(n19578), .B(n19577), .Z(n19582) );
  NANDN U20543 ( .A(n19580), .B(n19579), .Z(n19581) );
  NAND U20544 ( .A(n19582), .B(n19581), .Z(n19608) );
  XNOR U20545 ( .A(n19609), .B(n19608), .Z(n19594) );
  NANDN U20546 ( .A(n19584), .B(n19583), .Z(n19588) );
  OR U20547 ( .A(n19586), .B(n19585), .Z(n19587) );
  NAND U20548 ( .A(n19588), .B(n19587), .Z(n19595) );
  XNOR U20549 ( .A(n19594), .B(n19595), .Z(n19596) );
  XOR U20550 ( .A(n19597), .B(n19596), .Z(n19593) );
  XNOR U20551 ( .A(sreg[1838]), .B(n19592), .Z(n19591) );
  XOR U20552 ( .A(n19593), .B(n19591), .Z(c[1838]) );
  NANDN U20553 ( .A(n19595), .B(n19594), .Z(n19599) );
  NAND U20554 ( .A(n19597), .B(n19596), .Z(n19598) );
  NAND U20555 ( .A(n19599), .B(n19598), .Z(n19615) );
  AND U20556 ( .A(b[2]), .B(a[817]), .Z(n19621) );
  AND U20557 ( .A(a[818]), .B(b[1]), .Z(n19619) );
  AND U20558 ( .A(a[816]), .B(b[3]), .Z(n19618) );
  XOR U20559 ( .A(n19619), .B(n19618), .Z(n19620) );
  XOR U20560 ( .A(n19621), .B(n19620), .Z(n19624) );
  NAND U20561 ( .A(b[0]), .B(a[819]), .Z(n19625) );
  XOR U20562 ( .A(n19624), .B(n19625), .Z(n19627) );
  OR U20563 ( .A(n19601), .B(n19600), .Z(n19605) );
  NANDN U20564 ( .A(n19603), .B(n19602), .Z(n19604) );
  NAND U20565 ( .A(n19605), .B(n19604), .Z(n19626) );
  XNOR U20566 ( .A(n19627), .B(n19626), .Z(n19612) );
  NANDN U20567 ( .A(n19607), .B(n19606), .Z(n19611) );
  OR U20568 ( .A(n19609), .B(n19608), .Z(n19610) );
  NAND U20569 ( .A(n19611), .B(n19610), .Z(n19613) );
  XNOR U20570 ( .A(n19612), .B(n19613), .Z(n19614) );
  XNOR U20571 ( .A(n19615), .B(n19614), .Z(n19630) );
  XNOR U20572 ( .A(n19630), .B(sreg[1839]), .Z(n19631) );
  XOR U20573 ( .A(n19632), .B(n19631), .Z(c[1839]) );
  NANDN U20574 ( .A(n19613), .B(n19612), .Z(n19617) );
  NAND U20575 ( .A(n19615), .B(n19614), .Z(n19616) );
  NAND U20576 ( .A(n19617), .B(n19616), .Z(n19641) );
  AND U20577 ( .A(b[2]), .B(a[818]), .Z(n19653) );
  AND U20578 ( .A(a[819]), .B(b[1]), .Z(n19651) );
  AND U20579 ( .A(a[817]), .B(b[3]), .Z(n19650) );
  XOR U20580 ( .A(n19651), .B(n19650), .Z(n19652) );
  XOR U20581 ( .A(n19653), .B(n19652), .Z(n19644) );
  NAND U20582 ( .A(b[0]), .B(a[820]), .Z(n19645) );
  XOR U20583 ( .A(n19644), .B(n19645), .Z(n19647) );
  OR U20584 ( .A(n19619), .B(n19618), .Z(n19623) );
  NANDN U20585 ( .A(n19621), .B(n19620), .Z(n19622) );
  NAND U20586 ( .A(n19623), .B(n19622), .Z(n19646) );
  XNOR U20587 ( .A(n19647), .B(n19646), .Z(n19638) );
  NANDN U20588 ( .A(n19625), .B(n19624), .Z(n19629) );
  OR U20589 ( .A(n19627), .B(n19626), .Z(n19628) );
  NAND U20590 ( .A(n19629), .B(n19628), .Z(n19639) );
  XNOR U20591 ( .A(n19638), .B(n19639), .Z(n19640) );
  XOR U20592 ( .A(n19641), .B(n19640), .Z(n19637) );
  NAND U20593 ( .A(n19630), .B(sreg[1839]), .Z(n19634) );
  OR U20594 ( .A(n19632), .B(n19631), .Z(n19633) );
  NAND U20595 ( .A(n19634), .B(n19633), .Z(n19636) );
  XNOR U20596 ( .A(sreg[1840]), .B(n19636), .Z(n19635) );
  XOR U20597 ( .A(n19637), .B(n19635), .Z(c[1840]) );
  NANDN U20598 ( .A(n19639), .B(n19638), .Z(n19643) );
  NAND U20599 ( .A(n19641), .B(n19640), .Z(n19642) );
  NAND U20600 ( .A(n19643), .B(n19642), .Z(n19671) );
  NANDN U20601 ( .A(n19645), .B(n19644), .Z(n19649) );
  OR U20602 ( .A(n19647), .B(n19646), .Z(n19648) );
  NAND U20603 ( .A(n19649), .B(n19648), .Z(n19668) );
  AND U20604 ( .A(b[2]), .B(a[819]), .Z(n19659) );
  AND U20605 ( .A(a[820]), .B(b[1]), .Z(n19657) );
  AND U20606 ( .A(a[818]), .B(b[3]), .Z(n19656) );
  XOR U20607 ( .A(n19657), .B(n19656), .Z(n19658) );
  XOR U20608 ( .A(n19659), .B(n19658), .Z(n19662) );
  NAND U20609 ( .A(b[0]), .B(a[821]), .Z(n19663) );
  XNOR U20610 ( .A(n19662), .B(n19663), .Z(n19664) );
  OR U20611 ( .A(n19651), .B(n19650), .Z(n19655) );
  NANDN U20612 ( .A(n19653), .B(n19652), .Z(n19654) );
  AND U20613 ( .A(n19655), .B(n19654), .Z(n19665) );
  XNOR U20614 ( .A(n19664), .B(n19665), .Z(n19669) );
  XNOR U20615 ( .A(n19668), .B(n19669), .Z(n19670) );
  XNOR U20616 ( .A(n19671), .B(n19670), .Z(n19674) );
  XNOR U20617 ( .A(sreg[1841]), .B(n19674), .Z(n19675) );
  XOR U20618 ( .A(n19676), .B(n19675), .Z(c[1841]) );
  AND U20619 ( .A(b[2]), .B(a[820]), .Z(n19691) );
  AND U20620 ( .A(a[821]), .B(b[1]), .Z(n19689) );
  AND U20621 ( .A(a[819]), .B(b[3]), .Z(n19688) );
  XOR U20622 ( .A(n19689), .B(n19688), .Z(n19690) );
  XOR U20623 ( .A(n19691), .B(n19690), .Z(n19694) );
  NAND U20624 ( .A(b[0]), .B(a[822]), .Z(n19695) );
  XOR U20625 ( .A(n19694), .B(n19695), .Z(n19697) );
  OR U20626 ( .A(n19657), .B(n19656), .Z(n19661) );
  NANDN U20627 ( .A(n19659), .B(n19658), .Z(n19660) );
  NAND U20628 ( .A(n19661), .B(n19660), .Z(n19696) );
  XNOR U20629 ( .A(n19697), .B(n19696), .Z(n19682) );
  NANDN U20630 ( .A(n19663), .B(n19662), .Z(n19667) );
  NAND U20631 ( .A(n19665), .B(n19664), .Z(n19666) );
  NAND U20632 ( .A(n19667), .B(n19666), .Z(n19683) );
  XNOR U20633 ( .A(n19682), .B(n19683), .Z(n19684) );
  NANDN U20634 ( .A(n19669), .B(n19668), .Z(n19673) );
  NANDN U20635 ( .A(n19671), .B(n19670), .Z(n19672) );
  AND U20636 ( .A(n19673), .B(n19672), .Z(n19685) );
  XNOR U20637 ( .A(n19684), .B(n19685), .Z(n19681) );
  NAND U20638 ( .A(sreg[1841]), .B(n19674), .Z(n19678) );
  OR U20639 ( .A(n19676), .B(n19675), .Z(n19677) );
  AND U20640 ( .A(n19678), .B(n19677), .Z(n19680) );
  XNOR U20641 ( .A(n19680), .B(sreg[1842]), .Z(n19679) );
  XOR U20642 ( .A(n19681), .B(n19679), .Z(c[1842]) );
  NANDN U20643 ( .A(n19683), .B(n19682), .Z(n19687) );
  NAND U20644 ( .A(n19685), .B(n19684), .Z(n19686) );
  NAND U20645 ( .A(n19687), .B(n19686), .Z(n19720) );
  AND U20646 ( .A(b[2]), .B(a[821]), .Z(n19714) );
  AND U20647 ( .A(a[822]), .B(b[1]), .Z(n19712) );
  AND U20648 ( .A(a[820]), .B(b[3]), .Z(n19711) );
  XOR U20649 ( .A(n19712), .B(n19711), .Z(n19713) );
  XOR U20650 ( .A(n19714), .B(n19713), .Z(n19705) );
  NAND U20651 ( .A(b[0]), .B(a[823]), .Z(n19706) );
  XOR U20652 ( .A(n19705), .B(n19706), .Z(n19708) );
  OR U20653 ( .A(n19689), .B(n19688), .Z(n19693) );
  NANDN U20654 ( .A(n19691), .B(n19690), .Z(n19692) );
  NAND U20655 ( .A(n19693), .B(n19692), .Z(n19707) );
  XNOR U20656 ( .A(n19708), .B(n19707), .Z(n19717) );
  NANDN U20657 ( .A(n19695), .B(n19694), .Z(n19699) );
  OR U20658 ( .A(n19697), .B(n19696), .Z(n19698) );
  NAND U20659 ( .A(n19699), .B(n19698), .Z(n19718) );
  XNOR U20660 ( .A(n19717), .B(n19718), .Z(n19719) );
  XNOR U20661 ( .A(n19720), .B(n19719), .Z(n19700) );
  XNOR U20662 ( .A(n19700), .B(sreg[1843]), .Z(n19702) );
  XNOR U20663 ( .A(n19701), .B(n19702), .Z(c[1843]) );
  NAND U20664 ( .A(n19700), .B(sreg[1843]), .Z(n19704) );
  NANDN U20665 ( .A(n19702), .B(n19701), .Z(n19703) );
  NAND U20666 ( .A(n19704), .B(n19703), .Z(n19742) );
  NANDN U20667 ( .A(n19706), .B(n19705), .Z(n19710) );
  OR U20668 ( .A(n19708), .B(n19707), .Z(n19709) );
  NAND U20669 ( .A(n19710), .B(n19709), .Z(n19736) );
  AND U20670 ( .A(b[2]), .B(a[822]), .Z(n19727) );
  AND U20671 ( .A(a[823]), .B(b[1]), .Z(n19725) );
  AND U20672 ( .A(a[821]), .B(b[3]), .Z(n19724) );
  XOR U20673 ( .A(n19725), .B(n19724), .Z(n19726) );
  XOR U20674 ( .A(n19727), .B(n19726), .Z(n19730) );
  NAND U20675 ( .A(b[0]), .B(a[824]), .Z(n19731) );
  XNOR U20676 ( .A(n19730), .B(n19731), .Z(n19732) );
  OR U20677 ( .A(n19712), .B(n19711), .Z(n19716) );
  NANDN U20678 ( .A(n19714), .B(n19713), .Z(n19715) );
  AND U20679 ( .A(n19716), .B(n19715), .Z(n19733) );
  XNOR U20680 ( .A(n19732), .B(n19733), .Z(n19737) );
  XNOR U20681 ( .A(n19736), .B(n19737), .Z(n19738) );
  NANDN U20682 ( .A(n19718), .B(n19717), .Z(n19722) );
  NAND U20683 ( .A(n19720), .B(n19719), .Z(n19721) );
  AND U20684 ( .A(n19722), .B(n19721), .Z(n19739) );
  XNOR U20685 ( .A(n19738), .B(n19739), .Z(n19743) );
  XOR U20686 ( .A(sreg[1844]), .B(n19743), .Z(n19723) );
  XNOR U20687 ( .A(n19742), .B(n19723), .Z(c[1844]) );
  AND U20688 ( .A(b[2]), .B(a[823]), .Z(n19756) );
  AND U20689 ( .A(a[824]), .B(b[1]), .Z(n19754) );
  AND U20690 ( .A(a[822]), .B(b[3]), .Z(n19753) );
  XOR U20691 ( .A(n19754), .B(n19753), .Z(n19755) );
  XOR U20692 ( .A(n19756), .B(n19755), .Z(n19759) );
  NAND U20693 ( .A(b[0]), .B(a[825]), .Z(n19760) );
  XOR U20694 ( .A(n19759), .B(n19760), .Z(n19762) );
  OR U20695 ( .A(n19725), .B(n19724), .Z(n19729) );
  NANDN U20696 ( .A(n19727), .B(n19726), .Z(n19728) );
  NAND U20697 ( .A(n19729), .B(n19728), .Z(n19761) );
  XNOR U20698 ( .A(n19762), .B(n19761), .Z(n19747) );
  NANDN U20699 ( .A(n19731), .B(n19730), .Z(n19735) );
  NAND U20700 ( .A(n19733), .B(n19732), .Z(n19734) );
  NAND U20701 ( .A(n19735), .B(n19734), .Z(n19748) );
  XNOR U20702 ( .A(n19747), .B(n19748), .Z(n19749) );
  NANDN U20703 ( .A(n19737), .B(n19736), .Z(n19741) );
  NAND U20704 ( .A(n19739), .B(n19738), .Z(n19740) );
  AND U20705 ( .A(n19741), .B(n19740), .Z(n19750) );
  XNOR U20706 ( .A(n19749), .B(n19750), .Z(n19746) );
  XOR U20707 ( .A(n19745), .B(sreg[1845]), .Z(n19744) );
  XOR U20708 ( .A(n19746), .B(n19744), .Z(c[1845]) );
  NANDN U20709 ( .A(n19748), .B(n19747), .Z(n19752) );
  NAND U20710 ( .A(n19750), .B(n19749), .Z(n19751) );
  NAND U20711 ( .A(n19752), .B(n19751), .Z(n19785) );
  AND U20712 ( .A(b[2]), .B(a[824]), .Z(n19779) );
  AND U20713 ( .A(a[825]), .B(b[1]), .Z(n19777) );
  AND U20714 ( .A(a[823]), .B(b[3]), .Z(n19776) );
  XOR U20715 ( .A(n19777), .B(n19776), .Z(n19778) );
  XOR U20716 ( .A(n19779), .B(n19778), .Z(n19770) );
  NAND U20717 ( .A(b[0]), .B(a[826]), .Z(n19771) );
  XOR U20718 ( .A(n19770), .B(n19771), .Z(n19773) );
  OR U20719 ( .A(n19754), .B(n19753), .Z(n19758) );
  NANDN U20720 ( .A(n19756), .B(n19755), .Z(n19757) );
  NAND U20721 ( .A(n19758), .B(n19757), .Z(n19772) );
  XNOR U20722 ( .A(n19773), .B(n19772), .Z(n19782) );
  NANDN U20723 ( .A(n19760), .B(n19759), .Z(n19764) );
  OR U20724 ( .A(n19762), .B(n19761), .Z(n19763) );
  NAND U20725 ( .A(n19764), .B(n19763), .Z(n19783) );
  XNOR U20726 ( .A(n19782), .B(n19783), .Z(n19784) );
  XNOR U20727 ( .A(n19785), .B(n19784), .Z(n19765) );
  XNOR U20728 ( .A(n19765), .B(sreg[1846]), .Z(n19767) );
  XNOR U20729 ( .A(n19766), .B(n19767), .Z(c[1846]) );
  NAND U20730 ( .A(n19765), .B(sreg[1846]), .Z(n19769) );
  NANDN U20731 ( .A(n19767), .B(n19766), .Z(n19768) );
  NAND U20732 ( .A(n19769), .B(n19768), .Z(n19807) );
  NANDN U20733 ( .A(n19771), .B(n19770), .Z(n19775) );
  OR U20734 ( .A(n19773), .B(n19772), .Z(n19774) );
  NAND U20735 ( .A(n19775), .B(n19774), .Z(n19801) );
  AND U20736 ( .A(b[2]), .B(a[825]), .Z(n19792) );
  AND U20737 ( .A(a[826]), .B(b[1]), .Z(n19790) );
  AND U20738 ( .A(a[824]), .B(b[3]), .Z(n19789) );
  XOR U20739 ( .A(n19790), .B(n19789), .Z(n19791) );
  XOR U20740 ( .A(n19792), .B(n19791), .Z(n19795) );
  NAND U20741 ( .A(b[0]), .B(a[827]), .Z(n19796) );
  XNOR U20742 ( .A(n19795), .B(n19796), .Z(n19797) );
  OR U20743 ( .A(n19777), .B(n19776), .Z(n19781) );
  NANDN U20744 ( .A(n19779), .B(n19778), .Z(n19780) );
  AND U20745 ( .A(n19781), .B(n19780), .Z(n19798) );
  XNOR U20746 ( .A(n19797), .B(n19798), .Z(n19802) );
  XNOR U20747 ( .A(n19801), .B(n19802), .Z(n19803) );
  NANDN U20748 ( .A(n19783), .B(n19782), .Z(n19787) );
  NAND U20749 ( .A(n19785), .B(n19784), .Z(n19786) );
  AND U20750 ( .A(n19787), .B(n19786), .Z(n19804) );
  XNOR U20751 ( .A(n19803), .B(n19804), .Z(n19808) );
  XOR U20752 ( .A(sreg[1847]), .B(n19808), .Z(n19788) );
  XNOR U20753 ( .A(n19807), .B(n19788), .Z(c[1847]) );
  AND U20754 ( .A(b[2]), .B(a[826]), .Z(n19821) );
  AND U20755 ( .A(a[827]), .B(b[1]), .Z(n19819) );
  AND U20756 ( .A(a[825]), .B(b[3]), .Z(n19818) );
  XOR U20757 ( .A(n19819), .B(n19818), .Z(n19820) );
  XOR U20758 ( .A(n19821), .B(n19820), .Z(n19824) );
  NAND U20759 ( .A(b[0]), .B(a[828]), .Z(n19825) );
  XOR U20760 ( .A(n19824), .B(n19825), .Z(n19827) );
  OR U20761 ( .A(n19790), .B(n19789), .Z(n19794) );
  NANDN U20762 ( .A(n19792), .B(n19791), .Z(n19793) );
  NAND U20763 ( .A(n19794), .B(n19793), .Z(n19826) );
  XNOR U20764 ( .A(n19827), .B(n19826), .Z(n19812) );
  NANDN U20765 ( .A(n19796), .B(n19795), .Z(n19800) );
  NAND U20766 ( .A(n19798), .B(n19797), .Z(n19799) );
  NAND U20767 ( .A(n19800), .B(n19799), .Z(n19813) );
  XNOR U20768 ( .A(n19812), .B(n19813), .Z(n19814) );
  NANDN U20769 ( .A(n19802), .B(n19801), .Z(n19806) );
  NAND U20770 ( .A(n19804), .B(n19803), .Z(n19805) );
  AND U20771 ( .A(n19806), .B(n19805), .Z(n19815) );
  XNOR U20772 ( .A(n19814), .B(n19815), .Z(n19811) );
  XOR U20773 ( .A(n19810), .B(sreg[1848]), .Z(n19809) );
  XOR U20774 ( .A(n19811), .B(n19809), .Z(c[1848]) );
  NANDN U20775 ( .A(n19813), .B(n19812), .Z(n19817) );
  NAND U20776 ( .A(n19815), .B(n19814), .Z(n19816) );
  NAND U20777 ( .A(n19817), .B(n19816), .Z(n19850) );
  AND U20778 ( .A(b[2]), .B(a[827]), .Z(n19844) );
  AND U20779 ( .A(a[828]), .B(b[1]), .Z(n19842) );
  AND U20780 ( .A(a[826]), .B(b[3]), .Z(n19841) );
  XOR U20781 ( .A(n19842), .B(n19841), .Z(n19843) );
  XOR U20782 ( .A(n19844), .B(n19843), .Z(n19835) );
  NAND U20783 ( .A(b[0]), .B(a[829]), .Z(n19836) );
  XOR U20784 ( .A(n19835), .B(n19836), .Z(n19838) );
  OR U20785 ( .A(n19819), .B(n19818), .Z(n19823) );
  NANDN U20786 ( .A(n19821), .B(n19820), .Z(n19822) );
  NAND U20787 ( .A(n19823), .B(n19822), .Z(n19837) );
  XNOR U20788 ( .A(n19838), .B(n19837), .Z(n19847) );
  NANDN U20789 ( .A(n19825), .B(n19824), .Z(n19829) );
  OR U20790 ( .A(n19827), .B(n19826), .Z(n19828) );
  NAND U20791 ( .A(n19829), .B(n19828), .Z(n19848) );
  XNOR U20792 ( .A(n19847), .B(n19848), .Z(n19849) );
  XNOR U20793 ( .A(n19850), .B(n19849), .Z(n19830) );
  XNOR U20794 ( .A(n19830), .B(sreg[1849]), .Z(n19832) );
  XNOR U20795 ( .A(n19831), .B(n19832), .Z(c[1849]) );
  NAND U20796 ( .A(n19830), .B(sreg[1849]), .Z(n19834) );
  NANDN U20797 ( .A(n19832), .B(n19831), .Z(n19833) );
  NAND U20798 ( .A(n19834), .B(n19833), .Z(n19854) );
  NANDN U20799 ( .A(n19836), .B(n19835), .Z(n19840) );
  OR U20800 ( .A(n19838), .B(n19837), .Z(n19839) );
  NAND U20801 ( .A(n19840), .B(n19839), .Z(n19868) );
  AND U20802 ( .A(b[2]), .B(a[828]), .Z(n19859) );
  AND U20803 ( .A(a[829]), .B(b[1]), .Z(n19857) );
  AND U20804 ( .A(a[827]), .B(b[3]), .Z(n19856) );
  XOR U20805 ( .A(n19857), .B(n19856), .Z(n19858) );
  XOR U20806 ( .A(n19859), .B(n19858), .Z(n19862) );
  NAND U20807 ( .A(b[0]), .B(a[830]), .Z(n19863) );
  XNOR U20808 ( .A(n19862), .B(n19863), .Z(n19864) );
  OR U20809 ( .A(n19842), .B(n19841), .Z(n19846) );
  NANDN U20810 ( .A(n19844), .B(n19843), .Z(n19845) );
  AND U20811 ( .A(n19846), .B(n19845), .Z(n19865) );
  XNOR U20812 ( .A(n19864), .B(n19865), .Z(n19869) );
  XNOR U20813 ( .A(n19868), .B(n19869), .Z(n19870) );
  NANDN U20814 ( .A(n19848), .B(n19847), .Z(n19852) );
  NAND U20815 ( .A(n19850), .B(n19849), .Z(n19851) );
  AND U20816 ( .A(n19852), .B(n19851), .Z(n19871) );
  XNOR U20817 ( .A(n19870), .B(n19871), .Z(n19855) );
  XOR U20818 ( .A(sreg[1850]), .B(n19855), .Z(n19853) );
  XNOR U20819 ( .A(n19854), .B(n19853), .Z(c[1850]) );
  AND U20820 ( .A(b[2]), .B(a[829]), .Z(n19883) );
  AND U20821 ( .A(a[830]), .B(b[1]), .Z(n19881) );
  AND U20822 ( .A(a[828]), .B(b[3]), .Z(n19880) );
  XOR U20823 ( .A(n19881), .B(n19880), .Z(n19882) );
  XOR U20824 ( .A(n19883), .B(n19882), .Z(n19886) );
  NAND U20825 ( .A(b[0]), .B(a[831]), .Z(n19887) );
  XOR U20826 ( .A(n19886), .B(n19887), .Z(n19889) );
  OR U20827 ( .A(n19857), .B(n19856), .Z(n19861) );
  NANDN U20828 ( .A(n19859), .B(n19858), .Z(n19860) );
  NAND U20829 ( .A(n19861), .B(n19860), .Z(n19888) );
  XNOR U20830 ( .A(n19889), .B(n19888), .Z(n19874) );
  NANDN U20831 ( .A(n19863), .B(n19862), .Z(n19867) );
  NAND U20832 ( .A(n19865), .B(n19864), .Z(n19866) );
  NAND U20833 ( .A(n19867), .B(n19866), .Z(n19875) );
  XNOR U20834 ( .A(n19874), .B(n19875), .Z(n19876) );
  NANDN U20835 ( .A(n19869), .B(n19868), .Z(n19873) );
  NAND U20836 ( .A(n19871), .B(n19870), .Z(n19872) );
  NAND U20837 ( .A(n19873), .B(n19872), .Z(n19877) );
  XOR U20838 ( .A(n19876), .B(n19877), .Z(n19892) );
  XNOR U20839 ( .A(n19892), .B(sreg[1851]), .Z(n19893) );
  XOR U20840 ( .A(n19894), .B(n19893), .Z(c[1851]) );
  NANDN U20841 ( .A(n19875), .B(n19874), .Z(n19879) );
  NANDN U20842 ( .A(n19877), .B(n19876), .Z(n19878) );
  NAND U20843 ( .A(n19879), .B(n19878), .Z(n19900) );
  AND U20844 ( .A(b[2]), .B(a[830]), .Z(n19906) );
  AND U20845 ( .A(a[831]), .B(b[1]), .Z(n19904) );
  AND U20846 ( .A(a[829]), .B(b[3]), .Z(n19903) );
  XOR U20847 ( .A(n19904), .B(n19903), .Z(n19905) );
  XOR U20848 ( .A(n19906), .B(n19905), .Z(n19909) );
  NAND U20849 ( .A(b[0]), .B(a[832]), .Z(n19910) );
  XOR U20850 ( .A(n19909), .B(n19910), .Z(n19912) );
  OR U20851 ( .A(n19881), .B(n19880), .Z(n19885) );
  NANDN U20852 ( .A(n19883), .B(n19882), .Z(n19884) );
  NAND U20853 ( .A(n19885), .B(n19884), .Z(n19911) );
  XNOR U20854 ( .A(n19912), .B(n19911), .Z(n19897) );
  NANDN U20855 ( .A(n19887), .B(n19886), .Z(n19891) );
  OR U20856 ( .A(n19889), .B(n19888), .Z(n19890) );
  NAND U20857 ( .A(n19891), .B(n19890), .Z(n19898) );
  XNOR U20858 ( .A(n19897), .B(n19898), .Z(n19899) );
  XNOR U20859 ( .A(n19900), .B(n19899), .Z(n19915) );
  XNOR U20860 ( .A(n19915), .B(sreg[1852]), .Z(n19917) );
  NAND U20861 ( .A(n19892), .B(sreg[1851]), .Z(n19896) );
  OR U20862 ( .A(n19894), .B(n19893), .Z(n19895) );
  AND U20863 ( .A(n19896), .B(n19895), .Z(n19916) );
  XOR U20864 ( .A(n19917), .B(n19916), .Z(c[1852]) );
  NANDN U20865 ( .A(n19898), .B(n19897), .Z(n19902) );
  NAND U20866 ( .A(n19900), .B(n19899), .Z(n19901) );
  NAND U20867 ( .A(n19902), .B(n19901), .Z(n19926) );
  AND U20868 ( .A(b[2]), .B(a[831]), .Z(n19932) );
  AND U20869 ( .A(a[832]), .B(b[1]), .Z(n19930) );
  AND U20870 ( .A(a[830]), .B(b[3]), .Z(n19929) );
  XOR U20871 ( .A(n19930), .B(n19929), .Z(n19931) );
  XOR U20872 ( .A(n19932), .B(n19931), .Z(n19935) );
  NAND U20873 ( .A(b[0]), .B(a[833]), .Z(n19936) );
  XOR U20874 ( .A(n19935), .B(n19936), .Z(n19938) );
  OR U20875 ( .A(n19904), .B(n19903), .Z(n19908) );
  NANDN U20876 ( .A(n19906), .B(n19905), .Z(n19907) );
  NAND U20877 ( .A(n19908), .B(n19907), .Z(n19937) );
  XNOR U20878 ( .A(n19938), .B(n19937), .Z(n19923) );
  NANDN U20879 ( .A(n19910), .B(n19909), .Z(n19914) );
  OR U20880 ( .A(n19912), .B(n19911), .Z(n19913) );
  NAND U20881 ( .A(n19914), .B(n19913), .Z(n19924) );
  XNOR U20882 ( .A(n19923), .B(n19924), .Z(n19925) );
  XOR U20883 ( .A(n19926), .B(n19925), .Z(n19922) );
  NAND U20884 ( .A(n19915), .B(sreg[1852]), .Z(n19919) );
  OR U20885 ( .A(n19917), .B(n19916), .Z(n19918) );
  NAND U20886 ( .A(n19919), .B(n19918), .Z(n19921) );
  XNOR U20887 ( .A(sreg[1853]), .B(n19921), .Z(n19920) );
  XOR U20888 ( .A(n19922), .B(n19920), .Z(c[1853]) );
  NANDN U20889 ( .A(n19924), .B(n19923), .Z(n19928) );
  NAND U20890 ( .A(n19926), .B(n19925), .Z(n19927) );
  NAND U20891 ( .A(n19928), .B(n19927), .Z(n19944) );
  AND U20892 ( .A(b[2]), .B(a[832]), .Z(n19950) );
  AND U20893 ( .A(a[833]), .B(b[1]), .Z(n19948) );
  AND U20894 ( .A(a[831]), .B(b[3]), .Z(n19947) );
  XOR U20895 ( .A(n19948), .B(n19947), .Z(n19949) );
  XOR U20896 ( .A(n19950), .B(n19949), .Z(n19953) );
  NAND U20897 ( .A(b[0]), .B(a[834]), .Z(n19954) );
  XOR U20898 ( .A(n19953), .B(n19954), .Z(n19956) );
  OR U20899 ( .A(n19930), .B(n19929), .Z(n19934) );
  NANDN U20900 ( .A(n19932), .B(n19931), .Z(n19933) );
  NAND U20901 ( .A(n19934), .B(n19933), .Z(n19955) );
  XNOR U20902 ( .A(n19956), .B(n19955), .Z(n19941) );
  NANDN U20903 ( .A(n19936), .B(n19935), .Z(n19940) );
  OR U20904 ( .A(n19938), .B(n19937), .Z(n19939) );
  NAND U20905 ( .A(n19940), .B(n19939), .Z(n19942) );
  XNOR U20906 ( .A(n19941), .B(n19942), .Z(n19943) );
  XNOR U20907 ( .A(n19944), .B(n19943), .Z(n19959) );
  XNOR U20908 ( .A(n19959), .B(sreg[1854]), .Z(n19960) );
  XOR U20909 ( .A(n19961), .B(n19960), .Z(c[1854]) );
  NANDN U20910 ( .A(n19942), .B(n19941), .Z(n19946) );
  NAND U20911 ( .A(n19944), .B(n19943), .Z(n19945) );
  NAND U20912 ( .A(n19946), .B(n19945), .Z(n19972) );
  AND U20913 ( .A(b[2]), .B(a[833]), .Z(n19978) );
  AND U20914 ( .A(a[834]), .B(b[1]), .Z(n19976) );
  AND U20915 ( .A(a[832]), .B(b[3]), .Z(n19975) );
  XOR U20916 ( .A(n19976), .B(n19975), .Z(n19977) );
  XOR U20917 ( .A(n19978), .B(n19977), .Z(n19981) );
  NAND U20918 ( .A(b[0]), .B(a[835]), .Z(n19982) );
  XOR U20919 ( .A(n19981), .B(n19982), .Z(n19984) );
  OR U20920 ( .A(n19948), .B(n19947), .Z(n19952) );
  NANDN U20921 ( .A(n19950), .B(n19949), .Z(n19951) );
  NAND U20922 ( .A(n19952), .B(n19951), .Z(n19983) );
  XNOR U20923 ( .A(n19984), .B(n19983), .Z(n19969) );
  NANDN U20924 ( .A(n19954), .B(n19953), .Z(n19958) );
  OR U20925 ( .A(n19956), .B(n19955), .Z(n19957) );
  NAND U20926 ( .A(n19958), .B(n19957), .Z(n19970) );
  XNOR U20927 ( .A(n19969), .B(n19970), .Z(n19971) );
  XNOR U20928 ( .A(n19972), .B(n19971), .Z(n19964) );
  XOR U20929 ( .A(sreg[1855]), .B(n19964), .Z(n19965) );
  NAND U20930 ( .A(n19959), .B(sreg[1854]), .Z(n19963) );
  OR U20931 ( .A(n19961), .B(n19960), .Z(n19962) );
  NAND U20932 ( .A(n19963), .B(n19962), .Z(n19966) );
  XOR U20933 ( .A(n19965), .B(n19966), .Z(c[1855]) );
  OR U20934 ( .A(n19964), .B(sreg[1855]), .Z(n19968) );
  NANDN U20935 ( .A(n19966), .B(n19965), .Z(n19967) );
  AND U20936 ( .A(n19968), .B(n19967), .Z(n20006) );
  NANDN U20937 ( .A(n19970), .B(n19969), .Z(n19974) );
  NAND U20938 ( .A(n19972), .B(n19971), .Z(n19973) );
  NAND U20939 ( .A(n19974), .B(n19973), .Z(n19991) );
  AND U20940 ( .A(b[2]), .B(a[834]), .Z(n19997) );
  AND U20941 ( .A(a[835]), .B(b[1]), .Z(n19995) );
  AND U20942 ( .A(a[833]), .B(b[3]), .Z(n19994) );
  XOR U20943 ( .A(n19995), .B(n19994), .Z(n19996) );
  XOR U20944 ( .A(n19997), .B(n19996), .Z(n20000) );
  NAND U20945 ( .A(b[0]), .B(a[836]), .Z(n20001) );
  XOR U20946 ( .A(n20000), .B(n20001), .Z(n20003) );
  OR U20947 ( .A(n19976), .B(n19975), .Z(n19980) );
  NANDN U20948 ( .A(n19978), .B(n19977), .Z(n19979) );
  NAND U20949 ( .A(n19980), .B(n19979), .Z(n20002) );
  XNOR U20950 ( .A(n20003), .B(n20002), .Z(n19988) );
  NANDN U20951 ( .A(n19982), .B(n19981), .Z(n19986) );
  OR U20952 ( .A(n19984), .B(n19983), .Z(n19985) );
  NAND U20953 ( .A(n19986), .B(n19985), .Z(n19989) );
  XNOR U20954 ( .A(n19988), .B(n19989), .Z(n19990) );
  XNOR U20955 ( .A(n19991), .B(n19990), .Z(n20007) );
  XOR U20956 ( .A(sreg[1856]), .B(n20007), .Z(n19987) );
  XOR U20957 ( .A(n20006), .B(n19987), .Z(c[1856]) );
  NANDN U20958 ( .A(n19989), .B(n19988), .Z(n19993) );
  NAND U20959 ( .A(n19991), .B(n19990), .Z(n19992) );
  NAND U20960 ( .A(n19993), .B(n19992), .Z(n20012) );
  AND U20961 ( .A(b[2]), .B(a[835]), .Z(n20018) );
  AND U20962 ( .A(a[836]), .B(b[1]), .Z(n20016) );
  AND U20963 ( .A(a[834]), .B(b[3]), .Z(n20015) );
  XOR U20964 ( .A(n20016), .B(n20015), .Z(n20017) );
  XOR U20965 ( .A(n20018), .B(n20017), .Z(n20021) );
  NAND U20966 ( .A(b[0]), .B(a[837]), .Z(n20022) );
  XOR U20967 ( .A(n20021), .B(n20022), .Z(n20024) );
  OR U20968 ( .A(n19995), .B(n19994), .Z(n19999) );
  NANDN U20969 ( .A(n19997), .B(n19996), .Z(n19998) );
  NAND U20970 ( .A(n19999), .B(n19998), .Z(n20023) );
  XNOR U20971 ( .A(n20024), .B(n20023), .Z(n20009) );
  NANDN U20972 ( .A(n20001), .B(n20000), .Z(n20005) );
  OR U20973 ( .A(n20003), .B(n20002), .Z(n20004) );
  NAND U20974 ( .A(n20005), .B(n20004), .Z(n20010) );
  XNOR U20975 ( .A(n20009), .B(n20010), .Z(n20011) );
  XOR U20976 ( .A(n20012), .B(n20011), .Z(n20028) );
  XOR U20977 ( .A(sreg[1857]), .B(n20027), .Z(n20008) );
  XOR U20978 ( .A(n20028), .B(n20008), .Z(c[1857]) );
  NANDN U20979 ( .A(n20010), .B(n20009), .Z(n20014) );
  NAND U20980 ( .A(n20012), .B(n20011), .Z(n20013) );
  NAND U20981 ( .A(n20014), .B(n20013), .Z(n20035) );
  AND U20982 ( .A(b[2]), .B(a[836]), .Z(n20041) );
  AND U20983 ( .A(a[837]), .B(b[1]), .Z(n20039) );
  AND U20984 ( .A(a[835]), .B(b[3]), .Z(n20038) );
  XOR U20985 ( .A(n20039), .B(n20038), .Z(n20040) );
  XOR U20986 ( .A(n20041), .B(n20040), .Z(n20044) );
  NAND U20987 ( .A(b[0]), .B(a[838]), .Z(n20045) );
  XOR U20988 ( .A(n20044), .B(n20045), .Z(n20047) );
  OR U20989 ( .A(n20016), .B(n20015), .Z(n20020) );
  NANDN U20990 ( .A(n20018), .B(n20017), .Z(n20019) );
  NAND U20991 ( .A(n20020), .B(n20019), .Z(n20046) );
  XNOR U20992 ( .A(n20047), .B(n20046), .Z(n20032) );
  NANDN U20993 ( .A(n20022), .B(n20021), .Z(n20026) );
  OR U20994 ( .A(n20024), .B(n20023), .Z(n20025) );
  NAND U20995 ( .A(n20026), .B(n20025), .Z(n20033) );
  XNOR U20996 ( .A(n20032), .B(n20033), .Z(n20034) );
  XNOR U20997 ( .A(n20035), .B(n20034), .Z(n20031) );
  XOR U20998 ( .A(n20030), .B(sreg[1858]), .Z(n20029) );
  XOR U20999 ( .A(n20031), .B(n20029), .Z(c[1858]) );
  NANDN U21000 ( .A(n20033), .B(n20032), .Z(n20037) );
  NAND U21001 ( .A(n20035), .B(n20034), .Z(n20036) );
  NAND U21002 ( .A(n20037), .B(n20036), .Z(n20053) );
  AND U21003 ( .A(b[2]), .B(a[837]), .Z(n20059) );
  AND U21004 ( .A(a[838]), .B(b[1]), .Z(n20057) );
  AND U21005 ( .A(a[836]), .B(b[3]), .Z(n20056) );
  XOR U21006 ( .A(n20057), .B(n20056), .Z(n20058) );
  XOR U21007 ( .A(n20059), .B(n20058), .Z(n20062) );
  NAND U21008 ( .A(b[0]), .B(a[839]), .Z(n20063) );
  XOR U21009 ( .A(n20062), .B(n20063), .Z(n20065) );
  OR U21010 ( .A(n20039), .B(n20038), .Z(n20043) );
  NANDN U21011 ( .A(n20041), .B(n20040), .Z(n20042) );
  NAND U21012 ( .A(n20043), .B(n20042), .Z(n20064) );
  XNOR U21013 ( .A(n20065), .B(n20064), .Z(n20050) );
  NANDN U21014 ( .A(n20045), .B(n20044), .Z(n20049) );
  OR U21015 ( .A(n20047), .B(n20046), .Z(n20048) );
  NAND U21016 ( .A(n20049), .B(n20048), .Z(n20051) );
  XNOR U21017 ( .A(n20050), .B(n20051), .Z(n20052) );
  XNOR U21018 ( .A(n20053), .B(n20052), .Z(n20068) );
  XNOR U21019 ( .A(n20068), .B(sreg[1859]), .Z(n20070) );
  XNOR U21020 ( .A(n20069), .B(n20070), .Z(c[1859]) );
  NANDN U21021 ( .A(n20051), .B(n20050), .Z(n20055) );
  NAND U21022 ( .A(n20053), .B(n20052), .Z(n20054) );
  NAND U21023 ( .A(n20055), .B(n20054), .Z(n20081) );
  AND U21024 ( .A(b[2]), .B(a[838]), .Z(n20087) );
  AND U21025 ( .A(a[839]), .B(b[1]), .Z(n20085) );
  AND U21026 ( .A(a[837]), .B(b[3]), .Z(n20084) );
  XOR U21027 ( .A(n20085), .B(n20084), .Z(n20086) );
  XOR U21028 ( .A(n20087), .B(n20086), .Z(n20090) );
  NAND U21029 ( .A(b[0]), .B(a[840]), .Z(n20091) );
  XOR U21030 ( .A(n20090), .B(n20091), .Z(n20093) );
  OR U21031 ( .A(n20057), .B(n20056), .Z(n20061) );
  NANDN U21032 ( .A(n20059), .B(n20058), .Z(n20060) );
  NAND U21033 ( .A(n20061), .B(n20060), .Z(n20092) );
  XNOR U21034 ( .A(n20093), .B(n20092), .Z(n20078) );
  NANDN U21035 ( .A(n20063), .B(n20062), .Z(n20067) );
  OR U21036 ( .A(n20065), .B(n20064), .Z(n20066) );
  NAND U21037 ( .A(n20067), .B(n20066), .Z(n20079) );
  XNOR U21038 ( .A(n20078), .B(n20079), .Z(n20080) );
  XNOR U21039 ( .A(n20081), .B(n20080), .Z(n20073) );
  XOR U21040 ( .A(sreg[1860]), .B(n20073), .Z(n20074) );
  NAND U21041 ( .A(n20068), .B(sreg[1859]), .Z(n20072) );
  NANDN U21042 ( .A(n20070), .B(n20069), .Z(n20071) );
  NAND U21043 ( .A(n20072), .B(n20071), .Z(n20075) );
  XOR U21044 ( .A(n20074), .B(n20075), .Z(c[1860]) );
  OR U21045 ( .A(n20073), .B(sreg[1860]), .Z(n20077) );
  NANDN U21046 ( .A(n20075), .B(n20074), .Z(n20076) );
  AND U21047 ( .A(n20077), .B(n20076), .Z(n20097) );
  NANDN U21048 ( .A(n20079), .B(n20078), .Z(n20083) );
  NAND U21049 ( .A(n20081), .B(n20080), .Z(n20082) );
  NAND U21050 ( .A(n20083), .B(n20082), .Z(n20102) );
  AND U21051 ( .A(b[2]), .B(a[839]), .Z(n20108) );
  AND U21052 ( .A(a[840]), .B(b[1]), .Z(n20106) );
  AND U21053 ( .A(a[838]), .B(b[3]), .Z(n20105) );
  XOR U21054 ( .A(n20106), .B(n20105), .Z(n20107) );
  XOR U21055 ( .A(n20108), .B(n20107), .Z(n20111) );
  NAND U21056 ( .A(b[0]), .B(a[841]), .Z(n20112) );
  XOR U21057 ( .A(n20111), .B(n20112), .Z(n20114) );
  OR U21058 ( .A(n20085), .B(n20084), .Z(n20089) );
  NANDN U21059 ( .A(n20087), .B(n20086), .Z(n20088) );
  NAND U21060 ( .A(n20089), .B(n20088), .Z(n20113) );
  XNOR U21061 ( .A(n20114), .B(n20113), .Z(n20099) );
  NANDN U21062 ( .A(n20091), .B(n20090), .Z(n20095) );
  OR U21063 ( .A(n20093), .B(n20092), .Z(n20094) );
  NAND U21064 ( .A(n20095), .B(n20094), .Z(n20100) );
  XNOR U21065 ( .A(n20099), .B(n20100), .Z(n20101) );
  XNOR U21066 ( .A(n20102), .B(n20101), .Z(n20098) );
  XOR U21067 ( .A(sreg[1861]), .B(n20098), .Z(n20096) );
  XOR U21068 ( .A(n20097), .B(n20096), .Z(c[1861]) );
  NANDN U21069 ( .A(n20100), .B(n20099), .Z(n20104) );
  NAND U21070 ( .A(n20102), .B(n20101), .Z(n20103) );
  NAND U21071 ( .A(n20104), .B(n20103), .Z(n20120) );
  AND U21072 ( .A(b[2]), .B(a[840]), .Z(n20126) );
  AND U21073 ( .A(a[841]), .B(b[1]), .Z(n20124) );
  AND U21074 ( .A(a[839]), .B(b[3]), .Z(n20123) );
  XOR U21075 ( .A(n20124), .B(n20123), .Z(n20125) );
  XOR U21076 ( .A(n20126), .B(n20125), .Z(n20129) );
  NAND U21077 ( .A(b[0]), .B(a[842]), .Z(n20130) );
  XOR U21078 ( .A(n20129), .B(n20130), .Z(n20132) );
  OR U21079 ( .A(n20106), .B(n20105), .Z(n20110) );
  NANDN U21080 ( .A(n20108), .B(n20107), .Z(n20109) );
  NAND U21081 ( .A(n20110), .B(n20109), .Z(n20131) );
  XNOR U21082 ( .A(n20132), .B(n20131), .Z(n20117) );
  NANDN U21083 ( .A(n20112), .B(n20111), .Z(n20116) );
  OR U21084 ( .A(n20114), .B(n20113), .Z(n20115) );
  NAND U21085 ( .A(n20116), .B(n20115), .Z(n20118) );
  XNOR U21086 ( .A(n20117), .B(n20118), .Z(n20119) );
  XOR U21087 ( .A(n20120), .B(n20119), .Z(n20135) );
  XOR U21088 ( .A(sreg[1862]), .B(n20135), .Z(n20137) );
  XNOR U21089 ( .A(n20136), .B(n20137), .Z(c[1862]) );
  NANDN U21090 ( .A(n20118), .B(n20117), .Z(n20122) );
  NAND U21091 ( .A(n20120), .B(n20119), .Z(n20121) );
  NAND U21092 ( .A(n20122), .B(n20121), .Z(n20158) );
  AND U21093 ( .A(b[2]), .B(a[841]), .Z(n20152) );
  AND U21094 ( .A(a[842]), .B(b[1]), .Z(n20150) );
  AND U21095 ( .A(a[840]), .B(b[3]), .Z(n20149) );
  XOR U21096 ( .A(n20150), .B(n20149), .Z(n20151) );
  XOR U21097 ( .A(n20152), .B(n20151), .Z(n20143) );
  NAND U21098 ( .A(b[0]), .B(a[843]), .Z(n20144) );
  XOR U21099 ( .A(n20143), .B(n20144), .Z(n20146) );
  OR U21100 ( .A(n20124), .B(n20123), .Z(n20128) );
  NANDN U21101 ( .A(n20126), .B(n20125), .Z(n20127) );
  NAND U21102 ( .A(n20128), .B(n20127), .Z(n20145) );
  XNOR U21103 ( .A(n20146), .B(n20145), .Z(n20155) );
  NANDN U21104 ( .A(n20130), .B(n20129), .Z(n20134) );
  OR U21105 ( .A(n20132), .B(n20131), .Z(n20133) );
  NAND U21106 ( .A(n20134), .B(n20133), .Z(n20156) );
  XNOR U21107 ( .A(n20155), .B(n20156), .Z(n20157) );
  XOR U21108 ( .A(n20158), .B(n20157), .Z(n20142) );
  NANDN U21109 ( .A(n20135), .B(sreg[1862]), .Z(n20139) );
  NANDN U21110 ( .A(n20137), .B(n20136), .Z(n20138) );
  NAND U21111 ( .A(n20139), .B(n20138), .Z(n20141) );
  XNOR U21112 ( .A(sreg[1863]), .B(n20141), .Z(n20140) );
  XOR U21113 ( .A(n20142), .B(n20140), .Z(c[1863]) );
  NANDN U21114 ( .A(n20144), .B(n20143), .Z(n20148) );
  OR U21115 ( .A(n20146), .B(n20145), .Z(n20147) );
  NAND U21116 ( .A(n20148), .B(n20147), .Z(n20161) );
  AND U21117 ( .A(b[2]), .B(a[842]), .Z(n20170) );
  AND U21118 ( .A(a[843]), .B(b[1]), .Z(n20168) );
  AND U21119 ( .A(a[841]), .B(b[3]), .Z(n20167) );
  XOR U21120 ( .A(n20168), .B(n20167), .Z(n20169) );
  XOR U21121 ( .A(n20170), .B(n20169), .Z(n20173) );
  NAND U21122 ( .A(b[0]), .B(a[844]), .Z(n20174) );
  XNOR U21123 ( .A(n20173), .B(n20174), .Z(n20175) );
  OR U21124 ( .A(n20150), .B(n20149), .Z(n20154) );
  NANDN U21125 ( .A(n20152), .B(n20151), .Z(n20153) );
  AND U21126 ( .A(n20154), .B(n20153), .Z(n20176) );
  XNOR U21127 ( .A(n20175), .B(n20176), .Z(n20162) );
  XNOR U21128 ( .A(n20161), .B(n20162), .Z(n20163) );
  NANDN U21129 ( .A(n20156), .B(n20155), .Z(n20160) );
  NAND U21130 ( .A(n20158), .B(n20157), .Z(n20159) );
  NAND U21131 ( .A(n20160), .B(n20159), .Z(n20164) );
  XNOR U21132 ( .A(n20163), .B(n20164), .Z(n20179) );
  XOR U21133 ( .A(sreg[1864]), .B(n20179), .Z(n20181) );
  XNOR U21134 ( .A(n20180), .B(n20181), .Z(c[1864]) );
  NANDN U21135 ( .A(n20162), .B(n20161), .Z(n20166) );
  NANDN U21136 ( .A(n20164), .B(n20163), .Z(n20165) );
  NAND U21137 ( .A(n20166), .B(n20165), .Z(n20190) );
  AND U21138 ( .A(b[2]), .B(a[843]), .Z(n20196) );
  AND U21139 ( .A(a[844]), .B(b[1]), .Z(n20194) );
  AND U21140 ( .A(a[842]), .B(b[3]), .Z(n20193) );
  XOR U21141 ( .A(n20194), .B(n20193), .Z(n20195) );
  XOR U21142 ( .A(n20196), .B(n20195), .Z(n20199) );
  NAND U21143 ( .A(b[0]), .B(a[845]), .Z(n20200) );
  XOR U21144 ( .A(n20199), .B(n20200), .Z(n20202) );
  OR U21145 ( .A(n20168), .B(n20167), .Z(n20172) );
  NANDN U21146 ( .A(n20170), .B(n20169), .Z(n20171) );
  NAND U21147 ( .A(n20172), .B(n20171), .Z(n20201) );
  XNOR U21148 ( .A(n20202), .B(n20201), .Z(n20187) );
  NANDN U21149 ( .A(n20174), .B(n20173), .Z(n20178) );
  NAND U21150 ( .A(n20176), .B(n20175), .Z(n20177) );
  NAND U21151 ( .A(n20178), .B(n20177), .Z(n20188) );
  XNOR U21152 ( .A(n20187), .B(n20188), .Z(n20189) );
  XOR U21153 ( .A(n20190), .B(n20189), .Z(n20186) );
  OR U21154 ( .A(n20179), .B(sreg[1864]), .Z(n20183) );
  NAND U21155 ( .A(n20181), .B(n20180), .Z(n20182) );
  AND U21156 ( .A(n20183), .B(n20182), .Z(n20185) );
  XNOR U21157 ( .A(sreg[1865]), .B(n20185), .Z(n20184) );
  XNOR U21158 ( .A(n20186), .B(n20184), .Z(c[1865]) );
  NANDN U21159 ( .A(n20188), .B(n20187), .Z(n20192) );
  NANDN U21160 ( .A(n20190), .B(n20189), .Z(n20191) );
  NAND U21161 ( .A(n20192), .B(n20191), .Z(n20208) );
  AND U21162 ( .A(b[2]), .B(a[844]), .Z(n20220) );
  AND U21163 ( .A(a[845]), .B(b[1]), .Z(n20218) );
  AND U21164 ( .A(a[843]), .B(b[3]), .Z(n20217) );
  XOR U21165 ( .A(n20218), .B(n20217), .Z(n20219) );
  XOR U21166 ( .A(n20220), .B(n20219), .Z(n20211) );
  NAND U21167 ( .A(b[0]), .B(a[846]), .Z(n20212) );
  XOR U21168 ( .A(n20211), .B(n20212), .Z(n20214) );
  OR U21169 ( .A(n20194), .B(n20193), .Z(n20198) );
  NANDN U21170 ( .A(n20196), .B(n20195), .Z(n20197) );
  NAND U21171 ( .A(n20198), .B(n20197), .Z(n20213) );
  XNOR U21172 ( .A(n20214), .B(n20213), .Z(n20205) );
  NANDN U21173 ( .A(n20200), .B(n20199), .Z(n20204) );
  OR U21174 ( .A(n20202), .B(n20201), .Z(n20203) );
  NAND U21175 ( .A(n20204), .B(n20203), .Z(n20206) );
  XNOR U21176 ( .A(n20205), .B(n20206), .Z(n20207) );
  XNOR U21177 ( .A(n20208), .B(n20207), .Z(n20223) );
  XOR U21178 ( .A(sreg[1866]), .B(n20223), .Z(n20225) );
  XNOR U21179 ( .A(n20224), .B(n20225), .Z(c[1866]) );
  NANDN U21180 ( .A(n20206), .B(n20205), .Z(n20210) );
  NAND U21181 ( .A(n20208), .B(n20207), .Z(n20209) );
  NAND U21182 ( .A(n20210), .B(n20209), .Z(n20246) );
  NANDN U21183 ( .A(n20212), .B(n20211), .Z(n20216) );
  OR U21184 ( .A(n20214), .B(n20213), .Z(n20215) );
  NAND U21185 ( .A(n20216), .B(n20215), .Z(n20243) );
  AND U21186 ( .A(b[2]), .B(a[845]), .Z(n20234) );
  AND U21187 ( .A(a[846]), .B(b[1]), .Z(n20232) );
  AND U21188 ( .A(a[844]), .B(b[3]), .Z(n20231) );
  XOR U21189 ( .A(n20232), .B(n20231), .Z(n20233) );
  XOR U21190 ( .A(n20234), .B(n20233), .Z(n20237) );
  NAND U21191 ( .A(b[0]), .B(a[847]), .Z(n20238) );
  XNOR U21192 ( .A(n20237), .B(n20238), .Z(n20239) );
  OR U21193 ( .A(n20218), .B(n20217), .Z(n20222) );
  NANDN U21194 ( .A(n20220), .B(n20219), .Z(n20221) );
  AND U21195 ( .A(n20222), .B(n20221), .Z(n20240) );
  XNOR U21196 ( .A(n20239), .B(n20240), .Z(n20244) );
  XNOR U21197 ( .A(n20243), .B(n20244), .Z(n20245) );
  XOR U21198 ( .A(n20246), .B(n20245), .Z(n20230) );
  OR U21199 ( .A(n20223), .B(sreg[1866]), .Z(n20227) );
  NAND U21200 ( .A(n20225), .B(n20224), .Z(n20226) );
  AND U21201 ( .A(n20227), .B(n20226), .Z(n20229) );
  XOR U21202 ( .A(sreg[1867]), .B(n20229), .Z(n20228) );
  XNOR U21203 ( .A(n20230), .B(n20228), .Z(c[1867]) );
  AND U21204 ( .A(b[2]), .B(a[846]), .Z(n20258) );
  AND U21205 ( .A(a[847]), .B(b[1]), .Z(n20256) );
  AND U21206 ( .A(a[845]), .B(b[3]), .Z(n20255) );
  XOR U21207 ( .A(n20256), .B(n20255), .Z(n20257) );
  XOR U21208 ( .A(n20258), .B(n20257), .Z(n20261) );
  NAND U21209 ( .A(b[0]), .B(a[848]), .Z(n20262) );
  XOR U21210 ( .A(n20261), .B(n20262), .Z(n20264) );
  OR U21211 ( .A(n20232), .B(n20231), .Z(n20236) );
  NANDN U21212 ( .A(n20234), .B(n20233), .Z(n20235) );
  NAND U21213 ( .A(n20236), .B(n20235), .Z(n20263) );
  XNOR U21214 ( .A(n20264), .B(n20263), .Z(n20249) );
  NANDN U21215 ( .A(n20238), .B(n20237), .Z(n20242) );
  NAND U21216 ( .A(n20240), .B(n20239), .Z(n20241) );
  NAND U21217 ( .A(n20242), .B(n20241), .Z(n20250) );
  XNOR U21218 ( .A(n20249), .B(n20250), .Z(n20251) );
  NANDN U21219 ( .A(n20244), .B(n20243), .Z(n20248) );
  NANDN U21220 ( .A(n20246), .B(n20245), .Z(n20247) );
  NAND U21221 ( .A(n20248), .B(n20247), .Z(n20252) );
  XOR U21222 ( .A(n20251), .B(n20252), .Z(n20267) );
  XNOR U21223 ( .A(n20267), .B(sreg[1868]), .Z(n20269) );
  XNOR U21224 ( .A(n20268), .B(n20269), .Z(c[1868]) );
  NANDN U21225 ( .A(n20250), .B(n20249), .Z(n20254) );
  NANDN U21226 ( .A(n20252), .B(n20251), .Z(n20253) );
  NAND U21227 ( .A(n20254), .B(n20253), .Z(n20288) );
  AND U21228 ( .A(b[2]), .B(a[847]), .Z(n20282) );
  AND U21229 ( .A(a[848]), .B(b[1]), .Z(n20280) );
  AND U21230 ( .A(a[846]), .B(b[3]), .Z(n20279) );
  XOR U21231 ( .A(n20280), .B(n20279), .Z(n20281) );
  XOR U21232 ( .A(n20282), .B(n20281), .Z(n20273) );
  NAND U21233 ( .A(b[0]), .B(a[849]), .Z(n20274) );
  XOR U21234 ( .A(n20273), .B(n20274), .Z(n20276) );
  OR U21235 ( .A(n20256), .B(n20255), .Z(n20260) );
  NANDN U21236 ( .A(n20258), .B(n20257), .Z(n20259) );
  NAND U21237 ( .A(n20260), .B(n20259), .Z(n20275) );
  XNOR U21238 ( .A(n20276), .B(n20275), .Z(n20285) );
  NANDN U21239 ( .A(n20262), .B(n20261), .Z(n20266) );
  OR U21240 ( .A(n20264), .B(n20263), .Z(n20265) );
  NAND U21241 ( .A(n20266), .B(n20265), .Z(n20286) );
  XNOR U21242 ( .A(n20285), .B(n20286), .Z(n20287) );
  XNOR U21243 ( .A(n20288), .B(n20287), .Z(n20292) );
  NAND U21244 ( .A(n20267), .B(sreg[1868]), .Z(n20271) );
  NANDN U21245 ( .A(n20269), .B(n20268), .Z(n20270) );
  AND U21246 ( .A(n20271), .B(n20270), .Z(n20291) );
  XNOR U21247 ( .A(n20291), .B(sreg[1869]), .Z(n20272) );
  XOR U21248 ( .A(n20292), .B(n20272), .Z(c[1869]) );
  NANDN U21249 ( .A(n20274), .B(n20273), .Z(n20278) );
  OR U21250 ( .A(n20276), .B(n20275), .Z(n20277) );
  NAND U21251 ( .A(n20278), .B(n20277), .Z(n20296) );
  AND U21252 ( .A(b[2]), .B(a[848]), .Z(n20305) );
  AND U21253 ( .A(a[849]), .B(b[1]), .Z(n20303) );
  AND U21254 ( .A(a[847]), .B(b[3]), .Z(n20302) );
  XOR U21255 ( .A(n20303), .B(n20302), .Z(n20304) );
  XOR U21256 ( .A(n20305), .B(n20304), .Z(n20308) );
  NAND U21257 ( .A(b[0]), .B(a[850]), .Z(n20309) );
  XNOR U21258 ( .A(n20308), .B(n20309), .Z(n20310) );
  OR U21259 ( .A(n20280), .B(n20279), .Z(n20284) );
  NANDN U21260 ( .A(n20282), .B(n20281), .Z(n20283) );
  AND U21261 ( .A(n20284), .B(n20283), .Z(n20311) );
  XNOR U21262 ( .A(n20310), .B(n20311), .Z(n20297) );
  XNOR U21263 ( .A(n20296), .B(n20297), .Z(n20298) );
  NANDN U21264 ( .A(n20286), .B(n20285), .Z(n20290) );
  NAND U21265 ( .A(n20288), .B(n20287), .Z(n20289) );
  NAND U21266 ( .A(n20290), .B(n20289), .Z(n20299) );
  XOR U21267 ( .A(n20298), .B(n20299), .Z(n20295) );
  XOR U21268 ( .A(n20294), .B(sreg[1870]), .Z(n20293) );
  XNOR U21269 ( .A(n20295), .B(n20293), .Z(c[1870]) );
  NANDN U21270 ( .A(n20297), .B(n20296), .Z(n20301) );
  NANDN U21271 ( .A(n20299), .B(n20298), .Z(n20300) );
  NAND U21272 ( .A(n20301), .B(n20300), .Z(n20317) );
  AND U21273 ( .A(b[2]), .B(a[849]), .Z(n20323) );
  AND U21274 ( .A(a[850]), .B(b[1]), .Z(n20321) );
  AND U21275 ( .A(a[848]), .B(b[3]), .Z(n20320) );
  XOR U21276 ( .A(n20321), .B(n20320), .Z(n20322) );
  XOR U21277 ( .A(n20323), .B(n20322), .Z(n20326) );
  NAND U21278 ( .A(b[0]), .B(a[851]), .Z(n20327) );
  XOR U21279 ( .A(n20326), .B(n20327), .Z(n20329) );
  OR U21280 ( .A(n20303), .B(n20302), .Z(n20307) );
  NANDN U21281 ( .A(n20305), .B(n20304), .Z(n20306) );
  NAND U21282 ( .A(n20307), .B(n20306), .Z(n20328) );
  XNOR U21283 ( .A(n20329), .B(n20328), .Z(n20314) );
  NANDN U21284 ( .A(n20309), .B(n20308), .Z(n20313) );
  NAND U21285 ( .A(n20311), .B(n20310), .Z(n20312) );
  NAND U21286 ( .A(n20313), .B(n20312), .Z(n20315) );
  XNOR U21287 ( .A(n20314), .B(n20315), .Z(n20316) );
  XOR U21288 ( .A(n20317), .B(n20316), .Z(n20332) );
  XNOR U21289 ( .A(n20332), .B(sreg[1871]), .Z(n20334) );
  XNOR U21290 ( .A(n20333), .B(n20334), .Z(c[1871]) );
  NANDN U21291 ( .A(n20315), .B(n20314), .Z(n20319) );
  NANDN U21292 ( .A(n20317), .B(n20316), .Z(n20318) );
  NAND U21293 ( .A(n20319), .B(n20318), .Z(n20355) );
  AND U21294 ( .A(b[2]), .B(a[850]), .Z(n20349) );
  AND U21295 ( .A(a[851]), .B(b[1]), .Z(n20347) );
  AND U21296 ( .A(a[849]), .B(b[3]), .Z(n20346) );
  XOR U21297 ( .A(n20347), .B(n20346), .Z(n20348) );
  XOR U21298 ( .A(n20349), .B(n20348), .Z(n20340) );
  NAND U21299 ( .A(b[0]), .B(a[852]), .Z(n20341) );
  XOR U21300 ( .A(n20340), .B(n20341), .Z(n20343) );
  OR U21301 ( .A(n20321), .B(n20320), .Z(n20325) );
  NANDN U21302 ( .A(n20323), .B(n20322), .Z(n20324) );
  NAND U21303 ( .A(n20325), .B(n20324), .Z(n20342) );
  XNOR U21304 ( .A(n20343), .B(n20342), .Z(n20352) );
  NANDN U21305 ( .A(n20327), .B(n20326), .Z(n20331) );
  OR U21306 ( .A(n20329), .B(n20328), .Z(n20330) );
  NAND U21307 ( .A(n20331), .B(n20330), .Z(n20353) );
  XNOR U21308 ( .A(n20352), .B(n20353), .Z(n20354) );
  XOR U21309 ( .A(n20355), .B(n20354), .Z(n20339) );
  NAND U21310 ( .A(n20332), .B(sreg[1871]), .Z(n20336) );
  NANDN U21311 ( .A(n20334), .B(n20333), .Z(n20335) );
  NAND U21312 ( .A(n20336), .B(n20335), .Z(n20338) );
  XNOR U21313 ( .A(sreg[1872]), .B(n20338), .Z(n20337) );
  XOR U21314 ( .A(n20339), .B(n20337), .Z(c[1872]) );
  NANDN U21315 ( .A(n20341), .B(n20340), .Z(n20345) );
  OR U21316 ( .A(n20343), .B(n20342), .Z(n20344) );
  NAND U21317 ( .A(n20345), .B(n20344), .Z(n20358) );
  AND U21318 ( .A(b[2]), .B(a[851]), .Z(n20367) );
  AND U21319 ( .A(a[852]), .B(b[1]), .Z(n20365) );
  AND U21320 ( .A(a[850]), .B(b[3]), .Z(n20364) );
  XOR U21321 ( .A(n20365), .B(n20364), .Z(n20366) );
  XOR U21322 ( .A(n20367), .B(n20366), .Z(n20370) );
  NAND U21323 ( .A(b[0]), .B(a[853]), .Z(n20371) );
  XNOR U21324 ( .A(n20370), .B(n20371), .Z(n20372) );
  OR U21325 ( .A(n20347), .B(n20346), .Z(n20351) );
  NANDN U21326 ( .A(n20349), .B(n20348), .Z(n20350) );
  AND U21327 ( .A(n20351), .B(n20350), .Z(n20373) );
  XNOR U21328 ( .A(n20372), .B(n20373), .Z(n20359) );
  XNOR U21329 ( .A(n20358), .B(n20359), .Z(n20360) );
  NANDN U21330 ( .A(n20353), .B(n20352), .Z(n20357) );
  NAND U21331 ( .A(n20355), .B(n20354), .Z(n20356) );
  NAND U21332 ( .A(n20357), .B(n20356), .Z(n20361) );
  XOR U21333 ( .A(n20360), .B(n20361), .Z(n20376) );
  XNOR U21334 ( .A(sreg[1873]), .B(n20376), .Z(n20377) );
  XNOR U21335 ( .A(n20378), .B(n20377), .Z(c[1873]) );
  NANDN U21336 ( .A(n20359), .B(n20358), .Z(n20363) );
  NANDN U21337 ( .A(n20361), .B(n20360), .Z(n20362) );
  NAND U21338 ( .A(n20363), .B(n20362), .Z(n20389) );
  AND U21339 ( .A(b[2]), .B(a[852]), .Z(n20395) );
  AND U21340 ( .A(a[853]), .B(b[1]), .Z(n20393) );
  AND U21341 ( .A(a[851]), .B(b[3]), .Z(n20392) );
  XOR U21342 ( .A(n20393), .B(n20392), .Z(n20394) );
  XOR U21343 ( .A(n20395), .B(n20394), .Z(n20398) );
  NAND U21344 ( .A(b[0]), .B(a[854]), .Z(n20399) );
  XOR U21345 ( .A(n20398), .B(n20399), .Z(n20401) );
  OR U21346 ( .A(n20365), .B(n20364), .Z(n20369) );
  NANDN U21347 ( .A(n20367), .B(n20366), .Z(n20368) );
  NAND U21348 ( .A(n20369), .B(n20368), .Z(n20400) );
  XNOR U21349 ( .A(n20401), .B(n20400), .Z(n20386) );
  NANDN U21350 ( .A(n20371), .B(n20370), .Z(n20375) );
  NAND U21351 ( .A(n20373), .B(n20372), .Z(n20374) );
  NAND U21352 ( .A(n20375), .B(n20374), .Z(n20387) );
  XNOR U21353 ( .A(n20386), .B(n20387), .Z(n20388) );
  XNOR U21354 ( .A(n20389), .B(n20388), .Z(n20381) );
  XOR U21355 ( .A(sreg[1874]), .B(n20381), .Z(n20383) );
  NANDN U21356 ( .A(sreg[1873]), .B(n20376), .Z(n20380) );
  NAND U21357 ( .A(n20378), .B(n20377), .Z(n20379) );
  AND U21358 ( .A(n20380), .B(n20379), .Z(n20382) );
  XNOR U21359 ( .A(n20383), .B(n20382), .Z(c[1874]) );
  NANDN U21360 ( .A(sreg[1874]), .B(n20381), .Z(n20385) );
  OR U21361 ( .A(n20383), .B(n20382), .Z(n20384) );
  AND U21362 ( .A(n20385), .B(n20384), .Z(n20405) );
  NANDN U21363 ( .A(n20387), .B(n20386), .Z(n20391) );
  NANDN U21364 ( .A(n20389), .B(n20388), .Z(n20390) );
  NAND U21365 ( .A(n20391), .B(n20390), .Z(n20422) );
  AND U21366 ( .A(b[2]), .B(a[853]), .Z(n20416) );
  AND U21367 ( .A(a[854]), .B(b[1]), .Z(n20414) );
  AND U21368 ( .A(a[852]), .B(b[3]), .Z(n20413) );
  XOR U21369 ( .A(n20414), .B(n20413), .Z(n20415) );
  XOR U21370 ( .A(n20416), .B(n20415), .Z(n20407) );
  NAND U21371 ( .A(b[0]), .B(a[855]), .Z(n20408) );
  XOR U21372 ( .A(n20407), .B(n20408), .Z(n20410) );
  OR U21373 ( .A(n20393), .B(n20392), .Z(n20397) );
  NANDN U21374 ( .A(n20395), .B(n20394), .Z(n20396) );
  NAND U21375 ( .A(n20397), .B(n20396), .Z(n20409) );
  XNOR U21376 ( .A(n20410), .B(n20409), .Z(n20419) );
  NANDN U21377 ( .A(n20399), .B(n20398), .Z(n20403) );
  OR U21378 ( .A(n20401), .B(n20400), .Z(n20402) );
  NAND U21379 ( .A(n20403), .B(n20402), .Z(n20420) );
  XNOR U21380 ( .A(n20419), .B(n20420), .Z(n20421) );
  XNOR U21381 ( .A(n20422), .B(n20421), .Z(n20406) );
  XOR U21382 ( .A(sreg[1875]), .B(n20406), .Z(n20404) );
  XOR U21383 ( .A(n20405), .B(n20404), .Z(c[1875]) );
  NANDN U21384 ( .A(n20408), .B(n20407), .Z(n20412) );
  OR U21385 ( .A(n20410), .B(n20409), .Z(n20411) );
  NAND U21386 ( .A(n20412), .B(n20411), .Z(n20425) );
  AND U21387 ( .A(b[2]), .B(a[854]), .Z(n20434) );
  AND U21388 ( .A(a[855]), .B(b[1]), .Z(n20432) );
  AND U21389 ( .A(a[853]), .B(b[3]), .Z(n20431) );
  XOR U21390 ( .A(n20432), .B(n20431), .Z(n20433) );
  XOR U21391 ( .A(n20434), .B(n20433), .Z(n20437) );
  NAND U21392 ( .A(b[0]), .B(a[856]), .Z(n20438) );
  XNOR U21393 ( .A(n20437), .B(n20438), .Z(n20439) );
  OR U21394 ( .A(n20414), .B(n20413), .Z(n20418) );
  NANDN U21395 ( .A(n20416), .B(n20415), .Z(n20417) );
  AND U21396 ( .A(n20418), .B(n20417), .Z(n20440) );
  XNOR U21397 ( .A(n20439), .B(n20440), .Z(n20426) );
  XNOR U21398 ( .A(n20425), .B(n20426), .Z(n20427) );
  NANDN U21399 ( .A(n20420), .B(n20419), .Z(n20424) );
  NAND U21400 ( .A(n20422), .B(n20421), .Z(n20423) );
  AND U21401 ( .A(n20424), .B(n20423), .Z(n20428) );
  XNOR U21402 ( .A(n20427), .B(n20428), .Z(n20443) );
  XOR U21403 ( .A(n20443), .B(sreg[1876]), .Z(n20445) );
  XNOR U21404 ( .A(n20444), .B(n20445), .Z(c[1876]) );
  NANDN U21405 ( .A(n20426), .B(n20425), .Z(n20430) );
  NAND U21406 ( .A(n20428), .B(n20427), .Z(n20429) );
  NAND U21407 ( .A(n20430), .B(n20429), .Z(n20456) );
  AND U21408 ( .A(b[2]), .B(a[855]), .Z(n20462) );
  AND U21409 ( .A(a[856]), .B(b[1]), .Z(n20460) );
  AND U21410 ( .A(a[854]), .B(b[3]), .Z(n20459) );
  XOR U21411 ( .A(n20460), .B(n20459), .Z(n20461) );
  XOR U21412 ( .A(n20462), .B(n20461), .Z(n20465) );
  NAND U21413 ( .A(b[0]), .B(a[857]), .Z(n20466) );
  XOR U21414 ( .A(n20465), .B(n20466), .Z(n20468) );
  OR U21415 ( .A(n20432), .B(n20431), .Z(n20436) );
  NANDN U21416 ( .A(n20434), .B(n20433), .Z(n20435) );
  NAND U21417 ( .A(n20436), .B(n20435), .Z(n20467) );
  XNOR U21418 ( .A(n20468), .B(n20467), .Z(n20453) );
  NANDN U21419 ( .A(n20438), .B(n20437), .Z(n20442) );
  NAND U21420 ( .A(n20440), .B(n20439), .Z(n20441) );
  NAND U21421 ( .A(n20442), .B(n20441), .Z(n20454) );
  XNOR U21422 ( .A(n20453), .B(n20454), .Z(n20455) );
  XNOR U21423 ( .A(n20456), .B(n20455), .Z(n20448) );
  XOR U21424 ( .A(sreg[1877]), .B(n20448), .Z(n20450) );
  NANDN U21425 ( .A(n20443), .B(sreg[1876]), .Z(n20447) );
  NANDN U21426 ( .A(n20445), .B(n20444), .Z(n20446) );
  NAND U21427 ( .A(n20447), .B(n20446), .Z(n20449) );
  XNOR U21428 ( .A(n20450), .B(n20449), .Z(c[1877]) );
  NANDN U21429 ( .A(sreg[1877]), .B(n20448), .Z(n20452) );
  OR U21430 ( .A(n20450), .B(n20449), .Z(n20451) );
  AND U21431 ( .A(n20452), .B(n20451), .Z(n20490) );
  NANDN U21432 ( .A(n20454), .B(n20453), .Z(n20458) );
  NANDN U21433 ( .A(n20456), .B(n20455), .Z(n20457) );
  NAND U21434 ( .A(n20458), .B(n20457), .Z(n20487) );
  AND U21435 ( .A(b[2]), .B(a[856]), .Z(n20481) );
  AND U21436 ( .A(a[857]), .B(b[1]), .Z(n20479) );
  AND U21437 ( .A(a[855]), .B(b[3]), .Z(n20478) );
  XOR U21438 ( .A(n20479), .B(n20478), .Z(n20480) );
  XOR U21439 ( .A(n20481), .B(n20480), .Z(n20472) );
  NAND U21440 ( .A(b[0]), .B(a[858]), .Z(n20473) );
  XOR U21441 ( .A(n20472), .B(n20473), .Z(n20475) );
  OR U21442 ( .A(n20460), .B(n20459), .Z(n20464) );
  NANDN U21443 ( .A(n20462), .B(n20461), .Z(n20463) );
  NAND U21444 ( .A(n20464), .B(n20463), .Z(n20474) );
  XNOR U21445 ( .A(n20475), .B(n20474), .Z(n20484) );
  NANDN U21446 ( .A(n20466), .B(n20465), .Z(n20470) );
  OR U21447 ( .A(n20468), .B(n20467), .Z(n20469) );
  NAND U21448 ( .A(n20470), .B(n20469), .Z(n20485) );
  XNOR U21449 ( .A(n20484), .B(n20485), .Z(n20486) );
  XNOR U21450 ( .A(n20487), .B(n20486), .Z(n20491) );
  XOR U21451 ( .A(sreg[1878]), .B(n20491), .Z(n20471) );
  XOR U21452 ( .A(n20490), .B(n20471), .Z(c[1878]) );
  NANDN U21453 ( .A(n20473), .B(n20472), .Z(n20477) );
  OR U21454 ( .A(n20475), .B(n20474), .Z(n20476) );
  NAND U21455 ( .A(n20477), .B(n20476), .Z(n20495) );
  AND U21456 ( .A(b[2]), .B(a[857]), .Z(n20504) );
  AND U21457 ( .A(a[858]), .B(b[1]), .Z(n20502) );
  AND U21458 ( .A(a[856]), .B(b[3]), .Z(n20501) );
  XOR U21459 ( .A(n20502), .B(n20501), .Z(n20503) );
  XOR U21460 ( .A(n20504), .B(n20503), .Z(n20507) );
  NAND U21461 ( .A(b[0]), .B(a[859]), .Z(n20508) );
  XNOR U21462 ( .A(n20507), .B(n20508), .Z(n20509) );
  OR U21463 ( .A(n20479), .B(n20478), .Z(n20483) );
  NANDN U21464 ( .A(n20481), .B(n20480), .Z(n20482) );
  AND U21465 ( .A(n20483), .B(n20482), .Z(n20510) );
  XNOR U21466 ( .A(n20509), .B(n20510), .Z(n20496) );
  XNOR U21467 ( .A(n20495), .B(n20496), .Z(n20497) );
  NANDN U21468 ( .A(n20485), .B(n20484), .Z(n20489) );
  NAND U21469 ( .A(n20487), .B(n20486), .Z(n20488) );
  NAND U21470 ( .A(n20489), .B(n20488), .Z(n20498) );
  XOR U21471 ( .A(n20497), .B(n20498), .Z(n20494) );
  XOR U21472 ( .A(n20493), .B(sreg[1879]), .Z(n20492) );
  XNOR U21473 ( .A(n20494), .B(n20492), .Z(c[1879]) );
  NANDN U21474 ( .A(n20496), .B(n20495), .Z(n20500) );
  NANDN U21475 ( .A(n20498), .B(n20497), .Z(n20499) );
  NAND U21476 ( .A(n20500), .B(n20499), .Z(n20516) );
  AND U21477 ( .A(b[2]), .B(a[858]), .Z(n20522) );
  AND U21478 ( .A(a[859]), .B(b[1]), .Z(n20520) );
  AND U21479 ( .A(a[857]), .B(b[3]), .Z(n20519) );
  XOR U21480 ( .A(n20520), .B(n20519), .Z(n20521) );
  XOR U21481 ( .A(n20522), .B(n20521), .Z(n20525) );
  NAND U21482 ( .A(b[0]), .B(a[860]), .Z(n20526) );
  XOR U21483 ( .A(n20525), .B(n20526), .Z(n20528) );
  OR U21484 ( .A(n20502), .B(n20501), .Z(n20506) );
  NANDN U21485 ( .A(n20504), .B(n20503), .Z(n20505) );
  NAND U21486 ( .A(n20506), .B(n20505), .Z(n20527) );
  XNOR U21487 ( .A(n20528), .B(n20527), .Z(n20513) );
  NANDN U21488 ( .A(n20508), .B(n20507), .Z(n20512) );
  NAND U21489 ( .A(n20510), .B(n20509), .Z(n20511) );
  NAND U21490 ( .A(n20512), .B(n20511), .Z(n20514) );
  XNOR U21491 ( .A(n20513), .B(n20514), .Z(n20515) );
  XOR U21492 ( .A(n20516), .B(n20515), .Z(n20531) );
  XNOR U21493 ( .A(n20531), .B(sreg[1880]), .Z(n20533) );
  XNOR U21494 ( .A(n20532), .B(n20533), .Z(c[1880]) );
  NANDN U21495 ( .A(n20514), .B(n20513), .Z(n20518) );
  NANDN U21496 ( .A(n20516), .B(n20515), .Z(n20517) );
  NAND U21497 ( .A(n20518), .B(n20517), .Z(n20544) );
  AND U21498 ( .A(b[2]), .B(a[859]), .Z(n20550) );
  AND U21499 ( .A(a[860]), .B(b[1]), .Z(n20548) );
  AND U21500 ( .A(a[858]), .B(b[3]), .Z(n20547) );
  XOR U21501 ( .A(n20548), .B(n20547), .Z(n20549) );
  XOR U21502 ( .A(n20550), .B(n20549), .Z(n20553) );
  NAND U21503 ( .A(b[0]), .B(a[861]), .Z(n20554) );
  XOR U21504 ( .A(n20553), .B(n20554), .Z(n20556) );
  OR U21505 ( .A(n20520), .B(n20519), .Z(n20524) );
  NANDN U21506 ( .A(n20522), .B(n20521), .Z(n20523) );
  NAND U21507 ( .A(n20524), .B(n20523), .Z(n20555) );
  XNOR U21508 ( .A(n20556), .B(n20555), .Z(n20541) );
  NANDN U21509 ( .A(n20526), .B(n20525), .Z(n20530) );
  OR U21510 ( .A(n20528), .B(n20527), .Z(n20529) );
  NAND U21511 ( .A(n20530), .B(n20529), .Z(n20542) );
  XNOR U21512 ( .A(n20541), .B(n20542), .Z(n20543) );
  XNOR U21513 ( .A(n20544), .B(n20543), .Z(n20536) );
  XNOR U21514 ( .A(n20536), .B(sreg[1881]), .Z(n20538) );
  NAND U21515 ( .A(n20531), .B(sreg[1880]), .Z(n20535) );
  NANDN U21516 ( .A(n20533), .B(n20532), .Z(n20534) );
  AND U21517 ( .A(n20535), .B(n20534), .Z(n20537) );
  XOR U21518 ( .A(n20538), .B(n20537), .Z(c[1881]) );
  NAND U21519 ( .A(n20536), .B(sreg[1881]), .Z(n20540) );
  OR U21520 ( .A(n20538), .B(n20537), .Z(n20539) );
  NAND U21521 ( .A(n20540), .B(n20539), .Z(n20561) );
  NANDN U21522 ( .A(n20542), .B(n20541), .Z(n20546) );
  NAND U21523 ( .A(n20544), .B(n20543), .Z(n20545) );
  AND U21524 ( .A(n20546), .B(n20545), .Z(n20565) );
  AND U21525 ( .A(b[2]), .B(a[860]), .Z(n20569) );
  AND U21526 ( .A(a[861]), .B(b[1]), .Z(n20567) );
  AND U21527 ( .A(a[859]), .B(b[3]), .Z(n20566) );
  XOR U21528 ( .A(n20567), .B(n20566), .Z(n20568) );
  XOR U21529 ( .A(n20569), .B(n20568), .Z(n20572) );
  NAND U21530 ( .A(b[0]), .B(a[862]), .Z(n20573) );
  XOR U21531 ( .A(n20572), .B(n20573), .Z(n20574) );
  OR U21532 ( .A(n20548), .B(n20547), .Z(n20552) );
  NANDN U21533 ( .A(n20550), .B(n20549), .Z(n20551) );
  AND U21534 ( .A(n20552), .B(n20551), .Z(n20575) );
  XOR U21535 ( .A(n20574), .B(n20575), .Z(n20563) );
  NANDN U21536 ( .A(n20554), .B(n20553), .Z(n20558) );
  OR U21537 ( .A(n20556), .B(n20555), .Z(n20557) );
  AND U21538 ( .A(n20558), .B(n20557), .Z(n20564) );
  XOR U21539 ( .A(n20563), .B(n20564), .Z(n20559) );
  XNOR U21540 ( .A(n20565), .B(n20559), .Z(n20562) );
  XOR U21541 ( .A(sreg[1882]), .B(n20562), .Z(n20560) );
  XNOR U21542 ( .A(n20561), .B(n20560), .Z(c[1882]) );
  AND U21543 ( .A(b[2]), .B(a[861]), .Z(n20585) );
  AND U21544 ( .A(a[862]), .B(b[1]), .Z(n20583) );
  AND U21545 ( .A(a[860]), .B(b[3]), .Z(n20582) );
  XOR U21546 ( .A(n20583), .B(n20582), .Z(n20584) );
  XOR U21547 ( .A(n20585), .B(n20584), .Z(n20588) );
  NAND U21548 ( .A(b[0]), .B(a[863]), .Z(n20589) );
  XOR U21549 ( .A(n20588), .B(n20589), .Z(n20591) );
  OR U21550 ( .A(n20567), .B(n20566), .Z(n20571) );
  NANDN U21551 ( .A(n20569), .B(n20568), .Z(n20570) );
  NAND U21552 ( .A(n20571), .B(n20570), .Z(n20590) );
  XNOR U21553 ( .A(n20591), .B(n20590), .Z(n20576) );
  XNOR U21554 ( .A(n20576), .B(n20577), .Z(n20579) );
  XOR U21555 ( .A(n20578), .B(n20579), .Z(n20594) );
  XOR U21556 ( .A(n20594), .B(sreg[1883]), .Z(n20595) );
  XOR U21557 ( .A(n20596), .B(n20595), .Z(c[1883]) );
  NANDN U21558 ( .A(n20577), .B(n20576), .Z(n20581) );
  NAND U21559 ( .A(n20579), .B(n20578), .Z(n20580) );
  NAND U21560 ( .A(n20581), .B(n20580), .Z(n20605) );
  AND U21561 ( .A(b[2]), .B(a[862]), .Z(n20617) );
  AND U21562 ( .A(a[863]), .B(b[1]), .Z(n20615) );
  AND U21563 ( .A(a[861]), .B(b[3]), .Z(n20614) );
  XOR U21564 ( .A(n20615), .B(n20614), .Z(n20616) );
  XOR U21565 ( .A(n20617), .B(n20616), .Z(n20608) );
  NAND U21566 ( .A(b[0]), .B(a[864]), .Z(n20609) );
  XOR U21567 ( .A(n20608), .B(n20609), .Z(n20611) );
  OR U21568 ( .A(n20583), .B(n20582), .Z(n20587) );
  NANDN U21569 ( .A(n20585), .B(n20584), .Z(n20586) );
  NAND U21570 ( .A(n20587), .B(n20586), .Z(n20610) );
  XNOR U21571 ( .A(n20611), .B(n20610), .Z(n20602) );
  NANDN U21572 ( .A(n20589), .B(n20588), .Z(n20593) );
  OR U21573 ( .A(n20591), .B(n20590), .Z(n20592) );
  NAND U21574 ( .A(n20593), .B(n20592), .Z(n20603) );
  XNOR U21575 ( .A(n20602), .B(n20603), .Z(n20604) );
  XOR U21576 ( .A(n20605), .B(n20604), .Z(n20601) );
  NANDN U21577 ( .A(n20594), .B(sreg[1883]), .Z(n20598) );
  OR U21578 ( .A(n20596), .B(n20595), .Z(n20597) );
  NAND U21579 ( .A(n20598), .B(n20597), .Z(n20600) );
  XNOR U21580 ( .A(sreg[1884]), .B(n20600), .Z(n20599) );
  XOR U21581 ( .A(n20601), .B(n20599), .Z(c[1884]) );
  NANDN U21582 ( .A(n20603), .B(n20602), .Z(n20607) );
  NAND U21583 ( .A(n20605), .B(n20604), .Z(n20606) );
  AND U21584 ( .A(n20607), .B(n20606), .Z(n20623) );
  NANDN U21585 ( .A(n20609), .B(n20608), .Z(n20613) );
  OR U21586 ( .A(n20611), .B(n20610), .Z(n20612) );
  AND U21587 ( .A(n20613), .B(n20612), .Z(n20622) );
  AND U21588 ( .A(b[2]), .B(a[863]), .Z(n20627) );
  AND U21589 ( .A(a[864]), .B(b[1]), .Z(n20625) );
  AND U21590 ( .A(a[862]), .B(b[3]), .Z(n20624) );
  XOR U21591 ( .A(n20625), .B(n20624), .Z(n20626) );
  XOR U21592 ( .A(n20627), .B(n20626), .Z(n20630) );
  NAND U21593 ( .A(b[0]), .B(a[865]), .Z(n20631) );
  XOR U21594 ( .A(n20630), .B(n20631), .Z(n20633) );
  OR U21595 ( .A(n20615), .B(n20614), .Z(n20619) );
  NANDN U21596 ( .A(n20617), .B(n20616), .Z(n20618) );
  NAND U21597 ( .A(n20619), .B(n20618), .Z(n20632) );
  XOR U21598 ( .A(n20633), .B(n20632), .Z(n20621) );
  XNOR U21599 ( .A(n20622), .B(n20621), .Z(n20620) );
  XOR U21600 ( .A(n20623), .B(n20620), .Z(n20636) );
  XNOR U21601 ( .A(sreg[1885]), .B(n20636), .Z(n20637) );
  XOR U21602 ( .A(n20638), .B(n20637), .Z(c[1885]) );
  AND U21603 ( .A(b[2]), .B(a[864]), .Z(n20651) );
  AND U21604 ( .A(a[865]), .B(b[1]), .Z(n20649) );
  AND U21605 ( .A(a[863]), .B(b[3]), .Z(n20648) );
  XOR U21606 ( .A(n20649), .B(n20648), .Z(n20650) );
  XOR U21607 ( .A(n20651), .B(n20650), .Z(n20654) );
  NAND U21608 ( .A(b[0]), .B(a[866]), .Z(n20655) );
  XOR U21609 ( .A(n20654), .B(n20655), .Z(n20657) );
  OR U21610 ( .A(n20625), .B(n20624), .Z(n20629) );
  NANDN U21611 ( .A(n20627), .B(n20626), .Z(n20628) );
  NAND U21612 ( .A(n20629), .B(n20628), .Z(n20656) );
  XNOR U21613 ( .A(n20657), .B(n20656), .Z(n20642) );
  NANDN U21614 ( .A(n20631), .B(n20630), .Z(n20635) );
  OR U21615 ( .A(n20633), .B(n20632), .Z(n20634) );
  NAND U21616 ( .A(n20635), .B(n20634), .Z(n20643) );
  XNOR U21617 ( .A(n20642), .B(n20643), .Z(n20644) );
  XOR U21618 ( .A(n20645), .B(n20644), .Z(n20661) );
  NAND U21619 ( .A(sreg[1885]), .B(n20636), .Z(n20640) );
  OR U21620 ( .A(n20638), .B(n20637), .Z(n20639) );
  NAND U21621 ( .A(n20640), .B(n20639), .Z(n20660) );
  XNOR U21622 ( .A(sreg[1886]), .B(n20660), .Z(n20641) );
  XNOR U21623 ( .A(n20661), .B(n20641), .Z(c[1886]) );
  NANDN U21624 ( .A(n20643), .B(n20642), .Z(n20647) );
  NANDN U21625 ( .A(n20645), .B(n20644), .Z(n20646) );
  NAND U21626 ( .A(n20647), .B(n20646), .Z(n20666) );
  AND U21627 ( .A(b[2]), .B(a[865]), .Z(n20672) );
  AND U21628 ( .A(a[866]), .B(b[1]), .Z(n20670) );
  AND U21629 ( .A(a[864]), .B(b[3]), .Z(n20669) );
  XOR U21630 ( .A(n20670), .B(n20669), .Z(n20671) );
  XOR U21631 ( .A(n20672), .B(n20671), .Z(n20675) );
  NAND U21632 ( .A(b[0]), .B(a[867]), .Z(n20676) );
  XOR U21633 ( .A(n20675), .B(n20676), .Z(n20678) );
  OR U21634 ( .A(n20649), .B(n20648), .Z(n20653) );
  NANDN U21635 ( .A(n20651), .B(n20650), .Z(n20652) );
  NAND U21636 ( .A(n20653), .B(n20652), .Z(n20677) );
  XNOR U21637 ( .A(n20678), .B(n20677), .Z(n20663) );
  NANDN U21638 ( .A(n20655), .B(n20654), .Z(n20659) );
  OR U21639 ( .A(n20657), .B(n20656), .Z(n20658) );
  NAND U21640 ( .A(n20659), .B(n20658), .Z(n20664) );
  XNOR U21641 ( .A(n20663), .B(n20664), .Z(n20665) );
  XOR U21642 ( .A(n20666), .B(n20665), .Z(n20683) );
  XNOR U21643 ( .A(sreg[1887]), .B(n20682), .Z(n20662) );
  XOR U21644 ( .A(n20683), .B(n20662), .Z(c[1887]) );
  NANDN U21645 ( .A(n20664), .B(n20663), .Z(n20668) );
  NAND U21646 ( .A(n20666), .B(n20665), .Z(n20667) );
  NAND U21647 ( .A(n20668), .B(n20667), .Z(n20689) );
  AND U21648 ( .A(b[2]), .B(a[866]), .Z(n20697) );
  AND U21649 ( .A(a[867]), .B(b[1]), .Z(n20695) );
  AND U21650 ( .A(a[865]), .B(b[3]), .Z(n20694) );
  XOR U21651 ( .A(n20695), .B(n20694), .Z(n20696) );
  XOR U21652 ( .A(n20697), .B(n20696), .Z(n20690) );
  NAND U21653 ( .A(b[0]), .B(a[868]), .Z(n20691) );
  XOR U21654 ( .A(n20690), .B(n20691), .Z(n20692) );
  OR U21655 ( .A(n20670), .B(n20669), .Z(n20674) );
  NANDN U21656 ( .A(n20672), .B(n20671), .Z(n20673) );
  AND U21657 ( .A(n20674), .B(n20673), .Z(n20693) );
  XOR U21658 ( .A(n20692), .B(n20693), .Z(n20687) );
  NANDN U21659 ( .A(n20676), .B(n20675), .Z(n20680) );
  OR U21660 ( .A(n20678), .B(n20677), .Z(n20679) );
  AND U21661 ( .A(n20680), .B(n20679), .Z(n20688) );
  XOR U21662 ( .A(n20687), .B(n20688), .Z(n20681) );
  XOR U21663 ( .A(n20689), .B(n20681), .Z(n20686) );
  XOR U21664 ( .A(n20685), .B(sreg[1888]), .Z(n20684) );
  XNOR U21665 ( .A(n20686), .B(n20684), .Z(c[1888]) );
  AND U21666 ( .A(b[2]), .B(a[867]), .Z(n20703) );
  AND U21667 ( .A(a[868]), .B(b[1]), .Z(n20701) );
  AND U21668 ( .A(a[866]), .B(b[3]), .Z(n20700) );
  XOR U21669 ( .A(n20701), .B(n20700), .Z(n20702) );
  XOR U21670 ( .A(n20703), .B(n20702), .Z(n20706) );
  NAND U21671 ( .A(b[0]), .B(a[869]), .Z(n20707) );
  XNOR U21672 ( .A(n20706), .B(n20707), .Z(n20708) );
  OR U21673 ( .A(n20695), .B(n20694), .Z(n20699) );
  NANDN U21674 ( .A(n20697), .B(n20696), .Z(n20698) );
  AND U21675 ( .A(n20699), .B(n20698), .Z(n20709) );
  XNOR U21676 ( .A(n20708), .B(n20709), .Z(n20713) );
  XNOR U21677 ( .A(n20712), .B(n20713), .Z(n20714) );
  XNOR U21678 ( .A(n20715), .B(n20714), .Z(n20718) );
  XNOR U21679 ( .A(sreg[1889]), .B(n20718), .Z(n20720) );
  XNOR U21680 ( .A(n20719), .B(n20720), .Z(c[1889]) );
  AND U21681 ( .A(b[2]), .B(a[868]), .Z(n20735) );
  AND U21682 ( .A(a[869]), .B(b[1]), .Z(n20733) );
  AND U21683 ( .A(a[867]), .B(b[3]), .Z(n20732) );
  XOR U21684 ( .A(n20733), .B(n20732), .Z(n20734) );
  XOR U21685 ( .A(n20735), .B(n20734), .Z(n20738) );
  NAND U21686 ( .A(b[0]), .B(a[870]), .Z(n20739) );
  XOR U21687 ( .A(n20738), .B(n20739), .Z(n20741) );
  OR U21688 ( .A(n20701), .B(n20700), .Z(n20705) );
  NANDN U21689 ( .A(n20703), .B(n20702), .Z(n20704) );
  NAND U21690 ( .A(n20705), .B(n20704), .Z(n20740) );
  XNOR U21691 ( .A(n20741), .B(n20740), .Z(n20726) );
  NANDN U21692 ( .A(n20707), .B(n20706), .Z(n20711) );
  NAND U21693 ( .A(n20709), .B(n20708), .Z(n20710) );
  NAND U21694 ( .A(n20711), .B(n20710), .Z(n20727) );
  XNOR U21695 ( .A(n20726), .B(n20727), .Z(n20728) );
  NANDN U21696 ( .A(n20713), .B(n20712), .Z(n20717) );
  NANDN U21697 ( .A(n20715), .B(n20714), .Z(n20716) );
  NAND U21698 ( .A(n20717), .B(n20716), .Z(n20729) );
  XOR U21699 ( .A(n20728), .B(n20729), .Z(n20725) );
  NAND U21700 ( .A(sreg[1889]), .B(n20718), .Z(n20722) );
  NANDN U21701 ( .A(n20720), .B(n20719), .Z(n20721) );
  NAND U21702 ( .A(n20722), .B(n20721), .Z(n20724) );
  XNOR U21703 ( .A(sreg[1890]), .B(n20724), .Z(n20723) );
  XNOR U21704 ( .A(n20725), .B(n20723), .Z(c[1890]) );
  NANDN U21705 ( .A(n20727), .B(n20726), .Z(n20731) );
  NANDN U21706 ( .A(n20729), .B(n20728), .Z(n20730) );
  NAND U21707 ( .A(n20731), .B(n20730), .Z(n20759) );
  AND U21708 ( .A(b[2]), .B(a[869]), .Z(n20753) );
  AND U21709 ( .A(a[870]), .B(b[1]), .Z(n20751) );
  AND U21710 ( .A(a[868]), .B(b[3]), .Z(n20750) );
  XOR U21711 ( .A(n20751), .B(n20750), .Z(n20752) );
  XOR U21712 ( .A(n20753), .B(n20752), .Z(n20744) );
  NAND U21713 ( .A(b[0]), .B(a[871]), .Z(n20745) );
  XOR U21714 ( .A(n20744), .B(n20745), .Z(n20747) );
  OR U21715 ( .A(n20733), .B(n20732), .Z(n20737) );
  NANDN U21716 ( .A(n20735), .B(n20734), .Z(n20736) );
  NAND U21717 ( .A(n20737), .B(n20736), .Z(n20746) );
  XNOR U21718 ( .A(n20747), .B(n20746), .Z(n20756) );
  NANDN U21719 ( .A(n20739), .B(n20738), .Z(n20743) );
  OR U21720 ( .A(n20741), .B(n20740), .Z(n20742) );
  NAND U21721 ( .A(n20743), .B(n20742), .Z(n20757) );
  XNOR U21722 ( .A(n20756), .B(n20757), .Z(n20758) );
  XNOR U21723 ( .A(n20759), .B(n20758), .Z(n20762) );
  XOR U21724 ( .A(sreg[1891]), .B(n20762), .Z(n20764) );
  XNOR U21725 ( .A(n20763), .B(n20764), .Z(c[1891]) );
  NANDN U21726 ( .A(n20745), .B(n20744), .Z(n20749) );
  OR U21727 ( .A(n20747), .B(n20746), .Z(n20748) );
  NAND U21728 ( .A(n20749), .B(n20748), .Z(n20782) );
  AND U21729 ( .A(b[2]), .B(a[870]), .Z(n20773) );
  AND U21730 ( .A(a[871]), .B(b[1]), .Z(n20771) );
  AND U21731 ( .A(a[869]), .B(b[3]), .Z(n20770) );
  XOR U21732 ( .A(n20771), .B(n20770), .Z(n20772) );
  XOR U21733 ( .A(n20773), .B(n20772), .Z(n20776) );
  NAND U21734 ( .A(b[0]), .B(a[872]), .Z(n20777) );
  XNOR U21735 ( .A(n20776), .B(n20777), .Z(n20778) );
  OR U21736 ( .A(n20751), .B(n20750), .Z(n20755) );
  NANDN U21737 ( .A(n20753), .B(n20752), .Z(n20754) );
  AND U21738 ( .A(n20755), .B(n20754), .Z(n20779) );
  XNOR U21739 ( .A(n20778), .B(n20779), .Z(n20783) );
  XNOR U21740 ( .A(n20782), .B(n20783), .Z(n20784) );
  NANDN U21741 ( .A(n20757), .B(n20756), .Z(n20761) );
  NAND U21742 ( .A(n20759), .B(n20758), .Z(n20760) );
  NAND U21743 ( .A(n20761), .B(n20760), .Z(n20785) );
  XOR U21744 ( .A(n20784), .B(n20785), .Z(n20769) );
  OR U21745 ( .A(n20762), .B(sreg[1891]), .Z(n20766) );
  NAND U21746 ( .A(n20764), .B(n20763), .Z(n20765) );
  AND U21747 ( .A(n20766), .B(n20765), .Z(n20768) );
  XOR U21748 ( .A(sreg[1892]), .B(n20768), .Z(n20767) );
  XNOR U21749 ( .A(n20769), .B(n20767), .Z(c[1892]) );
  AND U21750 ( .A(b[2]), .B(a[871]), .Z(n20802) );
  AND U21751 ( .A(a[872]), .B(b[1]), .Z(n20800) );
  AND U21752 ( .A(a[870]), .B(b[3]), .Z(n20799) );
  XOR U21753 ( .A(n20800), .B(n20799), .Z(n20801) );
  XOR U21754 ( .A(n20802), .B(n20801), .Z(n20805) );
  NAND U21755 ( .A(b[0]), .B(a[873]), .Z(n20806) );
  XOR U21756 ( .A(n20805), .B(n20806), .Z(n20808) );
  OR U21757 ( .A(n20771), .B(n20770), .Z(n20775) );
  NANDN U21758 ( .A(n20773), .B(n20772), .Z(n20774) );
  NAND U21759 ( .A(n20775), .B(n20774), .Z(n20807) );
  XNOR U21760 ( .A(n20808), .B(n20807), .Z(n20793) );
  NANDN U21761 ( .A(n20777), .B(n20776), .Z(n20781) );
  NAND U21762 ( .A(n20779), .B(n20778), .Z(n20780) );
  NAND U21763 ( .A(n20781), .B(n20780), .Z(n20794) );
  XNOR U21764 ( .A(n20793), .B(n20794), .Z(n20795) );
  NANDN U21765 ( .A(n20783), .B(n20782), .Z(n20787) );
  NANDN U21766 ( .A(n20785), .B(n20784), .Z(n20786) );
  AND U21767 ( .A(n20787), .B(n20786), .Z(n20796) );
  XNOR U21768 ( .A(n20795), .B(n20796), .Z(n20788) );
  XOR U21769 ( .A(sreg[1893]), .B(n20788), .Z(n20789) );
  XOR U21770 ( .A(n20790), .B(n20789), .Z(c[1893]) );
  OR U21771 ( .A(n20788), .B(sreg[1893]), .Z(n20792) );
  NANDN U21772 ( .A(n20790), .B(n20789), .Z(n20791) );
  AND U21773 ( .A(n20792), .B(n20791), .Z(n20830) );
  NANDN U21774 ( .A(n20794), .B(n20793), .Z(n20798) );
  NAND U21775 ( .A(n20796), .B(n20795), .Z(n20797) );
  NAND U21776 ( .A(n20798), .B(n20797), .Z(n20815) );
  AND U21777 ( .A(b[2]), .B(a[872]), .Z(n20821) );
  AND U21778 ( .A(a[873]), .B(b[1]), .Z(n20819) );
  AND U21779 ( .A(a[871]), .B(b[3]), .Z(n20818) );
  XOR U21780 ( .A(n20819), .B(n20818), .Z(n20820) );
  XOR U21781 ( .A(n20821), .B(n20820), .Z(n20824) );
  NAND U21782 ( .A(b[0]), .B(a[874]), .Z(n20825) );
  XOR U21783 ( .A(n20824), .B(n20825), .Z(n20827) );
  OR U21784 ( .A(n20800), .B(n20799), .Z(n20804) );
  NANDN U21785 ( .A(n20802), .B(n20801), .Z(n20803) );
  NAND U21786 ( .A(n20804), .B(n20803), .Z(n20826) );
  XNOR U21787 ( .A(n20827), .B(n20826), .Z(n20812) );
  NANDN U21788 ( .A(n20806), .B(n20805), .Z(n20810) );
  OR U21789 ( .A(n20808), .B(n20807), .Z(n20809) );
  NAND U21790 ( .A(n20810), .B(n20809), .Z(n20813) );
  XNOR U21791 ( .A(n20812), .B(n20813), .Z(n20814) );
  XNOR U21792 ( .A(n20815), .B(n20814), .Z(n20831) );
  XOR U21793 ( .A(sreg[1894]), .B(n20831), .Z(n20811) );
  XOR U21794 ( .A(n20830), .B(n20811), .Z(c[1894]) );
  NANDN U21795 ( .A(n20813), .B(n20812), .Z(n20817) );
  NAND U21796 ( .A(n20815), .B(n20814), .Z(n20816) );
  NAND U21797 ( .A(n20817), .B(n20816), .Z(n20838) );
  AND U21798 ( .A(b[2]), .B(a[873]), .Z(n20844) );
  AND U21799 ( .A(a[874]), .B(b[1]), .Z(n20842) );
  AND U21800 ( .A(a[872]), .B(b[3]), .Z(n20841) );
  XOR U21801 ( .A(n20842), .B(n20841), .Z(n20843) );
  XOR U21802 ( .A(n20844), .B(n20843), .Z(n20847) );
  NAND U21803 ( .A(b[0]), .B(a[875]), .Z(n20848) );
  XOR U21804 ( .A(n20847), .B(n20848), .Z(n20850) );
  OR U21805 ( .A(n20819), .B(n20818), .Z(n20823) );
  NANDN U21806 ( .A(n20821), .B(n20820), .Z(n20822) );
  NAND U21807 ( .A(n20823), .B(n20822), .Z(n20849) );
  XNOR U21808 ( .A(n20850), .B(n20849), .Z(n20835) );
  NANDN U21809 ( .A(n20825), .B(n20824), .Z(n20829) );
  OR U21810 ( .A(n20827), .B(n20826), .Z(n20828) );
  NAND U21811 ( .A(n20829), .B(n20828), .Z(n20836) );
  XNOR U21812 ( .A(n20835), .B(n20836), .Z(n20837) );
  XNOR U21813 ( .A(n20838), .B(n20837), .Z(n20834) );
  XOR U21814 ( .A(n20833), .B(sreg[1895]), .Z(n20832) );
  XOR U21815 ( .A(n20834), .B(n20832), .Z(c[1895]) );
  NANDN U21816 ( .A(n20836), .B(n20835), .Z(n20840) );
  NAND U21817 ( .A(n20838), .B(n20837), .Z(n20839) );
  NAND U21818 ( .A(n20840), .B(n20839), .Z(n20856) );
  AND U21819 ( .A(b[2]), .B(a[874]), .Z(n20862) );
  AND U21820 ( .A(a[875]), .B(b[1]), .Z(n20860) );
  AND U21821 ( .A(a[873]), .B(b[3]), .Z(n20859) );
  XOR U21822 ( .A(n20860), .B(n20859), .Z(n20861) );
  XOR U21823 ( .A(n20862), .B(n20861), .Z(n20865) );
  NAND U21824 ( .A(b[0]), .B(a[876]), .Z(n20866) );
  XOR U21825 ( .A(n20865), .B(n20866), .Z(n20868) );
  OR U21826 ( .A(n20842), .B(n20841), .Z(n20846) );
  NANDN U21827 ( .A(n20844), .B(n20843), .Z(n20845) );
  NAND U21828 ( .A(n20846), .B(n20845), .Z(n20867) );
  XNOR U21829 ( .A(n20868), .B(n20867), .Z(n20853) );
  NANDN U21830 ( .A(n20848), .B(n20847), .Z(n20852) );
  OR U21831 ( .A(n20850), .B(n20849), .Z(n20851) );
  NAND U21832 ( .A(n20852), .B(n20851), .Z(n20854) );
  XNOR U21833 ( .A(n20853), .B(n20854), .Z(n20855) );
  XNOR U21834 ( .A(n20856), .B(n20855), .Z(n20871) );
  XNOR U21835 ( .A(n20871), .B(sreg[1896]), .Z(n20873) );
  XNOR U21836 ( .A(n20872), .B(n20873), .Z(c[1896]) );
  NANDN U21837 ( .A(n20854), .B(n20853), .Z(n20858) );
  NAND U21838 ( .A(n20856), .B(n20855), .Z(n20857) );
  NAND U21839 ( .A(n20858), .B(n20857), .Z(n20880) );
  AND U21840 ( .A(b[2]), .B(a[875]), .Z(n20886) );
  AND U21841 ( .A(a[876]), .B(b[1]), .Z(n20884) );
  AND U21842 ( .A(a[874]), .B(b[3]), .Z(n20883) );
  XOR U21843 ( .A(n20884), .B(n20883), .Z(n20885) );
  XOR U21844 ( .A(n20886), .B(n20885), .Z(n20889) );
  NAND U21845 ( .A(b[0]), .B(a[877]), .Z(n20890) );
  XOR U21846 ( .A(n20889), .B(n20890), .Z(n20892) );
  OR U21847 ( .A(n20860), .B(n20859), .Z(n20864) );
  NANDN U21848 ( .A(n20862), .B(n20861), .Z(n20863) );
  NAND U21849 ( .A(n20864), .B(n20863), .Z(n20891) );
  XNOR U21850 ( .A(n20892), .B(n20891), .Z(n20877) );
  NANDN U21851 ( .A(n20866), .B(n20865), .Z(n20870) );
  OR U21852 ( .A(n20868), .B(n20867), .Z(n20869) );
  NAND U21853 ( .A(n20870), .B(n20869), .Z(n20878) );
  XNOR U21854 ( .A(n20877), .B(n20878), .Z(n20879) );
  XOR U21855 ( .A(n20880), .B(n20879), .Z(n20896) );
  NAND U21856 ( .A(n20871), .B(sreg[1896]), .Z(n20875) );
  NANDN U21857 ( .A(n20873), .B(n20872), .Z(n20874) );
  NAND U21858 ( .A(n20875), .B(n20874), .Z(n20895) );
  XNOR U21859 ( .A(sreg[1897]), .B(n20895), .Z(n20876) );
  XOR U21860 ( .A(n20896), .B(n20876), .Z(c[1897]) );
  NANDN U21861 ( .A(n20878), .B(n20877), .Z(n20882) );
  NAND U21862 ( .A(n20880), .B(n20879), .Z(n20881) );
  NAND U21863 ( .A(n20882), .B(n20881), .Z(n20903) );
  AND U21864 ( .A(b[2]), .B(a[876]), .Z(n20909) );
  AND U21865 ( .A(a[877]), .B(b[1]), .Z(n20907) );
  AND U21866 ( .A(a[875]), .B(b[3]), .Z(n20906) );
  XOR U21867 ( .A(n20907), .B(n20906), .Z(n20908) );
  XOR U21868 ( .A(n20909), .B(n20908), .Z(n20912) );
  NAND U21869 ( .A(b[0]), .B(a[878]), .Z(n20913) );
  XOR U21870 ( .A(n20912), .B(n20913), .Z(n20915) );
  OR U21871 ( .A(n20884), .B(n20883), .Z(n20888) );
  NANDN U21872 ( .A(n20886), .B(n20885), .Z(n20887) );
  NAND U21873 ( .A(n20888), .B(n20887), .Z(n20914) );
  XNOR U21874 ( .A(n20915), .B(n20914), .Z(n20900) );
  NANDN U21875 ( .A(n20890), .B(n20889), .Z(n20894) );
  OR U21876 ( .A(n20892), .B(n20891), .Z(n20893) );
  NAND U21877 ( .A(n20894), .B(n20893), .Z(n20901) );
  XNOR U21878 ( .A(n20900), .B(n20901), .Z(n20902) );
  XOR U21879 ( .A(n20903), .B(n20902), .Z(n20899) );
  XNOR U21880 ( .A(sreg[1898]), .B(n20898), .Z(n20897) );
  XOR U21881 ( .A(n20899), .B(n20897), .Z(c[1898]) );
  NANDN U21882 ( .A(n20901), .B(n20900), .Z(n20905) );
  NAND U21883 ( .A(n20903), .B(n20902), .Z(n20904) );
  NAND U21884 ( .A(n20905), .B(n20904), .Z(n20921) );
  AND U21885 ( .A(b[2]), .B(a[877]), .Z(n20927) );
  AND U21886 ( .A(a[878]), .B(b[1]), .Z(n20925) );
  AND U21887 ( .A(a[876]), .B(b[3]), .Z(n20924) );
  XOR U21888 ( .A(n20925), .B(n20924), .Z(n20926) );
  XOR U21889 ( .A(n20927), .B(n20926), .Z(n20930) );
  NAND U21890 ( .A(b[0]), .B(a[879]), .Z(n20931) );
  XOR U21891 ( .A(n20930), .B(n20931), .Z(n20933) );
  OR U21892 ( .A(n20907), .B(n20906), .Z(n20911) );
  NANDN U21893 ( .A(n20909), .B(n20908), .Z(n20910) );
  NAND U21894 ( .A(n20911), .B(n20910), .Z(n20932) );
  XNOR U21895 ( .A(n20933), .B(n20932), .Z(n20918) );
  NANDN U21896 ( .A(n20913), .B(n20912), .Z(n20917) );
  OR U21897 ( .A(n20915), .B(n20914), .Z(n20916) );
  NAND U21898 ( .A(n20917), .B(n20916), .Z(n20919) );
  XNOR U21899 ( .A(n20918), .B(n20919), .Z(n20920) );
  XNOR U21900 ( .A(n20921), .B(n20920), .Z(n20936) );
  XNOR U21901 ( .A(n20936), .B(sreg[1899]), .Z(n20937) );
  XOR U21902 ( .A(n20938), .B(n20937), .Z(c[1899]) );
  NANDN U21903 ( .A(n20919), .B(n20918), .Z(n20923) );
  NAND U21904 ( .A(n20921), .B(n20920), .Z(n20922) );
  NAND U21905 ( .A(n20923), .B(n20922), .Z(n20947) );
  AND U21906 ( .A(b[2]), .B(a[878]), .Z(n20953) );
  AND U21907 ( .A(a[879]), .B(b[1]), .Z(n20951) );
  AND U21908 ( .A(a[877]), .B(b[3]), .Z(n20950) );
  XOR U21909 ( .A(n20951), .B(n20950), .Z(n20952) );
  XOR U21910 ( .A(n20953), .B(n20952), .Z(n20956) );
  NAND U21911 ( .A(b[0]), .B(a[880]), .Z(n20957) );
  XOR U21912 ( .A(n20956), .B(n20957), .Z(n20959) );
  OR U21913 ( .A(n20925), .B(n20924), .Z(n20929) );
  NANDN U21914 ( .A(n20927), .B(n20926), .Z(n20928) );
  NAND U21915 ( .A(n20929), .B(n20928), .Z(n20958) );
  XNOR U21916 ( .A(n20959), .B(n20958), .Z(n20944) );
  NANDN U21917 ( .A(n20931), .B(n20930), .Z(n20935) );
  OR U21918 ( .A(n20933), .B(n20932), .Z(n20934) );
  NAND U21919 ( .A(n20935), .B(n20934), .Z(n20945) );
  XNOR U21920 ( .A(n20944), .B(n20945), .Z(n20946) );
  XOR U21921 ( .A(n20947), .B(n20946), .Z(n20943) );
  NAND U21922 ( .A(n20936), .B(sreg[1899]), .Z(n20940) );
  OR U21923 ( .A(n20938), .B(n20937), .Z(n20939) );
  NAND U21924 ( .A(n20940), .B(n20939), .Z(n20942) );
  XNOR U21925 ( .A(sreg[1900]), .B(n20942), .Z(n20941) );
  XOR U21926 ( .A(n20943), .B(n20941), .Z(c[1900]) );
  NANDN U21927 ( .A(n20945), .B(n20944), .Z(n20949) );
  NAND U21928 ( .A(n20947), .B(n20946), .Z(n20948) );
  NAND U21929 ( .A(n20949), .B(n20948), .Z(n20965) );
  AND U21930 ( .A(b[2]), .B(a[879]), .Z(n20971) );
  AND U21931 ( .A(a[880]), .B(b[1]), .Z(n20969) );
  AND U21932 ( .A(a[878]), .B(b[3]), .Z(n20968) );
  XOR U21933 ( .A(n20969), .B(n20968), .Z(n20970) );
  XOR U21934 ( .A(n20971), .B(n20970), .Z(n20974) );
  NAND U21935 ( .A(b[0]), .B(a[881]), .Z(n20975) );
  XOR U21936 ( .A(n20974), .B(n20975), .Z(n20977) );
  OR U21937 ( .A(n20951), .B(n20950), .Z(n20955) );
  NANDN U21938 ( .A(n20953), .B(n20952), .Z(n20954) );
  NAND U21939 ( .A(n20955), .B(n20954), .Z(n20976) );
  XNOR U21940 ( .A(n20977), .B(n20976), .Z(n20962) );
  NANDN U21941 ( .A(n20957), .B(n20956), .Z(n20961) );
  OR U21942 ( .A(n20959), .B(n20958), .Z(n20960) );
  NAND U21943 ( .A(n20961), .B(n20960), .Z(n20963) );
  XNOR U21944 ( .A(n20962), .B(n20963), .Z(n20964) );
  XNOR U21945 ( .A(n20965), .B(n20964), .Z(n20980) );
  XNOR U21946 ( .A(n20980), .B(sreg[1901]), .Z(n20981) );
  XOR U21947 ( .A(n20982), .B(n20981), .Z(c[1901]) );
  NANDN U21948 ( .A(n20963), .B(n20962), .Z(n20967) );
  NAND U21949 ( .A(n20965), .B(n20964), .Z(n20966) );
  NAND U21950 ( .A(n20967), .B(n20966), .Z(n20991) );
  AND U21951 ( .A(b[2]), .B(a[880]), .Z(n20997) );
  AND U21952 ( .A(a[881]), .B(b[1]), .Z(n20995) );
  AND U21953 ( .A(a[879]), .B(b[3]), .Z(n20994) );
  XOR U21954 ( .A(n20995), .B(n20994), .Z(n20996) );
  XOR U21955 ( .A(n20997), .B(n20996), .Z(n21000) );
  NAND U21956 ( .A(b[0]), .B(a[882]), .Z(n21001) );
  XOR U21957 ( .A(n21000), .B(n21001), .Z(n21003) );
  OR U21958 ( .A(n20969), .B(n20968), .Z(n20973) );
  NANDN U21959 ( .A(n20971), .B(n20970), .Z(n20972) );
  NAND U21960 ( .A(n20973), .B(n20972), .Z(n21002) );
  XNOR U21961 ( .A(n21003), .B(n21002), .Z(n20988) );
  NANDN U21962 ( .A(n20975), .B(n20974), .Z(n20979) );
  OR U21963 ( .A(n20977), .B(n20976), .Z(n20978) );
  NAND U21964 ( .A(n20979), .B(n20978), .Z(n20989) );
  XNOR U21965 ( .A(n20988), .B(n20989), .Z(n20990) );
  XOR U21966 ( .A(n20991), .B(n20990), .Z(n20987) );
  NAND U21967 ( .A(n20980), .B(sreg[1901]), .Z(n20984) );
  OR U21968 ( .A(n20982), .B(n20981), .Z(n20983) );
  NAND U21969 ( .A(n20984), .B(n20983), .Z(n20986) );
  XNOR U21970 ( .A(sreg[1902]), .B(n20986), .Z(n20985) );
  XOR U21971 ( .A(n20987), .B(n20985), .Z(c[1902]) );
  NANDN U21972 ( .A(n20989), .B(n20988), .Z(n20993) );
  NAND U21973 ( .A(n20991), .B(n20990), .Z(n20992) );
  NAND U21974 ( .A(n20993), .B(n20992), .Z(n21009) );
  AND U21975 ( .A(b[2]), .B(a[881]), .Z(n21015) );
  AND U21976 ( .A(a[882]), .B(b[1]), .Z(n21013) );
  AND U21977 ( .A(a[880]), .B(b[3]), .Z(n21012) );
  XOR U21978 ( .A(n21013), .B(n21012), .Z(n21014) );
  XOR U21979 ( .A(n21015), .B(n21014), .Z(n21018) );
  NAND U21980 ( .A(b[0]), .B(a[883]), .Z(n21019) );
  XOR U21981 ( .A(n21018), .B(n21019), .Z(n21021) );
  OR U21982 ( .A(n20995), .B(n20994), .Z(n20999) );
  NANDN U21983 ( .A(n20997), .B(n20996), .Z(n20998) );
  NAND U21984 ( .A(n20999), .B(n20998), .Z(n21020) );
  XNOR U21985 ( .A(n21021), .B(n21020), .Z(n21006) );
  NANDN U21986 ( .A(n21001), .B(n21000), .Z(n21005) );
  OR U21987 ( .A(n21003), .B(n21002), .Z(n21004) );
  NAND U21988 ( .A(n21005), .B(n21004), .Z(n21007) );
  XNOR U21989 ( .A(n21006), .B(n21007), .Z(n21008) );
  XNOR U21990 ( .A(n21009), .B(n21008), .Z(n21024) );
  XNOR U21991 ( .A(n21024), .B(sreg[1903]), .Z(n21025) );
  XOR U21992 ( .A(n21026), .B(n21025), .Z(c[1903]) );
  NANDN U21993 ( .A(n21007), .B(n21006), .Z(n21011) );
  NAND U21994 ( .A(n21009), .B(n21008), .Z(n21010) );
  NAND U21995 ( .A(n21011), .B(n21010), .Z(n21037) );
  AND U21996 ( .A(b[2]), .B(a[882]), .Z(n21043) );
  AND U21997 ( .A(a[883]), .B(b[1]), .Z(n21041) );
  AND U21998 ( .A(a[881]), .B(b[3]), .Z(n21040) );
  XOR U21999 ( .A(n21041), .B(n21040), .Z(n21042) );
  XOR U22000 ( .A(n21043), .B(n21042), .Z(n21046) );
  NAND U22001 ( .A(b[0]), .B(a[884]), .Z(n21047) );
  XOR U22002 ( .A(n21046), .B(n21047), .Z(n21049) );
  OR U22003 ( .A(n21013), .B(n21012), .Z(n21017) );
  NANDN U22004 ( .A(n21015), .B(n21014), .Z(n21016) );
  NAND U22005 ( .A(n21017), .B(n21016), .Z(n21048) );
  XNOR U22006 ( .A(n21049), .B(n21048), .Z(n21034) );
  NANDN U22007 ( .A(n21019), .B(n21018), .Z(n21023) );
  OR U22008 ( .A(n21021), .B(n21020), .Z(n21022) );
  NAND U22009 ( .A(n21023), .B(n21022), .Z(n21035) );
  XNOR U22010 ( .A(n21034), .B(n21035), .Z(n21036) );
  XNOR U22011 ( .A(n21037), .B(n21036), .Z(n21029) );
  XOR U22012 ( .A(sreg[1904]), .B(n21029), .Z(n21030) );
  NAND U22013 ( .A(n21024), .B(sreg[1903]), .Z(n21028) );
  OR U22014 ( .A(n21026), .B(n21025), .Z(n21027) );
  NAND U22015 ( .A(n21028), .B(n21027), .Z(n21031) );
  XOR U22016 ( .A(n21030), .B(n21031), .Z(c[1904]) );
  OR U22017 ( .A(n21029), .B(sreg[1904]), .Z(n21033) );
  NANDN U22018 ( .A(n21031), .B(n21030), .Z(n21032) );
  AND U22019 ( .A(n21033), .B(n21032), .Z(n21071) );
  NANDN U22020 ( .A(n21035), .B(n21034), .Z(n21039) );
  NAND U22021 ( .A(n21037), .B(n21036), .Z(n21038) );
  NAND U22022 ( .A(n21039), .B(n21038), .Z(n21056) );
  AND U22023 ( .A(b[2]), .B(a[883]), .Z(n21062) );
  AND U22024 ( .A(a[884]), .B(b[1]), .Z(n21060) );
  AND U22025 ( .A(a[882]), .B(b[3]), .Z(n21059) );
  XOR U22026 ( .A(n21060), .B(n21059), .Z(n21061) );
  XOR U22027 ( .A(n21062), .B(n21061), .Z(n21065) );
  NAND U22028 ( .A(b[0]), .B(a[885]), .Z(n21066) );
  XOR U22029 ( .A(n21065), .B(n21066), .Z(n21068) );
  OR U22030 ( .A(n21041), .B(n21040), .Z(n21045) );
  NANDN U22031 ( .A(n21043), .B(n21042), .Z(n21044) );
  NAND U22032 ( .A(n21045), .B(n21044), .Z(n21067) );
  XNOR U22033 ( .A(n21068), .B(n21067), .Z(n21053) );
  NANDN U22034 ( .A(n21047), .B(n21046), .Z(n21051) );
  OR U22035 ( .A(n21049), .B(n21048), .Z(n21050) );
  NAND U22036 ( .A(n21051), .B(n21050), .Z(n21054) );
  XNOR U22037 ( .A(n21053), .B(n21054), .Z(n21055) );
  XNOR U22038 ( .A(n21056), .B(n21055), .Z(n21072) );
  XOR U22039 ( .A(sreg[1905]), .B(n21072), .Z(n21052) );
  XOR U22040 ( .A(n21071), .B(n21052), .Z(c[1905]) );
  NANDN U22041 ( .A(n21054), .B(n21053), .Z(n21058) );
  NAND U22042 ( .A(n21056), .B(n21055), .Z(n21057) );
  NAND U22043 ( .A(n21058), .B(n21057), .Z(n21079) );
  AND U22044 ( .A(b[2]), .B(a[884]), .Z(n21085) );
  AND U22045 ( .A(a[885]), .B(b[1]), .Z(n21083) );
  AND U22046 ( .A(a[883]), .B(b[3]), .Z(n21082) );
  XOR U22047 ( .A(n21083), .B(n21082), .Z(n21084) );
  XOR U22048 ( .A(n21085), .B(n21084), .Z(n21088) );
  NAND U22049 ( .A(b[0]), .B(a[886]), .Z(n21089) );
  XOR U22050 ( .A(n21088), .B(n21089), .Z(n21091) );
  OR U22051 ( .A(n21060), .B(n21059), .Z(n21064) );
  NANDN U22052 ( .A(n21062), .B(n21061), .Z(n21063) );
  NAND U22053 ( .A(n21064), .B(n21063), .Z(n21090) );
  XNOR U22054 ( .A(n21091), .B(n21090), .Z(n21076) );
  NANDN U22055 ( .A(n21066), .B(n21065), .Z(n21070) );
  OR U22056 ( .A(n21068), .B(n21067), .Z(n21069) );
  NAND U22057 ( .A(n21070), .B(n21069), .Z(n21077) );
  XNOR U22058 ( .A(n21076), .B(n21077), .Z(n21078) );
  XNOR U22059 ( .A(n21079), .B(n21078), .Z(n21075) );
  XOR U22060 ( .A(n21074), .B(sreg[1906]), .Z(n21073) );
  XOR U22061 ( .A(n21075), .B(n21073), .Z(c[1906]) );
  NANDN U22062 ( .A(n21077), .B(n21076), .Z(n21081) );
  NAND U22063 ( .A(n21079), .B(n21078), .Z(n21080) );
  NAND U22064 ( .A(n21081), .B(n21080), .Z(n21102) );
  AND U22065 ( .A(b[2]), .B(a[885]), .Z(n21108) );
  AND U22066 ( .A(a[886]), .B(b[1]), .Z(n21106) );
  AND U22067 ( .A(a[884]), .B(b[3]), .Z(n21105) );
  XOR U22068 ( .A(n21106), .B(n21105), .Z(n21107) );
  XOR U22069 ( .A(n21108), .B(n21107), .Z(n21111) );
  NAND U22070 ( .A(b[0]), .B(a[887]), .Z(n21112) );
  XOR U22071 ( .A(n21111), .B(n21112), .Z(n21114) );
  OR U22072 ( .A(n21083), .B(n21082), .Z(n21087) );
  NANDN U22073 ( .A(n21085), .B(n21084), .Z(n21086) );
  NAND U22074 ( .A(n21087), .B(n21086), .Z(n21113) );
  XNOR U22075 ( .A(n21114), .B(n21113), .Z(n21099) );
  NANDN U22076 ( .A(n21089), .B(n21088), .Z(n21093) );
  OR U22077 ( .A(n21091), .B(n21090), .Z(n21092) );
  NAND U22078 ( .A(n21093), .B(n21092), .Z(n21100) );
  XNOR U22079 ( .A(n21099), .B(n21100), .Z(n21101) );
  XNOR U22080 ( .A(n21102), .B(n21101), .Z(n21094) );
  XNOR U22081 ( .A(n21094), .B(sreg[1907]), .Z(n21096) );
  XNOR U22082 ( .A(n21095), .B(n21096), .Z(c[1907]) );
  NAND U22083 ( .A(n21094), .B(sreg[1907]), .Z(n21098) );
  NANDN U22084 ( .A(n21096), .B(n21095), .Z(n21097) );
  AND U22085 ( .A(n21098), .B(n21097), .Z(n21137) );
  NANDN U22086 ( .A(n21100), .B(n21099), .Z(n21104) );
  NAND U22087 ( .A(n21102), .B(n21101), .Z(n21103) );
  NAND U22088 ( .A(n21104), .B(n21103), .Z(n21121) );
  AND U22089 ( .A(b[2]), .B(a[886]), .Z(n21127) );
  AND U22090 ( .A(a[887]), .B(b[1]), .Z(n21125) );
  AND U22091 ( .A(a[885]), .B(b[3]), .Z(n21124) );
  XOR U22092 ( .A(n21125), .B(n21124), .Z(n21126) );
  XOR U22093 ( .A(n21127), .B(n21126), .Z(n21130) );
  NAND U22094 ( .A(b[0]), .B(a[888]), .Z(n21131) );
  XOR U22095 ( .A(n21130), .B(n21131), .Z(n21133) );
  OR U22096 ( .A(n21106), .B(n21105), .Z(n21110) );
  NANDN U22097 ( .A(n21108), .B(n21107), .Z(n21109) );
  NAND U22098 ( .A(n21110), .B(n21109), .Z(n21132) );
  XNOR U22099 ( .A(n21133), .B(n21132), .Z(n21118) );
  NANDN U22100 ( .A(n21112), .B(n21111), .Z(n21116) );
  OR U22101 ( .A(n21114), .B(n21113), .Z(n21115) );
  NAND U22102 ( .A(n21116), .B(n21115), .Z(n21119) );
  XNOR U22103 ( .A(n21118), .B(n21119), .Z(n21120) );
  XNOR U22104 ( .A(n21121), .B(n21120), .Z(n21136) );
  XNOR U22105 ( .A(sreg[1908]), .B(n21136), .Z(n21117) );
  XOR U22106 ( .A(n21137), .B(n21117), .Z(c[1908]) );
  NANDN U22107 ( .A(n21119), .B(n21118), .Z(n21123) );
  NAND U22108 ( .A(n21121), .B(n21120), .Z(n21122) );
  NAND U22109 ( .A(n21123), .B(n21122), .Z(n21144) );
  AND U22110 ( .A(b[2]), .B(a[887]), .Z(n21150) );
  AND U22111 ( .A(a[888]), .B(b[1]), .Z(n21148) );
  AND U22112 ( .A(a[886]), .B(b[3]), .Z(n21147) );
  XOR U22113 ( .A(n21148), .B(n21147), .Z(n21149) );
  XOR U22114 ( .A(n21150), .B(n21149), .Z(n21153) );
  NAND U22115 ( .A(b[0]), .B(a[889]), .Z(n21154) );
  XOR U22116 ( .A(n21153), .B(n21154), .Z(n21156) );
  OR U22117 ( .A(n21125), .B(n21124), .Z(n21129) );
  NANDN U22118 ( .A(n21127), .B(n21126), .Z(n21128) );
  NAND U22119 ( .A(n21129), .B(n21128), .Z(n21155) );
  XNOR U22120 ( .A(n21156), .B(n21155), .Z(n21141) );
  NANDN U22121 ( .A(n21131), .B(n21130), .Z(n21135) );
  OR U22122 ( .A(n21133), .B(n21132), .Z(n21134) );
  NAND U22123 ( .A(n21135), .B(n21134), .Z(n21142) );
  XNOR U22124 ( .A(n21141), .B(n21142), .Z(n21143) );
  XNOR U22125 ( .A(n21144), .B(n21143), .Z(n21140) );
  XOR U22126 ( .A(n21139), .B(sreg[1909]), .Z(n21138) );
  XOR U22127 ( .A(n21140), .B(n21138), .Z(c[1909]) );
  NANDN U22128 ( .A(n21142), .B(n21141), .Z(n21146) );
  NAND U22129 ( .A(n21144), .B(n21143), .Z(n21145) );
  NAND U22130 ( .A(n21146), .B(n21145), .Z(n21162) );
  AND U22131 ( .A(b[2]), .B(a[888]), .Z(n21168) );
  AND U22132 ( .A(a[889]), .B(b[1]), .Z(n21166) );
  AND U22133 ( .A(a[887]), .B(b[3]), .Z(n21165) );
  XOR U22134 ( .A(n21166), .B(n21165), .Z(n21167) );
  XOR U22135 ( .A(n21168), .B(n21167), .Z(n21171) );
  NAND U22136 ( .A(b[0]), .B(a[890]), .Z(n21172) );
  XOR U22137 ( .A(n21171), .B(n21172), .Z(n21174) );
  OR U22138 ( .A(n21148), .B(n21147), .Z(n21152) );
  NANDN U22139 ( .A(n21150), .B(n21149), .Z(n21151) );
  NAND U22140 ( .A(n21152), .B(n21151), .Z(n21173) );
  XNOR U22141 ( .A(n21174), .B(n21173), .Z(n21159) );
  NANDN U22142 ( .A(n21154), .B(n21153), .Z(n21158) );
  OR U22143 ( .A(n21156), .B(n21155), .Z(n21157) );
  NAND U22144 ( .A(n21158), .B(n21157), .Z(n21160) );
  XNOR U22145 ( .A(n21159), .B(n21160), .Z(n21161) );
  XNOR U22146 ( .A(n21162), .B(n21161), .Z(n21177) );
  XNOR U22147 ( .A(n21177), .B(sreg[1910]), .Z(n21179) );
  XNOR U22148 ( .A(n21178), .B(n21179), .Z(c[1910]) );
  NANDN U22149 ( .A(n21160), .B(n21159), .Z(n21164) );
  NAND U22150 ( .A(n21162), .B(n21161), .Z(n21163) );
  NAND U22151 ( .A(n21164), .B(n21163), .Z(n21186) );
  AND U22152 ( .A(b[2]), .B(a[889]), .Z(n21192) );
  AND U22153 ( .A(a[890]), .B(b[1]), .Z(n21190) );
  AND U22154 ( .A(a[888]), .B(b[3]), .Z(n21189) );
  XOR U22155 ( .A(n21190), .B(n21189), .Z(n21191) );
  XOR U22156 ( .A(n21192), .B(n21191), .Z(n21195) );
  NAND U22157 ( .A(b[0]), .B(a[891]), .Z(n21196) );
  XOR U22158 ( .A(n21195), .B(n21196), .Z(n21198) );
  OR U22159 ( .A(n21166), .B(n21165), .Z(n21170) );
  NANDN U22160 ( .A(n21168), .B(n21167), .Z(n21169) );
  NAND U22161 ( .A(n21170), .B(n21169), .Z(n21197) );
  XNOR U22162 ( .A(n21198), .B(n21197), .Z(n21183) );
  NANDN U22163 ( .A(n21172), .B(n21171), .Z(n21176) );
  OR U22164 ( .A(n21174), .B(n21173), .Z(n21175) );
  NAND U22165 ( .A(n21176), .B(n21175), .Z(n21184) );
  XNOR U22166 ( .A(n21183), .B(n21184), .Z(n21185) );
  XNOR U22167 ( .A(n21186), .B(n21185), .Z(n21202) );
  NAND U22168 ( .A(n21177), .B(sreg[1910]), .Z(n21181) );
  NANDN U22169 ( .A(n21179), .B(n21178), .Z(n21180) );
  AND U22170 ( .A(n21181), .B(n21180), .Z(n21201) );
  XNOR U22171 ( .A(n21201), .B(sreg[1911]), .Z(n21182) );
  XOR U22172 ( .A(n21202), .B(n21182), .Z(c[1911]) );
  NANDN U22173 ( .A(n21184), .B(n21183), .Z(n21188) );
  NAND U22174 ( .A(n21186), .B(n21185), .Z(n21187) );
  NAND U22175 ( .A(n21188), .B(n21187), .Z(n21209) );
  AND U22176 ( .A(b[2]), .B(a[890]), .Z(n21215) );
  AND U22177 ( .A(a[891]), .B(b[1]), .Z(n21213) );
  AND U22178 ( .A(a[889]), .B(b[3]), .Z(n21212) );
  XOR U22179 ( .A(n21213), .B(n21212), .Z(n21214) );
  XOR U22180 ( .A(n21215), .B(n21214), .Z(n21218) );
  NAND U22181 ( .A(b[0]), .B(a[892]), .Z(n21219) );
  XOR U22182 ( .A(n21218), .B(n21219), .Z(n21221) );
  OR U22183 ( .A(n21190), .B(n21189), .Z(n21194) );
  NANDN U22184 ( .A(n21192), .B(n21191), .Z(n21193) );
  NAND U22185 ( .A(n21194), .B(n21193), .Z(n21220) );
  XNOR U22186 ( .A(n21221), .B(n21220), .Z(n21206) );
  NANDN U22187 ( .A(n21196), .B(n21195), .Z(n21200) );
  OR U22188 ( .A(n21198), .B(n21197), .Z(n21199) );
  NAND U22189 ( .A(n21200), .B(n21199), .Z(n21207) );
  XNOR U22190 ( .A(n21206), .B(n21207), .Z(n21208) );
  XNOR U22191 ( .A(n21209), .B(n21208), .Z(n21205) );
  XOR U22192 ( .A(n21204), .B(sreg[1912]), .Z(n21203) );
  XOR U22193 ( .A(n21205), .B(n21203), .Z(c[1912]) );
  NANDN U22194 ( .A(n21207), .B(n21206), .Z(n21211) );
  NAND U22195 ( .A(n21209), .B(n21208), .Z(n21210) );
  NAND U22196 ( .A(n21211), .B(n21210), .Z(n21232) );
  AND U22197 ( .A(b[2]), .B(a[891]), .Z(n21238) );
  AND U22198 ( .A(a[892]), .B(b[1]), .Z(n21236) );
  AND U22199 ( .A(a[890]), .B(b[3]), .Z(n21235) );
  XOR U22200 ( .A(n21236), .B(n21235), .Z(n21237) );
  XOR U22201 ( .A(n21238), .B(n21237), .Z(n21241) );
  NAND U22202 ( .A(b[0]), .B(a[893]), .Z(n21242) );
  XOR U22203 ( .A(n21241), .B(n21242), .Z(n21244) );
  OR U22204 ( .A(n21213), .B(n21212), .Z(n21217) );
  NANDN U22205 ( .A(n21215), .B(n21214), .Z(n21216) );
  NAND U22206 ( .A(n21217), .B(n21216), .Z(n21243) );
  XNOR U22207 ( .A(n21244), .B(n21243), .Z(n21229) );
  NANDN U22208 ( .A(n21219), .B(n21218), .Z(n21223) );
  OR U22209 ( .A(n21221), .B(n21220), .Z(n21222) );
  NAND U22210 ( .A(n21223), .B(n21222), .Z(n21230) );
  XNOR U22211 ( .A(n21229), .B(n21230), .Z(n21231) );
  XNOR U22212 ( .A(n21232), .B(n21231), .Z(n21224) );
  XNOR U22213 ( .A(n21224), .B(sreg[1913]), .Z(n21226) );
  XNOR U22214 ( .A(n21225), .B(n21226), .Z(c[1913]) );
  NAND U22215 ( .A(n21224), .B(sreg[1913]), .Z(n21228) );
  NANDN U22216 ( .A(n21226), .B(n21225), .Z(n21227) );
  AND U22217 ( .A(n21228), .B(n21227), .Z(n21267) );
  NANDN U22218 ( .A(n21230), .B(n21229), .Z(n21234) );
  NAND U22219 ( .A(n21232), .B(n21231), .Z(n21233) );
  NAND U22220 ( .A(n21234), .B(n21233), .Z(n21251) );
  AND U22221 ( .A(b[2]), .B(a[892]), .Z(n21257) );
  AND U22222 ( .A(a[893]), .B(b[1]), .Z(n21255) );
  AND U22223 ( .A(a[891]), .B(b[3]), .Z(n21254) );
  XOR U22224 ( .A(n21255), .B(n21254), .Z(n21256) );
  XOR U22225 ( .A(n21257), .B(n21256), .Z(n21260) );
  NAND U22226 ( .A(b[0]), .B(a[894]), .Z(n21261) );
  XOR U22227 ( .A(n21260), .B(n21261), .Z(n21263) );
  OR U22228 ( .A(n21236), .B(n21235), .Z(n21240) );
  NANDN U22229 ( .A(n21238), .B(n21237), .Z(n21239) );
  NAND U22230 ( .A(n21240), .B(n21239), .Z(n21262) );
  XNOR U22231 ( .A(n21263), .B(n21262), .Z(n21248) );
  NANDN U22232 ( .A(n21242), .B(n21241), .Z(n21246) );
  OR U22233 ( .A(n21244), .B(n21243), .Z(n21245) );
  NAND U22234 ( .A(n21246), .B(n21245), .Z(n21249) );
  XNOR U22235 ( .A(n21248), .B(n21249), .Z(n21250) );
  XNOR U22236 ( .A(n21251), .B(n21250), .Z(n21266) );
  XNOR U22237 ( .A(sreg[1914]), .B(n21266), .Z(n21247) );
  XOR U22238 ( .A(n21267), .B(n21247), .Z(c[1914]) );
  NANDN U22239 ( .A(n21249), .B(n21248), .Z(n21253) );
  NAND U22240 ( .A(n21251), .B(n21250), .Z(n21252) );
  NAND U22241 ( .A(n21253), .B(n21252), .Z(n21272) );
  AND U22242 ( .A(b[2]), .B(a[893]), .Z(n21278) );
  AND U22243 ( .A(a[894]), .B(b[1]), .Z(n21276) );
  AND U22244 ( .A(a[892]), .B(b[3]), .Z(n21275) );
  XOR U22245 ( .A(n21276), .B(n21275), .Z(n21277) );
  XOR U22246 ( .A(n21278), .B(n21277), .Z(n21281) );
  NAND U22247 ( .A(b[0]), .B(a[895]), .Z(n21282) );
  XOR U22248 ( .A(n21281), .B(n21282), .Z(n21284) );
  OR U22249 ( .A(n21255), .B(n21254), .Z(n21259) );
  NANDN U22250 ( .A(n21257), .B(n21256), .Z(n21258) );
  NAND U22251 ( .A(n21259), .B(n21258), .Z(n21283) );
  XNOR U22252 ( .A(n21284), .B(n21283), .Z(n21269) );
  NANDN U22253 ( .A(n21261), .B(n21260), .Z(n21265) );
  OR U22254 ( .A(n21263), .B(n21262), .Z(n21264) );
  NAND U22255 ( .A(n21265), .B(n21264), .Z(n21270) );
  XNOR U22256 ( .A(n21269), .B(n21270), .Z(n21271) );
  XOR U22257 ( .A(n21272), .B(n21271), .Z(n21288) );
  XNOR U22258 ( .A(sreg[1915]), .B(n21287), .Z(n21268) );
  XOR U22259 ( .A(n21288), .B(n21268), .Z(c[1915]) );
  NANDN U22260 ( .A(n21270), .B(n21269), .Z(n21274) );
  NAND U22261 ( .A(n21272), .B(n21271), .Z(n21273) );
  NAND U22262 ( .A(n21274), .B(n21273), .Z(n21295) );
  AND U22263 ( .A(b[2]), .B(a[894]), .Z(n21301) );
  AND U22264 ( .A(a[895]), .B(b[1]), .Z(n21299) );
  AND U22265 ( .A(a[893]), .B(b[3]), .Z(n21298) );
  XOR U22266 ( .A(n21299), .B(n21298), .Z(n21300) );
  XOR U22267 ( .A(n21301), .B(n21300), .Z(n21304) );
  NAND U22268 ( .A(b[0]), .B(a[896]), .Z(n21305) );
  XOR U22269 ( .A(n21304), .B(n21305), .Z(n21307) );
  OR U22270 ( .A(n21276), .B(n21275), .Z(n21280) );
  NANDN U22271 ( .A(n21278), .B(n21277), .Z(n21279) );
  NAND U22272 ( .A(n21280), .B(n21279), .Z(n21306) );
  XNOR U22273 ( .A(n21307), .B(n21306), .Z(n21292) );
  NANDN U22274 ( .A(n21282), .B(n21281), .Z(n21286) );
  OR U22275 ( .A(n21284), .B(n21283), .Z(n21285) );
  NAND U22276 ( .A(n21286), .B(n21285), .Z(n21293) );
  XNOR U22277 ( .A(n21292), .B(n21293), .Z(n21294) );
  XOR U22278 ( .A(n21295), .B(n21294), .Z(n21291) );
  XNOR U22279 ( .A(sreg[1916]), .B(n21290), .Z(n21289) );
  XOR U22280 ( .A(n21291), .B(n21289), .Z(c[1916]) );
  NANDN U22281 ( .A(n21293), .B(n21292), .Z(n21297) );
  NAND U22282 ( .A(n21295), .B(n21294), .Z(n21296) );
  NAND U22283 ( .A(n21297), .B(n21296), .Z(n21313) );
  AND U22284 ( .A(b[2]), .B(a[895]), .Z(n21319) );
  AND U22285 ( .A(a[896]), .B(b[1]), .Z(n21317) );
  AND U22286 ( .A(a[894]), .B(b[3]), .Z(n21316) );
  XOR U22287 ( .A(n21317), .B(n21316), .Z(n21318) );
  XOR U22288 ( .A(n21319), .B(n21318), .Z(n21322) );
  NAND U22289 ( .A(b[0]), .B(a[897]), .Z(n21323) );
  XOR U22290 ( .A(n21322), .B(n21323), .Z(n21325) );
  OR U22291 ( .A(n21299), .B(n21298), .Z(n21303) );
  NANDN U22292 ( .A(n21301), .B(n21300), .Z(n21302) );
  NAND U22293 ( .A(n21303), .B(n21302), .Z(n21324) );
  XNOR U22294 ( .A(n21325), .B(n21324), .Z(n21310) );
  NANDN U22295 ( .A(n21305), .B(n21304), .Z(n21309) );
  OR U22296 ( .A(n21307), .B(n21306), .Z(n21308) );
  NAND U22297 ( .A(n21309), .B(n21308), .Z(n21311) );
  XNOR U22298 ( .A(n21310), .B(n21311), .Z(n21312) );
  XNOR U22299 ( .A(n21313), .B(n21312), .Z(n21328) );
  XNOR U22300 ( .A(n21328), .B(sreg[1917]), .Z(n21329) );
  XOR U22301 ( .A(n21330), .B(n21329), .Z(c[1917]) );
  NANDN U22302 ( .A(n21311), .B(n21310), .Z(n21315) );
  NAND U22303 ( .A(n21313), .B(n21312), .Z(n21314) );
  NAND U22304 ( .A(n21315), .B(n21314), .Z(n21339) );
  AND U22305 ( .A(b[2]), .B(a[896]), .Z(n21345) );
  AND U22306 ( .A(a[897]), .B(b[1]), .Z(n21343) );
  AND U22307 ( .A(a[895]), .B(b[3]), .Z(n21342) );
  XOR U22308 ( .A(n21343), .B(n21342), .Z(n21344) );
  XOR U22309 ( .A(n21345), .B(n21344), .Z(n21348) );
  NAND U22310 ( .A(b[0]), .B(a[898]), .Z(n21349) );
  XOR U22311 ( .A(n21348), .B(n21349), .Z(n21351) );
  OR U22312 ( .A(n21317), .B(n21316), .Z(n21321) );
  NANDN U22313 ( .A(n21319), .B(n21318), .Z(n21320) );
  NAND U22314 ( .A(n21321), .B(n21320), .Z(n21350) );
  XNOR U22315 ( .A(n21351), .B(n21350), .Z(n21336) );
  NANDN U22316 ( .A(n21323), .B(n21322), .Z(n21327) );
  OR U22317 ( .A(n21325), .B(n21324), .Z(n21326) );
  NAND U22318 ( .A(n21327), .B(n21326), .Z(n21337) );
  XNOR U22319 ( .A(n21336), .B(n21337), .Z(n21338) );
  XOR U22320 ( .A(n21339), .B(n21338), .Z(n21335) );
  NAND U22321 ( .A(n21328), .B(sreg[1917]), .Z(n21332) );
  OR U22322 ( .A(n21330), .B(n21329), .Z(n21331) );
  NAND U22323 ( .A(n21332), .B(n21331), .Z(n21334) );
  XNOR U22324 ( .A(sreg[1918]), .B(n21334), .Z(n21333) );
  XOR U22325 ( .A(n21335), .B(n21333), .Z(c[1918]) );
  NANDN U22326 ( .A(n21337), .B(n21336), .Z(n21341) );
  NAND U22327 ( .A(n21339), .B(n21338), .Z(n21340) );
  NAND U22328 ( .A(n21341), .B(n21340), .Z(n21357) );
  AND U22329 ( .A(b[2]), .B(a[897]), .Z(n21363) );
  AND U22330 ( .A(a[898]), .B(b[1]), .Z(n21361) );
  AND U22331 ( .A(a[896]), .B(b[3]), .Z(n21360) );
  XOR U22332 ( .A(n21361), .B(n21360), .Z(n21362) );
  XOR U22333 ( .A(n21363), .B(n21362), .Z(n21366) );
  NAND U22334 ( .A(b[0]), .B(a[899]), .Z(n21367) );
  XOR U22335 ( .A(n21366), .B(n21367), .Z(n21369) );
  OR U22336 ( .A(n21343), .B(n21342), .Z(n21347) );
  NANDN U22337 ( .A(n21345), .B(n21344), .Z(n21346) );
  NAND U22338 ( .A(n21347), .B(n21346), .Z(n21368) );
  XNOR U22339 ( .A(n21369), .B(n21368), .Z(n21354) );
  NANDN U22340 ( .A(n21349), .B(n21348), .Z(n21353) );
  OR U22341 ( .A(n21351), .B(n21350), .Z(n21352) );
  NAND U22342 ( .A(n21353), .B(n21352), .Z(n21355) );
  XNOR U22343 ( .A(n21354), .B(n21355), .Z(n21356) );
  XNOR U22344 ( .A(n21357), .B(n21356), .Z(n21372) );
  XNOR U22345 ( .A(n21372), .B(sreg[1919]), .Z(n21373) );
  XOR U22346 ( .A(n21374), .B(n21373), .Z(c[1919]) );
  NANDN U22347 ( .A(n21355), .B(n21354), .Z(n21359) );
  NAND U22348 ( .A(n21357), .B(n21356), .Z(n21358) );
  NAND U22349 ( .A(n21359), .B(n21358), .Z(n21380) );
  AND U22350 ( .A(b[2]), .B(a[898]), .Z(n21386) );
  AND U22351 ( .A(a[899]), .B(b[1]), .Z(n21384) );
  AND U22352 ( .A(a[897]), .B(b[3]), .Z(n21383) );
  XOR U22353 ( .A(n21384), .B(n21383), .Z(n21385) );
  XOR U22354 ( .A(n21386), .B(n21385), .Z(n21389) );
  NAND U22355 ( .A(b[0]), .B(a[900]), .Z(n21390) );
  XOR U22356 ( .A(n21389), .B(n21390), .Z(n21392) );
  OR U22357 ( .A(n21361), .B(n21360), .Z(n21365) );
  NANDN U22358 ( .A(n21363), .B(n21362), .Z(n21364) );
  NAND U22359 ( .A(n21365), .B(n21364), .Z(n21391) );
  XNOR U22360 ( .A(n21392), .B(n21391), .Z(n21377) );
  NANDN U22361 ( .A(n21367), .B(n21366), .Z(n21371) );
  OR U22362 ( .A(n21369), .B(n21368), .Z(n21370) );
  NAND U22363 ( .A(n21371), .B(n21370), .Z(n21378) );
  XNOR U22364 ( .A(n21377), .B(n21378), .Z(n21379) );
  XNOR U22365 ( .A(n21380), .B(n21379), .Z(n21395) );
  XNOR U22366 ( .A(n21395), .B(sreg[1920]), .Z(n21397) );
  NAND U22367 ( .A(n21372), .B(sreg[1919]), .Z(n21376) );
  OR U22368 ( .A(n21374), .B(n21373), .Z(n21375) );
  AND U22369 ( .A(n21376), .B(n21375), .Z(n21396) );
  XOR U22370 ( .A(n21397), .B(n21396), .Z(c[1920]) );
  NANDN U22371 ( .A(n21378), .B(n21377), .Z(n21382) );
  NAND U22372 ( .A(n21380), .B(n21379), .Z(n21381) );
  NAND U22373 ( .A(n21382), .B(n21381), .Z(n21404) );
  AND U22374 ( .A(b[2]), .B(a[899]), .Z(n21410) );
  AND U22375 ( .A(a[900]), .B(b[1]), .Z(n21408) );
  AND U22376 ( .A(a[898]), .B(b[3]), .Z(n21407) );
  XOR U22377 ( .A(n21408), .B(n21407), .Z(n21409) );
  XOR U22378 ( .A(n21410), .B(n21409), .Z(n21413) );
  NAND U22379 ( .A(b[0]), .B(a[901]), .Z(n21414) );
  XOR U22380 ( .A(n21413), .B(n21414), .Z(n21416) );
  OR U22381 ( .A(n21384), .B(n21383), .Z(n21388) );
  NANDN U22382 ( .A(n21386), .B(n21385), .Z(n21387) );
  NAND U22383 ( .A(n21388), .B(n21387), .Z(n21415) );
  XNOR U22384 ( .A(n21416), .B(n21415), .Z(n21401) );
  NANDN U22385 ( .A(n21390), .B(n21389), .Z(n21394) );
  OR U22386 ( .A(n21392), .B(n21391), .Z(n21393) );
  NAND U22387 ( .A(n21394), .B(n21393), .Z(n21402) );
  XNOR U22388 ( .A(n21401), .B(n21402), .Z(n21403) );
  XOR U22389 ( .A(n21404), .B(n21403), .Z(n21420) );
  NAND U22390 ( .A(n21395), .B(sreg[1920]), .Z(n21399) );
  OR U22391 ( .A(n21397), .B(n21396), .Z(n21398) );
  NAND U22392 ( .A(n21399), .B(n21398), .Z(n21419) );
  XNOR U22393 ( .A(sreg[1921]), .B(n21419), .Z(n21400) );
  XOR U22394 ( .A(n21420), .B(n21400), .Z(c[1921]) );
  NANDN U22395 ( .A(n21402), .B(n21401), .Z(n21406) );
  NAND U22396 ( .A(n21404), .B(n21403), .Z(n21405) );
  NAND U22397 ( .A(n21406), .B(n21405), .Z(n21437) );
  AND U22398 ( .A(b[2]), .B(a[900]), .Z(n21431) );
  AND U22399 ( .A(a[901]), .B(b[1]), .Z(n21429) );
  AND U22400 ( .A(a[899]), .B(b[3]), .Z(n21428) );
  XOR U22401 ( .A(n21429), .B(n21428), .Z(n21430) );
  XOR U22402 ( .A(n21431), .B(n21430), .Z(n21422) );
  NAND U22403 ( .A(b[0]), .B(a[902]), .Z(n21423) );
  XOR U22404 ( .A(n21422), .B(n21423), .Z(n21425) );
  OR U22405 ( .A(n21408), .B(n21407), .Z(n21412) );
  NANDN U22406 ( .A(n21410), .B(n21409), .Z(n21411) );
  NAND U22407 ( .A(n21412), .B(n21411), .Z(n21424) );
  XNOR U22408 ( .A(n21425), .B(n21424), .Z(n21434) );
  NANDN U22409 ( .A(n21414), .B(n21413), .Z(n21418) );
  OR U22410 ( .A(n21416), .B(n21415), .Z(n21417) );
  NAND U22411 ( .A(n21418), .B(n21417), .Z(n21435) );
  XNOR U22412 ( .A(n21434), .B(n21435), .Z(n21436) );
  XOR U22413 ( .A(n21437), .B(n21436), .Z(n21441) );
  XNOR U22414 ( .A(sreg[1922]), .B(n21440), .Z(n21421) );
  XOR U22415 ( .A(n21441), .B(n21421), .Z(c[1922]) );
  NANDN U22416 ( .A(n21423), .B(n21422), .Z(n21427) );
  OR U22417 ( .A(n21425), .B(n21424), .Z(n21426) );
  NAND U22418 ( .A(n21427), .B(n21426), .Z(n21445) );
  AND U22419 ( .A(b[2]), .B(a[901]), .Z(n21454) );
  AND U22420 ( .A(a[902]), .B(b[1]), .Z(n21452) );
  AND U22421 ( .A(a[900]), .B(b[3]), .Z(n21451) );
  XOR U22422 ( .A(n21452), .B(n21451), .Z(n21453) );
  XOR U22423 ( .A(n21454), .B(n21453), .Z(n21457) );
  NAND U22424 ( .A(b[0]), .B(a[903]), .Z(n21458) );
  XNOR U22425 ( .A(n21457), .B(n21458), .Z(n21459) );
  OR U22426 ( .A(n21429), .B(n21428), .Z(n21433) );
  NANDN U22427 ( .A(n21431), .B(n21430), .Z(n21432) );
  AND U22428 ( .A(n21433), .B(n21432), .Z(n21460) );
  XNOR U22429 ( .A(n21459), .B(n21460), .Z(n21446) );
  XNOR U22430 ( .A(n21445), .B(n21446), .Z(n21447) );
  NANDN U22431 ( .A(n21435), .B(n21434), .Z(n21439) );
  NAND U22432 ( .A(n21437), .B(n21436), .Z(n21438) );
  AND U22433 ( .A(n21439), .B(n21438), .Z(n21448) );
  XNOR U22434 ( .A(n21447), .B(n21448), .Z(n21444) );
  XNOR U22435 ( .A(sreg[1923]), .B(n21443), .Z(n21442) );
  XOR U22436 ( .A(n21444), .B(n21442), .Z(c[1923]) );
  NANDN U22437 ( .A(n21446), .B(n21445), .Z(n21450) );
  NAND U22438 ( .A(n21448), .B(n21447), .Z(n21449) );
  NAND U22439 ( .A(n21450), .B(n21449), .Z(n21466) );
  AND U22440 ( .A(b[2]), .B(a[902]), .Z(n21472) );
  AND U22441 ( .A(a[903]), .B(b[1]), .Z(n21470) );
  AND U22442 ( .A(a[901]), .B(b[3]), .Z(n21469) );
  XOR U22443 ( .A(n21470), .B(n21469), .Z(n21471) );
  XOR U22444 ( .A(n21472), .B(n21471), .Z(n21475) );
  NAND U22445 ( .A(b[0]), .B(a[904]), .Z(n21476) );
  XOR U22446 ( .A(n21475), .B(n21476), .Z(n21478) );
  OR U22447 ( .A(n21452), .B(n21451), .Z(n21456) );
  NANDN U22448 ( .A(n21454), .B(n21453), .Z(n21455) );
  NAND U22449 ( .A(n21456), .B(n21455), .Z(n21477) );
  XNOR U22450 ( .A(n21478), .B(n21477), .Z(n21463) );
  NANDN U22451 ( .A(n21458), .B(n21457), .Z(n21462) );
  NAND U22452 ( .A(n21460), .B(n21459), .Z(n21461) );
  NAND U22453 ( .A(n21462), .B(n21461), .Z(n21464) );
  XNOR U22454 ( .A(n21463), .B(n21464), .Z(n21465) );
  XOR U22455 ( .A(n21466), .B(n21465), .Z(n21481) );
  XNOR U22456 ( .A(n21481), .B(sreg[1924]), .Z(n21482) );
  XOR U22457 ( .A(n21483), .B(n21482), .Z(c[1924]) );
  NANDN U22458 ( .A(n21464), .B(n21463), .Z(n21468) );
  NANDN U22459 ( .A(n21466), .B(n21465), .Z(n21467) );
  NAND U22460 ( .A(n21468), .B(n21467), .Z(n21502) );
  AND U22461 ( .A(b[2]), .B(a[903]), .Z(n21496) );
  AND U22462 ( .A(a[904]), .B(b[1]), .Z(n21494) );
  AND U22463 ( .A(a[902]), .B(b[3]), .Z(n21493) );
  XOR U22464 ( .A(n21494), .B(n21493), .Z(n21495) );
  XOR U22465 ( .A(n21496), .B(n21495), .Z(n21487) );
  NAND U22466 ( .A(b[0]), .B(a[905]), .Z(n21488) );
  XOR U22467 ( .A(n21487), .B(n21488), .Z(n21490) );
  OR U22468 ( .A(n21470), .B(n21469), .Z(n21474) );
  NANDN U22469 ( .A(n21472), .B(n21471), .Z(n21473) );
  NAND U22470 ( .A(n21474), .B(n21473), .Z(n21489) );
  XNOR U22471 ( .A(n21490), .B(n21489), .Z(n21499) );
  NANDN U22472 ( .A(n21476), .B(n21475), .Z(n21480) );
  OR U22473 ( .A(n21478), .B(n21477), .Z(n21479) );
  NAND U22474 ( .A(n21480), .B(n21479), .Z(n21500) );
  XNOR U22475 ( .A(n21499), .B(n21500), .Z(n21501) );
  XNOR U22476 ( .A(n21502), .B(n21501), .Z(n21506) );
  NAND U22477 ( .A(n21481), .B(sreg[1924]), .Z(n21485) );
  OR U22478 ( .A(n21483), .B(n21482), .Z(n21484) );
  AND U22479 ( .A(n21485), .B(n21484), .Z(n21505) );
  XNOR U22480 ( .A(n21505), .B(sreg[1925]), .Z(n21486) );
  XOR U22481 ( .A(n21506), .B(n21486), .Z(c[1925]) );
  NANDN U22482 ( .A(n21488), .B(n21487), .Z(n21492) );
  OR U22483 ( .A(n21490), .B(n21489), .Z(n21491) );
  NAND U22484 ( .A(n21492), .B(n21491), .Z(n21508) );
  AND U22485 ( .A(b[2]), .B(a[904]), .Z(n21517) );
  AND U22486 ( .A(a[905]), .B(b[1]), .Z(n21515) );
  AND U22487 ( .A(a[903]), .B(b[3]), .Z(n21514) );
  XOR U22488 ( .A(n21515), .B(n21514), .Z(n21516) );
  XOR U22489 ( .A(n21517), .B(n21516), .Z(n21520) );
  NAND U22490 ( .A(b[0]), .B(a[906]), .Z(n21521) );
  XNOR U22491 ( .A(n21520), .B(n21521), .Z(n21522) );
  OR U22492 ( .A(n21494), .B(n21493), .Z(n21498) );
  NANDN U22493 ( .A(n21496), .B(n21495), .Z(n21497) );
  AND U22494 ( .A(n21498), .B(n21497), .Z(n21523) );
  XNOR U22495 ( .A(n21522), .B(n21523), .Z(n21509) );
  XNOR U22496 ( .A(n21508), .B(n21509), .Z(n21510) );
  NANDN U22497 ( .A(n21500), .B(n21499), .Z(n21504) );
  NAND U22498 ( .A(n21502), .B(n21501), .Z(n21503) );
  AND U22499 ( .A(n21504), .B(n21503), .Z(n21511) );
  XNOR U22500 ( .A(n21510), .B(n21511), .Z(n21527) );
  XNOR U22501 ( .A(n21526), .B(sreg[1926]), .Z(n21507) );
  XOR U22502 ( .A(n21527), .B(n21507), .Z(c[1926]) );
  NANDN U22503 ( .A(n21509), .B(n21508), .Z(n21513) );
  NAND U22504 ( .A(n21511), .B(n21510), .Z(n21512) );
  NAND U22505 ( .A(n21513), .B(n21512), .Z(n21532) );
  AND U22506 ( .A(b[2]), .B(a[905]), .Z(n21538) );
  AND U22507 ( .A(a[906]), .B(b[1]), .Z(n21536) );
  AND U22508 ( .A(a[904]), .B(b[3]), .Z(n21535) );
  XOR U22509 ( .A(n21536), .B(n21535), .Z(n21537) );
  XOR U22510 ( .A(n21538), .B(n21537), .Z(n21541) );
  NAND U22511 ( .A(b[0]), .B(a[907]), .Z(n21542) );
  XOR U22512 ( .A(n21541), .B(n21542), .Z(n21544) );
  OR U22513 ( .A(n21515), .B(n21514), .Z(n21519) );
  NANDN U22514 ( .A(n21517), .B(n21516), .Z(n21518) );
  NAND U22515 ( .A(n21519), .B(n21518), .Z(n21543) );
  XNOR U22516 ( .A(n21544), .B(n21543), .Z(n21529) );
  NANDN U22517 ( .A(n21521), .B(n21520), .Z(n21525) );
  NAND U22518 ( .A(n21523), .B(n21522), .Z(n21524) );
  NAND U22519 ( .A(n21525), .B(n21524), .Z(n21530) );
  XNOR U22520 ( .A(n21529), .B(n21530), .Z(n21531) );
  XNOR U22521 ( .A(n21532), .B(n21531), .Z(n21548) );
  XNOR U22522 ( .A(n21547), .B(sreg[1927]), .Z(n21528) );
  XNOR U22523 ( .A(n21548), .B(n21528), .Z(c[1927]) );
  NANDN U22524 ( .A(n21530), .B(n21529), .Z(n21534) );
  NANDN U22525 ( .A(n21532), .B(n21531), .Z(n21533) );
  NAND U22526 ( .A(n21534), .B(n21533), .Z(n21565) );
  AND U22527 ( .A(b[2]), .B(a[906]), .Z(n21559) );
  AND U22528 ( .A(a[907]), .B(b[1]), .Z(n21557) );
  AND U22529 ( .A(a[905]), .B(b[3]), .Z(n21556) );
  XOR U22530 ( .A(n21557), .B(n21556), .Z(n21558) );
  XOR U22531 ( .A(n21559), .B(n21558), .Z(n21550) );
  NAND U22532 ( .A(b[0]), .B(a[908]), .Z(n21551) );
  XOR U22533 ( .A(n21550), .B(n21551), .Z(n21553) );
  OR U22534 ( .A(n21536), .B(n21535), .Z(n21540) );
  NANDN U22535 ( .A(n21538), .B(n21537), .Z(n21539) );
  NAND U22536 ( .A(n21540), .B(n21539), .Z(n21552) );
  XNOR U22537 ( .A(n21553), .B(n21552), .Z(n21562) );
  NANDN U22538 ( .A(n21542), .B(n21541), .Z(n21546) );
  OR U22539 ( .A(n21544), .B(n21543), .Z(n21545) );
  NAND U22540 ( .A(n21546), .B(n21545), .Z(n21563) );
  XNOR U22541 ( .A(n21562), .B(n21563), .Z(n21564) );
  XOR U22542 ( .A(n21565), .B(n21564), .Z(n21569) );
  XOR U22543 ( .A(sreg[1928]), .B(n21568), .Z(n21549) );
  XOR U22544 ( .A(n21569), .B(n21549), .Z(c[1928]) );
  NANDN U22545 ( .A(n21551), .B(n21550), .Z(n21555) );
  OR U22546 ( .A(n21553), .B(n21552), .Z(n21554) );
  NAND U22547 ( .A(n21555), .B(n21554), .Z(n21573) );
  AND U22548 ( .A(b[2]), .B(a[907]), .Z(n21582) );
  AND U22549 ( .A(a[908]), .B(b[1]), .Z(n21580) );
  AND U22550 ( .A(a[906]), .B(b[3]), .Z(n21579) );
  XOR U22551 ( .A(n21580), .B(n21579), .Z(n21581) );
  XOR U22552 ( .A(n21582), .B(n21581), .Z(n21585) );
  NAND U22553 ( .A(b[0]), .B(a[909]), .Z(n21586) );
  XNOR U22554 ( .A(n21585), .B(n21586), .Z(n21587) );
  OR U22555 ( .A(n21557), .B(n21556), .Z(n21561) );
  NANDN U22556 ( .A(n21559), .B(n21558), .Z(n21560) );
  AND U22557 ( .A(n21561), .B(n21560), .Z(n21588) );
  XNOR U22558 ( .A(n21587), .B(n21588), .Z(n21574) );
  XNOR U22559 ( .A(n21573), .B(n21574), .Z(n21575) );
  NANDN U22560 ( .A(n21563), .B(n21562), .Z(n21567) );
  NAND U22561 ( .A(n21565), .B(n21564), .Z(n21566) );
  NAND U22562 ( .A(n21567), .B(n21566), .Z(n21576) );
  XOR U22563 ( .A(n21575), .B(n21576), .Z(n21572) );
  XOR U22564 ( .A(n21571), .B(sreg[1929]), .Z(n21570) );
  XNOR U22565 ( .A(n21572), .B(n21570), .Z(c[1929]) );
  NANDN U22566 ( .A(n21574), .B(n21573), .Z(n21578) );
  NANDN U22567 ( .A(n21576), .B(n21575), .Z(n21577) );
  NAND U22568 ( .A(n21578), .B(n21577), .Z(n21594) );
  AND U22569 ( .A(b[2]), .B(a[908]), .Z(n21600) );
  AND U22570 ( .A(a[909]), .B(b[1]), .Z(n21598) );
  AND U22571 ( .A(a[907]), .B(b[3]), .Z(n21597) );
  XOR U22572 ( .A(n21598), .B(n21597), .Z(n21599) );
  XOR U22573 ( .A(n21600), .B(n21599), .Z(n21603) );
  NAND U22574 ( .A(b[0]), .B(a[910]), .Z(n21604) );
  XOR U22575 ( .A(n21603), .B(n21604), .Z(n21606) );
  OR U22576 ( .A(n21580), .B(n21579), .Z(n21584) );
  NANDN U22577 ( .A(n21582), .B(n21581), .Z(n21583) );
  NAND U22578 ( .A(n21584), .B(n21583), .Z(n21605) );
  XNOR U22579 ( .A(n21606), .B(n21605), .Z(n21591) );
  NANDN U22580 ( .A(n21586), .B(n21585), .Z(n21590) );
  NAND U22581 ( .A(n21588), .B(n21587), .Z(n21589) );
  NAND U22582 ( .A(n21590), .B(n21589), .Z(n21592) );
  XNOR U22583 ( .A(n21591), .B(n21592), .Z(n21593) );
  XOR U22584 ( .A(n21594), .B(n21593), .Z(n21609) );
  XNOR U22585 ( .A(n21609), .B(sreg[1930]), .Z(n21611) );
  XNOR U22586 ( .A(n21610), .B(n21611), .Z(c[1930]) );
  NANDN U22587 ( .A(n21592), .B(n21591), .Z(n21596) );
  NANDN U22588 ( .A(n21594), .B(n21593), .Z(n21595) );
  NAND U22589 ( .A(n21596), .B(n21595), .Z(n21617) );
  AND U22590 ( .A(b[2]), .B(a[909]), .Z(n21623) );
  AND U22591 ( .A(a[910]), .B(b[1]), .Z(n21621) );
  AND U22592 ( .A(a[908]), .B(b[3]), .Z(n21620) );
  XOR U22593 ( .A(n21621), .B(n21620), .Z(n21622) );
  XOR U22594 ( .A(n21623), .B(n21622), .Z(n21626) );
  NAND U22595 ( .A(b[0]), .B(a[911]), .Z(n21627) );
  XOR U22596 ( .A(n21626), .B(n21627), .Z(n21629) );
  OR U22597 ( .A(n21598), .B(n21597), .Z(n21602) );
  NANDN U22598 ( .A(n21600), .B(n21599), .Z(n21601) );
  NAND U22599 ( .A(n21602), .B(n21601), .Z(n21628) );
  XNOR U22600 ( .A(n21629), .B(n21628), .Z(n21614) );
  NANDN U22601 ( .A(n21604), .B(n21603), .Z(n21608) );
  OR U22602 ( .A(n21606), .B(n21605), .Z(n21607) );
  NAND U22603 ( .A(n21608), .B(n21607), .Z(n21615) );
  XNOR U22604 ( .A(n21614), .B(n21615), .Z(n21616) );
  XNOR U22605 ( .A(n21617), .B(n21616), .Z(n21632) );
  XNOR U22606 ( .A(n21632), .B(sreg[1931]), .Z(n21634) );
  NAND U22607 ( .A(n21609), .B(sreg[1930]), .Z(n21613) );
  NANDN U22608 ( .A(n21611), .B(n21610), .Z(n21612) );
  AND U22609 ( .A(n21613), .B(n21612), .Z(n21633) );
  XOR U22610 ( .A(n21634), .B(n21633), .Z(c[1931]) );
  NANDN U22611 ( .A(n21615), .B(n21614), .Z(n21619) );
  NAND U22612 ( .A(n21617), .B(n21616), .Z(n21618) );
  NAND U22613 ( .A(n21619), .B(n21618), .Z(n21643) );
  AND U22614 ( .A(b[2]), .B(a[910]), .Z(n21649) );
  AND U22615 ( .A(a[911]), .B(b[1]), .Z(n21647) );
  AND U22616 ( .A(a[909]), .B(b[3]), .Z(n21646) );
  XOR U22617 ( .A(n21647), .B(n21646), .Z(n21648) );
  XOR U22618 ( .A(n21649), .B(n21648), .Z(n21652) );
  NAND U22619 ( .A(b[0]), .B(a[912]), .Z(n21653) );
  XOR U22620 ( .A(n21652), .B(n21653), .Z(n21655) );
  OR U22621 ( .A(n21621), .B(n21620), .Z(n21625) );
  NANDN U22622 ( .A(n21623), .B(n21622), .Z(n21624) );
  NAND U22623 ( .A(n21625), .B(n21624), .Z(n21654) );
  XNOR U22624 ( .A(n21655), .B(n21654), .Z(n21640) );
  NANDN U22625 ( .A(n21627), .B(n21626), .Z(n21631) );
  OR U22626 ( .A(n21629), .B(n21628), .Z(n21630) );
  NAND U22627 ( .A(n21631), .B(n21630), .Z(n21641) );
  XNOR U22628 ( .A(n21640), .B(n21641), .Z(n21642) );
  XOR U22629 ( .A(n21643), .B(n21642), .Z(n21639) );
  NAND U22630 ( .A(n21632), .B(sreg[1931]), .Z(n21636) );
  OR U22631 ( .A(n21634), .B(n21633), .Z(n21635) );
  NAND U22632 ( .A(n21636), .B(n21635), .Z(n21638) );
  XNOR U22633 ( .A(sreg[1932]), .B(n21638), .Z(n21637) );
  XOR U22634 ( .A(n21639), .B(n21637), .Z(c[1932]) );
  NANDN U22635 ( .A(n21641), .B(n21640), .Z(n21645) );
  NAND U22636 ( .A(n21643), .B(n21642), .Z(n21644) );
  NAND U22637 ( .A(n21645), .B(n21644), .Z(n21661) );
  AND U22638 ( .A(b[2]), .B(a[911]), .Z(n21673) );
  AND U22639 ( .A(a[912]), .B(b[1]), .Z(n21671) );
  AND U22640 ( .A(a[910]), .B(b[3]), .Z(n21670) );
  XOR U22641 ( .A(n21671), .B(n21670), .Z(n21672) );
  XOR U22642 ( .A(n21673), .B(n21672), .Z(n21664) );
  NAND U22643 ( .A(b[0]), .B(a[913]), .Z(n21665) );
  XOR U22644 ( .A(n21664), .B(n21665), .Z(n21667) );
  OR U22645 ( .A(n21647), .B(n21646), .Z(n21651) );
  NANDN U22646 ( .A(n21649), .B(n21648), .Z(n21650) );
  NAND U22647 ( .A(n21651), .B(n21650), .Z(n21666) );
  XNOR U22648 ( .A(n21667), .B(n21666), .Z(n21658) );
  NANDN U22649 ( .A(n21653), .B(n21652), .Z(n21657) );
  OR U22650 ( .A(n21655), .B(n21654), .Z(n21656) );
  NAND U22651 ( .A(n21657), .B(n21656), .Z(n21659) );
  XNOR U22652 ( .A(n21658), .B(n21659), .Z(n21660) );
  XNOR U22653 ( .A(n21661), .B(n21660), .Z(n21677) );
  XNOR U22654 ( .A(n21677), .B(sreg[1933]), .Z(n21678) );
  XOR U22655 ( .A(n21679), .B(n21678), .Z(c[1933]) );
  NANDN U22656 ( .A(n21659), .B(n21658), .Z(n21663) );
  NAND U22657 ( .A(n21661), .B(n21660), .Z(n21662) );
  AND U22658 ( .A(n21663), .B(n21662), .Z(n21684) );
  NANDN U22659 ( .A(n21665), .B(n21664), .Z(n21669) );
  OR U22660 ( .A(n21667), .B(n21666), .Z(n21668) );
  AND U22661 ( .A(n21669), .B(n21668), .Z(n21683) );
  AND U22662 ( .A(b[2]), .B(a[912]), .Z(n21688) );
  AND U22663 ( .A(a[913]), .B(b[1]), .Z(n21686) );
  AND U22664 ( .A(a[911]), .B(b[3]), .Z(n21685) );
  XOR U22665 ( .A(n21686), .B(n21685), .Z(n21687) );
  XOR U22666 ( .A(n21688), .B(n21687), .Z(n21691) );
  NAND U22667 ( .A(b[0]), .B(a[914]), .Z(n21692) );
  XOR U22668 ( .A(n21691), .B(n21692), .Z(n21694) );
  OR U22669 ( .A(n21671), .B(n21670), .Z(n21675) );
  NANDN U22670 ( .A(n21673), .B(n21672), .Z(n21674) );
  NAND U22671 ( .A(n21675), .B(n21674), .Z(n21693) );
  XOR U22672 ( .A(n21694), .B(n21693), .Z(n21682) );
  XNOR U22673 ( .A(n21683), .B(n21682), .Z(n21676) );
  XOR U22674 ( .A(n21684), .B(n21676), .Z(n21697) );
  XNOR U22675 ( .A(sreg[1934]), .B(n21697), .Z(n21699) );
  NAND U22676 ( .A(n21677), .B(sreg[1933]), .Z(n21681) );
  OR U22677 ( .A(n21679), .B(n21678), .Z(n21680) );
  AND U22678 ( .A(n21681), .B(n21680), .Z(n21698) );
  XOR U22679 ( .A(n21699), .B(n21698), .Z(c[1934]) );
  AND U22680 ( .A(b[2]), .B(a[913]), .Z(n21711) );
  AND U22681 ( .A(a[914]), .B(b[1]), .Z(n21709) );
  AND U22682 ( .A(a[912]), .B(b[3]), .Z(n21708) );
  XOR U22683 ( .A(n21709), .B(n21708), .Z(n21710) );
  XOR U22684 ( .A(n21711), .B(n21710), .Z(n21714) );
  NAND U22685 ( .A(b[0]), .B(a[915]), .Z(n21715) );
  XOR U22686 ( .A(n21714), .B(n21715), .Z(n21717) );
  OR U22687 ( .A(n21686), .B(n21685), .Z(n21690) );
  NANDN U22688 ( .A(n21688), .B(n21687), .Z(n21689) );
  NAND U22689 ( .A(n21690), .B(n21689), .Z(n21716) );
  XNOR U22690 ( .A(n21717), .B(n21716), .Z(n21702) );
  NANDN U22691 ( .A(n21692), .B(n21691), .Z(n21696) );
  OR U22692 ( .A(n21694), .B(n21693), .Z(n21695) );
  NAND U22693 ( .A(n21696), .B(n21695), .Z(n21703) );
  XNOR U22694 ( .A(n21702), .B(n21703), .Z(n21704) );
  XOR U22695 ( .A(n21705), .B(n21704), .Z(n21720) );
  XNOR U22696 ( .A(n21720), .B(sreg[1935]), .Z(n21722) );
  NAND U22697 ( .A(sreg[1934]), .B(n21697), .Z(n21701) );
  OR U22698 ( .A(n21699), .B(n21698), .Z(n21700) );
  AND U22699 ( .A(n21701), .B(n21700), .Z(n21721) );
  XOR U22700 ( .A(n21722), .B(n21721), .Z(c[1935]) );
  NANDN U22701 ( .A(n21703), .B(n21702), .Z(n21707) );
  NANDN U22702 ( .A(n21705), .B(n21704), .Z(n21706) );
  NAND U22703 ( .A(n21707), .B(n21706), .Z(n21728) );
  AND U22704 ( .A(b[2]), .B(a[914]), .Z(n21740) );
  AND U22705 ( .A(a[915]), .B(b[1]), .Z(n21738) );
  AND U22706 ( .A(a[913]), .B(b[3]), .Z(n21737) );
  XOR U22707 ( .A(n21738), .B(n21737), .Z(n21739) );
  XOR U22708 ( .A(n21740), .B(n21739), .Z(n21731) );
  NAND U22709 ( .A(b[0]), .B(a[916]), .Z(n21732) );
  XOR U22710 ( .A(n21731), .B(n21732), .Z(n21734) );
  OR U22711 ( .A(n21709), .B(n21708), .Z(n21713) );
  NANDN U22712 ( .A(n21711), .B(n21710), .Z(n21712) );
  NAND U22713 ( .A(n21713), .B(n21712), .Z(n21733) );
  XNOR U22714 ( .A(n21734), .B(n21733), .Z(n21725) );
  NANDN U22715 ( .A(n21715), .B(n21714), .Z(n21719) );
  OR U22716 ( .A(n21717), .B(n21716), .Z(n21718) );
  NAND U22717 ( .A(n21719), .B(n21718), .Z(n21726) );
  XNOR U22718 ( .A(n21725), .B(n21726), .Z(n21727) );
  XNOR U22719 ( .A(n21728), .B(n21727), .Z(n21743) );
  XOR U22720 ( .A(sreg[1936]), .B(n21743), .Z(n21744) );
  NAND U22721 ( .A(n21720), .B(sreg[1935]), .Z(n21724) );
  OR U22722 ( .A(n21722), .B(n21721), .Z(n21723) );
  NAND U22723 ( .A(n21724), .B(n21723), .Z(n21745) );
  XOR U22724 ( .A(n21744), .B(n21745), .Z(c[1936]) );
  NANDN U22725 ( .A(n21726), .B(n21725), .Z(n21730) );
  NAND U22726 ( .A(n21728), .B(n21727), .Z(n21729) );
  NAND U22727 ( .A(n21730), .B(n21729), .Z(n21766) );
  NANDN U22728 ( .A(n21732), .B(n21731), .Z(n21736) );
  OR U22729 ( .A(n21734), .B(n21733), .Z(n21735) );
  NAND U22730 ( .A(n21736), .B(n21735), .Z(n21763) );
  AND U22731 ( .A(b[2]), .B(a[915]), .Z(n21754) );
  AND U22732 ( .A(a[916]), .B(b[1]), .Z(n21752) );
  AND U22733 ( .A(a[914]), .B(b[3]), .Z(n21751) );
  XOR U22734 ( .A(n21752), .B(n21751), .Z(n21753) );
  XOR U22735 ( .A(n21754), .B(n21753), .Z(n21757) );
  NAND U22736 ( .A(b[0]), .B(a[917]), .Z(n21758) );
  XNOR U22737 ( .A(n21757), .B(n21758), .Z(n21759) );
  OR U22738 ( .A(n21738), .B(n21737), .Z(n21742) );
  NANDN U22739 ( .A(n21740), .B(n21739), .Z(n21741) );
  AND U22740 ( .A(n21742), .B(n21741), .Z(n21760) );
  XNOR U22741 ( .A(n21759), .B(n21760), .Z(n21764) );
  XNOR U22742 ( .A(n21763), .B(n21764), .Z(n21765) );
  XNOR U22743 ( .A(n21766), .B(n21765), .Z(n21750) );
  OR U22744 ( .A(n21743), .B(sreg[1936]), .Z(n21747) );
  NANDN U22745 ( .A(n21745), .B(n21744), .Z(n21746) );
  AND U22746 ( .A(n21747), .B(n21746), .Z(n21749) );
  XNOR U22747 ( .A(sreg[1937]), .B(n21749), .Z(n21748) );
  XNOR U22748 ( .A(n21750), .B(n21748), .Z(c[1937]) );
  AND U22749 ( .A(b[2]), .B(a[916]), .Z(n21778) );
  AND U22750 ( .A(a[917]), .B(b[1]), .Z(n21776) );
  AND U22751 ( .A(a[915]), .B(b[3]), .Z(n21775) );
  XOR U22752 ( .A(n21776), .B(n21775), .Z(n21777) );
  XOR U22753 ( .A(n21778), .B(n21777), .Z(n21781) );
  NAND U22754 ( .A(b[0]), .B(a[918]), .Z(n21782) );
  XOR U22755 ( .A(n21781), .B(n21782), .Z(n21784) );
  OR U22756 ( .A(n21752), .B(n21751), .Z(n21756) );
  NANDN U22757 ( .A(n21754), .B(n21753), .Z(n21755) );
  NAND U22758 ( .A(n21756), .B(n21755), .Z(n21783) );
  XNOR U22759 ( .A(n21784), .B(n21783), .Z(n21769) );
  NANDN U22760 ( .A(n21758), .B(n21757), .Z(n21762) );
  NAND U22761 ( .A(n21760), .B(n21759), .Z(n21761) );
  NAND U22762 ( .A(n21762), .B(n21761), .Z(n21770) );
  XNOR U22763 ( .A(n21769), .B(n21770), .Z(n21771) );
  NANDN U22764 ( .A(n21764), .B(n21763), .Z(n21768) );
  NANDN U22765 ( .A(n21766), .B(n21765), .Z(n21767) );
  NAND U22766 ( .A(n21768), .B(n21767), .Z(n21772) );
  XOR U22767 ( .A(n21771), .B(n21772), .Z(n21787) );
  XNOR U22768 ( .A(n21787), .B(sreg[1938]), .Z(n21788) );
  XOR U22769 ( .A(n21789), .B(n21788), .Z(c[1938]) );
  NANDN U22770 ( .A(n21770), .B(n21769), .Z(n21774) );
  NANDN U22771 ( .A(n21772), .B(n21771), .Z(n21773) );
  NAND U22772 ( .A(n21774), .B(n21773), .Z(n21810) );
  AND U22773 ( .A(b[2]), .B(a[917]), .Z(n21804) );
  AND U22774 ( .A(a[918]), .B(b[1]), .Z(n21802) );
  AND U22775 ( .A(a[916]), .B(b[3]), .Z(n21801) );
  XOR U22776 ( .A(n21802), .B(n21801), .Z(n21803) );
  XOR U22777 ( .A(n21804), .B(n21803), .Z(n21795) );
  NAND U22778 ( .A(b[0]), .B(a[919]), .Z(n21796) );
  XOR U22779 ( .A(n21795), .B(n21796), .Z(n21798) );
  OR U22780 ( .A(n21776), .B(n21775), .Z(n21780) );
  NANDN U22781 ( .A(n21778), .B(n21777), .Z(n21779) );
  NAND U22782 ( .A(n21780), .B(n21779), .Z(n21797) );
  XNOR U22783 ( .A(n21798), .B(n21797), .Z(n21807) );
  NANDN U22784 ( .A(n21782), .B(n21781), .Z(n21786) );
  OR U22785 ( .A(n21784), .B(n21783), .Z(n21785) );
  NAND U22786 ( .A(n21786), .B(n21785), .Z(n21808) );
  XNOR U22787 ( .A(n21807), .B(n21808), .Z(n21809) );
  XOR U22788 ( .A(n21810), .B(n21809), .Z(n21794) );
  NAND U22789 ( .A(n21787), .B(sreg[1938]), .Z(n21791) );
  OR U22790 ( .A(n21789), .B(n21788), .Z(n21790) );
  NAND U22791 ( .A(n21791), .B(n21790), .Z(n21793) );
  XNOR U22792 ( .A(sreg[1939]), .B(n21793), .Z(n21792) );
  XOR U22793 ( .A(n21794), .B(n21792), .Z(c[1939]) );
  NANDN U22794 ( .A(n21796), .B(n21795), .Z(n21800) );
  OR U22795 ( .A(n21798), .B(n21797), .Z(n21799) );
  NAND U22796 ( .A(n21800), .B(n21799), .Z(n21825) );
  AND U22797 ( .A(b[2]), .B(a[918]), .Z(n21816) );
  AND U22798 ( .A(a[919]), .B(b[1]), .Z(n21814) );
  AND U22799 ( .A(a[917]), .B(b[3]), .Z(n21813) );
  XOR U22800 ( .A(n21814), .B(n21813), .Z(n21815) );
  XOR U22801 ( .A(n21816), .B(n21815), .Z(n21819) );
  NAND U22802 ( .A(b[0]), .B(a[920]), .Z(n21820) );
  XNOR U22803 ( .A(n21819), .B(n21820), .Z(n21821) );
  OR U22804 ( .A(n21802), .B(n21801), .Z(n21806) );
  NANDN U22805 ( .A(n21804), .B(n21803), .Z(n21805) );
  AND U22806 ( .A(n21806), .B(n21805), .Z(n21822) );
  XNOR U22807 ( .A(n21821), .B(n21822), .Z(n21826) );
  XNOR U22808 ( .A(n21825), .B(n21826), .Z(n21827) );
  NANDN U22809 ( .A(n21808), .B(n21807), .Z(n21812) );
  NAND U22810 ( .A(n21810), .B(n21809), .Z(n21811) );
  NAND U22811 ( .A(n21812), .B(n21811), .Z(n21828) );
  XNOR U22812 ( .A(n21827), .B(n21828), .Z(n21831) );
  XOR U22813 ( .A(sreg[1940]), .B(n21831), .Z(n21833) );
  XNOR U22814 ( .A(n21832), .B(n21833), .Z(c[1940]) );
  AND U22815 ( .A(b[2]), .B(a[919]), .Z(n21848) );
  AND U22816 ( .A(a[920]), .B(b[1]), .Z(n21846) );
  AND U22817 ( .A(a[918]), .B(b[3]), .Z(n21845) );
  XOR U22818 ( .A(n21846), .B(n21845), .Z(n21847) );
  XOR U22819 ( .A(n21848), .B(n21847), .Z(n21851) );
  NAND U22820 ( .A(b[0]), .B(a[921]), .Z(n21852) );
  XOR U22821 ( .A(n21851), .B(n21852), .Z(n21854) );
  OR U22822 ( .A(n21814), .B(n21813), .Z(n21818) );
  NANDN U22823 ( .A(n21816), .B(n21815), .Z(n21817) );
  NAND U22824 ( .A(n21818), .B(n21817), .Z(n21853) );
  XNOR U22825 ( .A(n21854), .B(n21853), .Z(n21839) );
  NANDN U22826 ( .A(n21820), .B(n21819), .Z(n21824) );
  NAND U22827 ( .A(n21822), .B(n21821), .Z(n21823) );
  NAND U22828 ( .A(n21824), .B(n21823), .Z(n21840) );
  XNOR U22829 ( .A(n21839), .B(n21840), .Z(n21841) );
  NANDN U22830 ( .A(n21826), .B(n21825), .Z(n21830) );
  NANDN U22831 ( .A(n21828), .B(n21827), .Z(n21829) );
  NAND U22832 ( .A(n21830), .B(n21829), .Z(n21842) );
  XOR U22833 ( .A(n21841), .B(n21842), .Z(n21838) );
  OR U22834 ( .A(n21831), .B(sreg[1940]), .Z(n21835) );
  NAND U22835 ( .A(n21833), .B(n21832), .Z(n21834) );
  AND U22836 ( .A(n21835), .B(n21834), .Z(n21837) );
  XNOR U22837 ( .A(sreg[1941]), .B(n21837), .Z(n21836) );
  XNOR U22838 ( .A(n21838), .B(n21836), .Z(c[1941]) );
  NANDN U22839 ( .A(n21840), .B(n21839), .Z(n21844) );
  NANDN U22840 ( .A(n21842), .B(n21841), .Z(n21843) );
  NAND U22841 ( .A(n21844), .B(n21843), .Z(n21865) );
  AND U22842 ( .A(b[2]), .B(a[920]), .Z(n21871) );
  AND U22843 ( .A(a[921]), .B(b[1]), .Z(n21869) );
  AND U22844 ( .A(a[919]), .B(b[3]), .Z(n21868) );
  XOR U22845 ( .A(n21869), .B(n21868), .Z(n21870) );
  XOR U22846 ( .A(n21871), .B(n21870), .Z(n21874) );
  NAND U22847 ( .A(b[0]), .B(a[922]), .Z(n21875) );
  XOR U22848 ( .A(n21874), .B(n21875), .Z(n21877) );
  OR U22849 ( .A(n21846), .B(n21845), .Z(n21850) );
  NANDN U22850 ( .A(n21848), .B(n21847), .Z(n21849) );
  NAND U22851 ( .A(n21850), .B(n21849), .Z(n21876) );
  XNOR U22852 ( .A(n21877), .B(n21876), .Z(n21862) );
  NANDN U22853 ( .A(n21852), .B(n21851), .Z(n21856) );
  OR U22854 ( .A(n21854), .B(n21853), .Z(n21855) );
  NAND U22855 ( .A(n21856), .B(n21855), .Z(n21863) );
  XNOR U22856 ( .A(n21862), .B(n21863), .Z(n21864) );
  XNOR U22857 ( .A(n21865), .B(n21864), .Z(n21857) );
  XOR U22858 ( .A(sreg[1942]), .B(n21857), .Z(n21859) );
  XNOR U22859 ( .A(n21858), .B(n21859), .Z(c[1942]) );
  OR U22860 ( .A(n21857), .B(sreg[1942]), .Z(n21861) );
  NAND U22861 ( .A(n21859), .B(n21858), .Z(n21860) );
  AND U22862 ( .A(n21861), .B(n21860), .Z(n21881) );
  NANDN U22863 ( .A(n21863), .B(n21862), .Z(n21867) );
  NAND U22864 ( .A(n21865), .B(n21864), .Z(n21866) );
  NAND U22865 ( .A(n21867), .B(n21866), .Z(n21886) );
  AND U22866 ( .A(b[2]), .B(a[921]), .Z(n21892) );
  AND U22867 ( .A(a[922]), .B(b[1]), .Z(n21890) );
  AND U22868 ( .A(a[920]), .B(b[3]), .Z(n21889) );
  XOR U22869 ( .A(n21890), .B(n21889), .Z(n21891) );
  XOR U22870 ( .A(n21892), .B(n21891), .Z(n21895) );
  NAND U22871 ( .A(b[0]), .B(a[923]), .Z(n21896) );
  XOR U22872 ( .A(n21895), .B(n21896), .Z(n21898) );
  OR U22873 ( .A(n21869), .B(n21868), .Z(n21873) );
  NANDN U22874 ( .A(n21871), .B(n21870), .Z(n21872) );
  NAND U22875 ( .A(n21873), .B(n21872), .Z(n21897) );
  XNOR U22876 ( .A(n21898), .B(n21897), .Z(n21883) );
  NANDN U22877 ( .A(n21875), .B(n21874), .Z(n21879) );
  OR U22878 ( .A(n21877), .B(n21876), .Z(n21878) );
  NAND U22879 ( .A(n21879), .B(n21878), .Z(n21884) );
  XNOR U22880 ( .A(n21883), .B(n21884), .Z(n21885) );
  XNOR U22881 ( .A(n21886), .B(n21885), .Z(n21882) );
  XOR U22882 ( .A(sreg[1943]), .B(n21882), .Z(n21880) );
  XOR U22883 ( .A(n21881), .B(n21880), .Z(c[1943]) );
  NANDN U22884 ( .A(n21884), .B(n21883), .Z(n21888) );
  NAND U22885 ( .A(n21886), .B(n21885), .Z(n21887) );
  NAND U22886 ( .A(n21888), .B(n21887), .Z(n21909) );
  AND U22887 ( .A(b[2]), .B(a[922]), .Z(n21915) );
  AND U22888 ( .A(a[923]), .B(b[1]), .Z(n21913) );
  AND U22889 ( .A(a[921]), .B(b[3]), .Z(n21912) );
  XOR U22890 ( .A(n21913), .B(n21912), .Z(n21914) );
  XOR U22891 ( .A(n21915), .B(n21914), .Z(n21918) );
  NAND U22892 ( .A(b[0]), .B(a[924]), .Z(n21919) );
  XOR U22893 ( .A(n21918), .B(n21919), .Z(n21921) );
  OR U22894 ( .A(n21890), .B(n21889), .Z(n21894) );
  NANDN U22895 ( .A(n21892), .B(n21891), .Z(n21893) );
  NAND U22896 ( .A(n21894), .B(n21893), .Z(n21920) );
  XNOR U22897 ( .A(n21921), .B(n21920), .Z(n21906) );
  NANDN U22898 ( .A(n21896), .B(n21895), .Z(n21900) );
  OR U22899 ( .A(n21898), .B(n21897), .Z(n21899) );
  NAND U22900 ( .A(n21900), .B(n21899), .Z(n21907) );
  XNOR U22901 ( .A(n21906), .B(n21907), .Z(n21908) );
  XNOR U22902 ( .A(n21909), .B(n21908), .Z(n21901) );
  XOR U22903 ( .A(sreg[1944]), .B(n21901), .Z(n21902) );
  XOR U22904 ( .A(n21903), .B(n21902), .Z(c[1944]) );
  OR U22905 ( .A(n21901), .B(sreg[1944]), .Z(n21905) );
  NANDN U22906 ( .A(n21903), .B(n21902), .Z(n21904) );
  NAND U22907 ( .A(n21905), .B(n21904), .Z(n21926) );
  NANDN U22908 ( .A(n21907), .B(n21906), .Z(n21911) );
  NAND U22909 ( .A(n21909), .B(n21908), .Z(n21910) );
  NAND U22910 ( .A(n21911), .B(n21910), .Z(n21932) );
  AND U22911 ( .A(b[2]), .B(a[923]), .Z(n21938) );
  AND U22912 ( .A(a[924]), .B(b[1]), .Z(n21936) );
  AND U22913 ( .A(a[922]), .B(b[3]), .Z(n21935) );
  XOR U22914 ( .A(n21936), .B(n21935), .Z(n21937) );
  XOR U22915 ( .A(n21938), .B(n21937), .Z(n21941) );
  NAND U22916 ( .A(b[0]), .B(a[925]), .Z(n21942) );
  XOR U22917 ( .A(n21941), .B(n21942), .Z(n21944) );
  OR U22918 ( .A(n21913), .B(n21912), .Z(n21917) );
  NANDN U22919 ( .A(n21915), .B(n21914), .Z(n21916) );
  NAND U22920 ( .A(n21917), .B(n21916), .Z(n21943) );
  XNOR U22921 ( .A(n21944), .B(n21943), .Z(n21929) );
  NANDN U22922 ( .A(n21919), .B(n21918), .Z(n21923) );
  OR U22923 ( .A(n21921), .B(n21920), .Z(n21922) );
  NAND U22924 ( .A(n21923), .B(n21922), .Z(n21930) );
  XNOR U22925 ( .A(n21929), .B(n21930), .Z(n21931) );
  XNOR U22926 ( .A(n21932), .B(n21931), .Z(n21924) );
  XNOR U22927 ( .A(n21924), .B(sreg[1945]), .Z(n21925) );
  XOR U22928 ( .A(n21926), .B(n21925), .Z(c[1945]) );
  NAND U22929 ( .A(n21924), .B(sreg[1945]), .Z(n21928) );
  OR U22930 ( .A(n21926), .B(n21925), .Z(n21927) );
  AND U22931 ( .A(n21928), .B(n21927), .Z(n21967) );
  NANDN U22932 ( .A(n21930), .B(n21929), .Z(n21934) );
  NAND U22933 ( .A(n21932), .B(n21931), .Z(n21933) );
  NAND U22934 ( .A(n21934), .B(n21933), .Z(n21951) );
  AND U22935 ( .A(b[2]), .B(a[924]), .Z(n21957) );
  AND U22936 ( .A(a[925]), .B(b[1]), .Z(n21955) );
  AND U22937 ( .A(a[923]), .B(b[3]), .Z(n21954) );
  XOR U22938 ( .A(n21955), .B(n21954), .Z(n21956) );
  XOR U22939 ( .A(n21957), .B(n21956), .Z(n21960) );
  NAND U22940 ( .A(b[0]), .B(a[926]), .Z(n21961) );
  XOR U22941 ( .A(n21960), .B(n21961), .Z(n21963) );
  OR U22942 ( .A(n21936), .B(n21935), .Z(n21940) );
  NANDN U22943 ( .A(n21938), .B(n21937), .Z(n21939) );
  NAND U22944 ( .A(n21940), .B(n21939), .Z(n21962) );
  XNOR U22945 ( .A(n21963), .B(n21962), .Z(n21948) );
  NANDN U22946 ( .A(n21942), .B(n21941), .Z(n21946) );
  OR U22947 ( .A(n21944), .B(n21943), .Z(n21945) );
  NAND U22948 ( .A(n21946), .B(n21945), .Z(n21949) );
  XNOR U22949 ( .A(n21948), .B(n21949), .Z(n21950) );
  XNOR U22950 ( .A(n21951), .B(n21950), .Z(n21966) );
  XNOR U22951 ( .A(sreg[1946]), .B(n21966), .Z(n21947) );
  XOR U22952 ( .A(n21967), .B(n21947), .Z(c[1946]) );
  NANDN U22953 ( .A(n21949), .B(n21948), .Z(n21953) );
  NAND U22954 ( .A(n21951), .B(n21950), .Z(n21952) );
  NAND U22955 ( .A(n21953), .B(n21952), .Z(n21974) );
  AND U22956 ( .A(b[2]), .B(a[925]), .Z(n21980) );
  AND U22957 ( .A(a[926]), .B(b[1]), .Z(n21978) );
  AND U22958 ( .A(a[924]), .B(b[3]), .Z(n21977) );
  XOR U22959 ( .A(n21978), .B(n21977), .Z(n21979) );
  XOR U22960 ( .A(n21980), .B(n21979), .Z(n21983) );
  NAND U22961 ( .A(b[0]), .B(a[927]), .Z(n21984) );
  XOR U22962 ( .A(n21983), .B(n21984), .Z(n21986) );
  OR U22963 ( .A(n21955), .B(n21954), .Z(n21959) );
  NANDN U22964 ( .A(n21957), .B(n21956), .Z(n21958) );
  NAND U22965 ( .A(n21959), .B(n21958), .Z(n21985) );
  XNOR U22966 ( .A(n21986), .B(n21985), .Z(n21971) );
  NANDN U22967 ( .A(n21961), .B(n21960), .Z(n21965) );
  OR U22968 ( .A(n21963), .B(n21962), .Z(n21964) );
  NAND U22969 ( .A(n21965), .B(n21964), .Z(n21972) );
  XNOR U22970 ( .A(n21971), .B(n21972), .Z(n21973) );
  XNOR U22971 ( .A(n21974), .B(n21973), .Z(n21970) );
  XOR U22972 ( .A(n21969), .B(sreg[1947]), .Z(n21968) );
  XOR U22973 ( .A(n21970), .B(n21968), .Z(c[1947]) );
  NANDN U22974 ( .A(n21972), .B(n21971), .Z(n21976) );
  NAND U22975 ( .A(n21974), .B(n21973), .Z(n21975) );
  NAND U22976 ( .A(n21976), .B(n21975), .Z(n21992) );
  AND U22977 ( .A(b[2]), .B(a[926]), .Z(n21998) );
  AND U22978 ( .A(a[927]), .B(b[1]), .Z(n21996) );
  AND U22979 ( .A(a[925]), .B(b[3]), .Z(n21995) );
  XOR U22980 ( .A(n21996), .B(n21995), .Z(n21997) );
  XOR U22981 ( .A(n21998), .B(n21997), .Z(n22001) );
  NAND U22982 ( .A(b[0]), .B(a[928]), .Z(n22002) );
  XOR U22983 ( .A(n22001), .B(n22002), .Z(n22004) );
  OR U22984 ( .A(n21978), .B(n21977), .Z(n21982) );
  NANDN U22985 ( .A(n21980), .B(n21979), .Z(n21981) );
  NAND U22986 ( .A(n21982), .B(n21981), .Z(n22003) );
  XNOR U22987 ( .A(n22004), .B(n22003), .Z(n21989) );
  NANDN U22988 ( .A(n21984), .B(n21983), .Z(n21988) );
  OR U22989 ( .A(n21986), .B(n21985), .Z(n21987) );
  NAND U22990 ( .A(n21988), .B(n21987), .Z(n21990) );
  XNOR U22991 ( .A(n21989), .B(n21990), .Z(n21991) );
  XNOR U22992 ( .A(n21992), .B(n21991), .Z(n22007) );
  XNOR U22993 ( .A(n22007), .B(sreg[1948]), .Z(n22009) );
  XNOR U22994 ( .A(n22008), .B(n22009), .Z(c[1948]) );
  NANDN U22995 ( .A(n21990), .B(n21989), .Z(n21994) );
  NAND U22996 ( .A(n21992), .B(n21991), .Z(n21993) );
  NAND U22997 ( .A(n21994), .B(n21993), .Z(n22016) );
  AND U22998 ( .A(b[2]), .B(a[927]), .Z(n22028) );
  AND U22999 ( .A(a[928]), .B(b[1]), .Z(n22026) );
  AND U23000 ( .A(a[926]), .B(b[3]), .Z(n22025) );
  XOR U23001 ( .A(n22026), .B(n22025), .Z(n22027) );
  XOR U23002 ( .A(n22028), .B(n22027), .Z(n22019) );
  NAND U23003 ( .A(b[0]), .B(a[929]), .Z(n22020) );
  XOR U23004 ( .A(n22019), .B(n22020), .Z(n22022) );
  OR U23005 ( .A(n21996), .B(n21995), .Z(n22000) );
  NANDN U23006 ( .A(n21998), .B(n21997), .Z(n21999) );
  NAND U23007 ( .A(n22000), .B(n21999), .Z(n22021) );
  XNOR U23008 ( .A(n22022), .B(n22021), .Z(n22013) );
  NANDN U23009 ( .A(n22002), .B(n22001), .Z(n22006) );
  OR U23010 ( .A(n22004), .B(n22003), .Z(n22005) );
  NAND U23011 ( .A(n22006), .B(n22005), .Z(n22014) );
  XNOR U23012 ( .A(n22013), .B(n22014), .Z(n22015) );
  XNOR U23013 ( .A(n22016), .B(n22015), .Z(n22033) );
  NAND U23014 ( .A(n22007), .B(sreg[1948]), .Z(n22011) );
  NANDN U23015 ( .A(n22009), .B(n22008), .Z(n22010) );
  AND U23016 ( .A(n22011), .B(n22010), .Z(n22032) );
  XNOR U23017 ( .A(n22032), .B(sreg[1949]), .Z(n22012) );
  XOR U23018 ( .A(n22033), .B(n22012), .Z(c[1949]) );
  NANDN U23019 ( .A(n22014), .B(n22013), .Z(n22018) );
  NAND U23020 ( .A(n22016), .B(n22015), .Z(n22017) );
  NAND U23021 ( .A(n22018), .B(n22017), .Z(n22039) );
  NANDN U23022 ( .A(n22020), .B(n22019), .Z(n22024) );
  OR U23023 ( .A(n22022), .B(n22021), .Z(n22023) );
  AND U23024 ( .A(n22024), .B(n22023), .Z(n22038) );
  AND U23025 ( .A(b[2]), .B(a[928]), .Z(n22043) );
  AND U23026 ( .A(a[929]), .B(b[1]), .Z(n22041) );
  AND U23027 ( .A(a[927]), .B(b[3]), .Z(n22040) );
  XOR U23028 ( .A(n22041), .B(n22040), .Z(n22042) );
  XOR U23029 ( .A(n22043), .B(n22042), .Z(n22046) );
  NAND U23030 ( .A(b[0]), .B(a[930]), .Z(n22047) );
  XOR U23031 ( .A(n22046), .B(n22047), .Z(n22049) );
  OR U23032 ( .A(n22026), .B(n22025), .Z(n22030) );
  NANDN U23033 ( .A(n22028), .B(n22027), .Z(n22029) );
  NAND U23034 ( .A(n22030), .B(n22029), .Z(n22048) );
  XOR U23035 ( .A(n22049), .B(n22048), .Z(n22037) );
  XNOR U23036 ( .A(n22038), .B(n22037), .Z(n22031) );
  XNOR U23037 ( .A(n22039), .B(n22031), .Z(n22036) );
  XOR U23038 ( .A(n22035), .B(sreg[1950]), .Z(n22034) );
  XOR U23039 ( .A(n22036), .B(n22034), .Z(c[1950]) );
  AND U23040 ( .A(b[2]), .B(a[929]), .Z(n22061) );
  AND U23041 ( .A(a[930]), .B(b[1]), .Z(n22059) );
  AND U23042 ( .A(a[928]), .B(b[3]), .Z(n22058) );
  XOR U23043 ( .A(n22059), .B(n22058), .Z(n22060) );
  XOR U23044 ( .A(n22061), .B(n22060), .Z(n22064) );
  NAND U23045 ( .A(b[0]), .B(a[931]), .Z(n22065) );
  XOR U23046 ( .A(n22064), .B(n22065), .Z(n22067) );
  OR U23047 ( .A(n22041), .B(n22040), .Z(n22045) );
  NANDN U23048 ( .A(n22043), .B(n22042), .Z(n22044) );
  NAND U23049 ( .A(n22045), .B(n22044), .Z(n22066) );
  XNOR U23050 ( .A(n22067), .B(n22066), .Z(n22052) );
  NANDN U23051 ( .A(n22047), .B(n22046), .Z(n22051) );
  OR U23052 ( .A(n22049), .B(n22048), .Z(n22050) );
  NAND U23053 ( .A(n22051), .B(n22050), .Z(n22053) );
  XNOR U23054 ( .A(n22052), .B(n22053), .Z(n22054) );
  XOR U23055 ( .A(n22055), .B(n22054), .Z(n22070) );
  XNOR U23056 ( .A(n22070), .B(sreg[1951]), .Z(n22072) );
  XNOR U23057 ( .A(n22071), .B(n22072), .Z(c[1951]) );
  NANDN U23058 ( .A(n22053), .B(n22052), .Z(n22057) );
  NANDN U23059 ( .A(n22055), .B(n22054), .Z(n22056) );
  NAND U23060 ( .A(n22057), .B(n22056), .Z(n22078) );
  AND U23061 ( .A(b[2]), .B(a[930]), .Z(n22084) );
  AND U23062 ( .A(a[931]), .B(b[1]), .Z(n22082) );
  AND U23063 ( .A(a[929]), .B(b[3]), .Z(n22081) );
  XOR U23064 ( .A(n22082), .B(n22081), .Z(n22083) );
  XOR U23065 ( .A(n22084), .B(n22083), .Z(n22087) );
  NAND U23066 ( .A(b[0]), .B(a[932]), .Z(n22088) );
  XOR U23067 ( .A(n22087), .B(n22088), .Z(n22090) );
  OR U23068 ( .A(n22059), .B(n22058), .Z(n22063) );
  NANDN U23069 ( .A(n22061), .B(n22060), .Z(n22062) );
  NAND U23070 ( .A(n22063), .B(n22062), .Z(n22089) );
  XNOR U23071 ( .A(n22090), .B(n22089), .Z(n22075) );
  NANDN U23072 ( .A(n22065), .B(n22064), .Z(n22069) );
  OR U23073 ( .A(n22067), .B(n22066), .Z(n22068) );
  NAND U23074 ( .A(n22069), .B(n22068), .Z(n22076) );
  XNOR U23075 ( .A(n22075), .B(n22076), .Z(n22077) );
  XNOR U23076 ( .A(n22078), .B(n22077), .Z(n22094) );
  XNOR U23077 ( .A(n22094), .B(sreg[1952]), .Z(n22096) );
  NAND U23078 ( .A(n22070), .B(sreg[1951]), .Z(n22074) );
  NANDN U23079 ( .A(n22072), .B(n22071), .Z(n22073) );
  AND U23080 ( .A(n22074), .B(n22073), .Z(n22095) );
  XOR U23081 ( .A(n22096), .B(n22095), .Z(c[1952]) );
  NANDN U23082 ( .A(n22076), .B(n22075), .Z(n22080) );
  NAND U23083 ( .A(n22078), .B(n22077), .Z(n22079) );
  NAND U23084 ( .A(n22080), .B(n22079), .Z(n22104) );
  AND U23085 ( .A(b[2]), .B(a[931]), .Z(n22108) );
  AND U23086 ( .A(a[932]), .B(b[1]), .Z(n22106) );
  AND U23087 ( .A(a[930]), .B(b[3]), .Z(n22105) );
  XOR U23088 ( .A(n22106), .B(n22105), .Z(n22107) );
  XOR U23089 ( .A(n22108), .B(n22107), .Z(n22111) );
  NAND U23090 ( .A(b[0]), .B(a[933]), .Z(n22112) );
  XOR U23091 ( .A(n22111), .B(n22112), .Z(n22113) );
  OR U23092 ( .A(n22082), .B(n22081), .Z(n22086) );
  NANDN U23093 ( .A(n22084), .B(n22083), .Z(n22085) );
  AND U23094 ( .A(n22086), .B(n22085), .Z(n22114) );
  XOR U23095 ( .A(n22113), .B(n22114), .Z(n22102) );
  NANDN U23096 ( .A(n22088), .B(n22087), .Z(n22092) );
  OR U23097 ( .A(n22090), .B(n22089), .Z(n22091) );
  AND U23098 ( .A(n22092), .B(n22091), .Z(n22103) );
  XOR U23099 ( .A(n22102), .B(n22103), .Z(n22093) );
  XOR U23100 ( .A(n22104), .B(n22093), .Z(n22101) );
  NAND U23101 ( .A(n22094), .B(sreg[1952]), .Z(n22098) );
  OR U23102 ( .A(n22096), .B(n22095), .Z(n22097) );
  AND U23103 ( .A(n22098), .B(n22097), .Z(n22100) );
  XNOR U23104 ( .A(n22100), .B(sreg[1953]), .Z(n22099) );
  XNOR U23105 ( .A(n22101), .B(n22099), .Z(c[1953]) );
  AND U23106 ( .A(b[2]), .B(a[932]), .Z(n22124) );
  AND U23107 ( .A(a[933]), .B(b[1]), .Z(n22122) );
  AND U23108 ( .A(a[931]), .B(b[3]), .Z(n22121) );
  XOR U23109 ( .A(n22122), .B(n22121), .Z(n22123) );
  XOR U23110 ( .A(n22124), .B(n22123), .Z(n22127) );
  NAND U23111 ( .A(b[0]), .B(a[934]), .Z(n22128) );
  XOR U23112 ( .A(n22127), .B(n22128), .Z(n22130) );
  OR U23113 ( .A(n22106), .B(n22105), .Z(n22110) );
  NANDN U23114 ( .A(n22108), .B(n22107), .Z(n22109) );
  NAND U23115 ( .A(n22110), .B(n22109), .Z(n22129) );
  XNOR U23116 ( .A(n22130), .B(n22129), .Z(n22115) );
  XNOR U23117 ( .A(n22115), .B(n22116), .Z(n22118) );
  XOR U23118 ( .A(n22117), .B(n22118), .Z(n22133) );
  XOR U23119 ( .A(n22133), .B(sreg[1954]), .Z(n22135) );
  XNOR U23120 ( .A(n22134), .B(n22135), .Z(c[1954]) );
  NANDN U23121 ( .A(n22116), .B(n22115), .Z(n22120) );
  NAND U23122 ( .A(n22118), .B(n22117), .Z(n22119) );
  NAND U23123 ( .A(n22120), .B(n22119), .Z(n22153) );
  AND U23124 ( .A(b[2]), .B(a[933]), .Z(n22147) );
  AND U23125 ( .A(a[934]), .B(b[1]), .Z(n22145) );
  AND U23126 ( .A(a[932]), .B(b[3]), .Z(n22144) );
  XOR U23127 ( .A(n22145), .B(n22144), .Z(n22146) );
  XOR U23128 ( .A(n22147), .B(n22146), .Z(n22138) );
  NAND U23129 ( .A(b[0]), .B(a[935]), .Z(n22139) );
  XOR U23130 ( .A(n22138), .B(n22139), .Z(n22141) );
  OR U23131 ( .A(n22122), .B(n22121), .Z(n22126) );
  NANDN U23132 ( .A(n22124), .B(n22123), .Z(n22125) );
  NAND U23133 ( .A(n22126), .B(n22125), .Z(n22140) );
  XNOR U23134 ( .A(n22141), .B(n22140), .Z(n22150) );
  NANDN U23135 ( .A(n22128), .B(n22127), .Z(n22132) );
  OR U23136 ( .A(n22130), .B(n22129), .Z(n22131) );
  NAND U23137 ( .A(n22132), .B(n22131), .Z(n22151) );
  XNOR U23138 ( .A(n22150), .B(n22151), .Z(n22152) );
  XNOR U23139 ( .A(n22153), .B(n22152), .Z(n22156) );
  XOR U23140 ( .A(sreg[1955]), .B(n22156), .Z(n22157) );
  NANDN U23141 ( .A(n22133), .B(sreg[1954]), .Z(n22137) );
  NANDN U23142 ( .A(n22135), .B(n22134), .Z(n22136) );
  NAND U23143 ( .A(n22137), .B(n22136), .Z(n22158) );
  XOR U23144 ( .A(n22157), .B(n22158), .Z(c[1955]) );
  NANDN U23145 ( .A(n22139), .B(n22138), .Z(n22143) );
  OR U23146 ( .A(n22141), .B(n22140), .Z(n22142) );
  NAND U23147 ( .A(n22143), .B(n22142), .Z(n22162) );
  AND U23148 ( .A(b[2]), .B(a[934]), .Z(n22171) );
  AND U23149 ( .A(a[935]), .B(b[1]), .Z(n22169) );
  AND U23150 ( .A(a[933]), .B(b[3]), .Z(n22168) );
  XOR U23151 ( .A(n22169), .B(n22168), .Z(n22170) );
  XOR U23152 ( .A(n22171), .B(n22170), .Z(n22174) );
  NAND U23153 ( .A(b[0]), .B(a[936]), .Z(n22175) );
  XNOR U23154 ( .A(n22174), .B(n22175), .Z(n22176) );
  OR U23155 ( .A(n22145), .B(n22144), .Z(n22149) );
  NANDN U23156 ( .A(n22147), .B(n22146), .Z(n22148) );
  AND U23157 ( .A(n22149), .B(n22148), .Z(n22177) );
  XNOR U23158 ( .A(n22176), .B(n22177), .Z(n22163) );
  XNOR U23159 ( .A(n22162), .B(n22163), .Z(n22164) );
  NANDN U23160 ( .A(n22151), .B(n22150), .Z(n22155) );
  NAND U23161 ( .A(n22153), .B(n22152), .Z(n22154) );
  AND U23162 ( .A(n22155), .B(n22154), .Z(n22165) );
  XNOR U23163 ( .A(n22164), .B(n22165), .Z(n22181) );
  OR U23164 ( .A(n22156), .B(sreg[1955]), .Z(n22160) );
  NANDN U23165 ( .A(n22158), .B(n22157), .Z(n22159) );
  AND U23166 ( .A(n22160), .B(n22159), .Z(n22180) );
  XNOR U23167 ( .A(n22180), .B(sreg[1956]), .Z(n22161) );
  XOR U23168 ( .A(n22181), .B(n22161), .Z(c[1956]) );
  NANDN U23169 ( .A(n22163), .B(n22162), .Z(n22167) );
  NAND U23170 ( .A(n22165), .B(n22164), .Z(n22166) );
  NAND U23171 ( .A(n22167), .B(n22166), .Z(n22185) );
  AND U23172 ( .A(b[2]), .B(a[935]), .Z(n22191) );
  AND U23173 ( .A(a[936]), .B(b[1]), .Z(n22189) );
  AND U23174 ( .A(a[934]), .B(b[3]), .Z(n22188) );
  XOR U23175 ( .A(n22189), .B(n22188), .Z(n22190) );
  XOR U23176 ( .A(n22191), .B(n22190), .Z(n22194) );
  NAND U23177 ( .A(b[0]), .B(a[937]), .Z(n22195) );
  XOR U23178 ( .A(n22194), .B(n22195), .Z(n22197) );
  OR U23179 ( .A(n22169), .B(n22168), .Z(n22173) );
  NANDN U23180 ( .A(n22171), .B(n22170), .Z(n22172) );
  NAND U23181 ( .A(n22173), .B(n22172), .Z(n22196) );
  XNOR U23182 ( .A(n22197), .B(n22196), .Z(n22182) );
  NANDN U23183 ( .A(n22175), .B(n22174), .Z(n22179) );
  NAND U23184 ( .A(n22177), .B(n22176), .Z(n22178) );
  NAND U23185 ( .A(n22179), .B(n22178), .Z(n22183) );
  XNOR U23186 ( .A(n22182), .B(n22183), .Z(n22184) );
  XOR U23187 ( .A(n22185), .B(n22184), .Z(n22200) );
  XNOR U23188 ( .A(n22200), .B(sreg[1957]), .Z(n22202) );
  XOR U23189 ( .A(n22202), .B(n22201), .Z(c[1957]) );
  NANDN U23190 ( .A(n22183), .B(n22182), .Z(n22187) );
  NANDN U23191 ( .A(n22185), .B(n22184), .Z(n22186) );
  NAND U23192 ( .A(n22187), .B(n22186), .Z(n22208) );
  AND U23193 ( .A(b[2]), .B(a[936]), .Z(n22214) );
  AND U23194 ( .A(a[937]), .B(b[1]), .Z(n22212) );
  AND U23195 ( .A(a[935]), .B(b[3]), .Z(n22211) );
  XOR U23196 ( .A(n22212), .B(n22211), .Z(n22213) );
  XOR U23197 ( .A(n22214), .B(n22213), .Z(n22217) );
  NAND U23198 ( .A(b[0]), .B(a[938]), .Z(n22218) );
  XOR U23199 ( .A(n22217), .B(n22218), .Z(n22220) );
  OR U23200 ( .A(n22189), .B(n22188), .Z(n22193) );
  NANDN U23201 ( .A(n22191), .B(n22190), .Z(n22192) );
  NAND U23202 ( .A(n22193), .B(n22192), .Z(n22219) );
  XNOR U23203 ( .A(n22220), .B(n22219), .Z(n22205) );
  NANDN U23204 ( .A(n22195), .B(n22194), .Z(n22199) );
  OR U23205 ( .A(n22197), .B(n22196), .Z(n22198) );
  NAND U23206 ( .A(n22199), .B(n22198), .Z(n22206) );
  XNOR U23207 ( .A(n22205), .B(n22206), .Z(n22207) );
  XNOR U23208 ( .A(n22208), .B(n22207), .Z(n22223) );
  XNOR U23209 ( .A(n22223), .B(sreg[1958]), .Z(n22225) );
  NAND U23210 ( .A(n22200), .B(sreg[1957]), .Z(n22204) );
  OR U23211 ( .A(n22202), .B(n22201), .Z(n22203) );
  AND U23212 ( .A(n22204), .B(n22203), .Z(n22224) );
  XOR U23213 ( .A(n22225), .B(n22224), .Z(c[1958]) );
  NANDN U23214 ( .A(n22206), .B(n22205), .Z(n22210) );
  NAND U23215 ( .A(n22208), .B(n22207), .Z(n22209) );
  NAND U23216 ( .A(n22210), .B(n22209), .Z(n22231) );
  AND U23217 ( .A(b[2]), .B(a[937]), .Z(n22237) );
  AND U23218 ( .A(a[938]), .B(b[1]), .Z(n22235) );
  AND U23219 ( .A(a[936]), .B(b[3]), .Z(n22234) );
  XOR U23220 ( .A(n22235), .B(n22234), .Z(n22236) );
  XOR U23221 ( .A(n22237), .B(n22236), .Z(n22240) );
  NAND U23222 ( .A(b[0]), .B(a[939]), .Z(n22241) );
  XOR U23223 ( .A(n22240), .B(n22241), .Z(n22243) );
  OR U23224 ( .A(n22212), .B(n22211), .Z(n22216) );
  NANDN U23225 ( .A(n22214), .B(n22213), .Z(n22215) );
  NAND U23226 ( .A(n22216), .B(n22215), .Z(n22242) );
  XNOR U23227 ( .A(n22243), .B(n22242), .Z(n22228) );
  NANDN U23228 ( .A(n22218), .B(n22217), .Z(n22222) );
  OR U23229 ( .A(n22220), .B(n22219), .Z(n22221) );
  NAND U23230 ( .A(n22222), .B(n22221), .Z(n22229) );
  XNOR U23231 ( .A(n22228), .B(n22229), .Z(n22230) );
  XNOR U23232 ( .A(n22231), .B(n22230), .Z(n22246) );
  XNOR U23233 ( .A(n22246), .B(sreg[1959]), .Z(n22248) );
  NAND U23234 ( .A(n22223), .B(sreg[1958]), .Z(n22227) );
  OR U23235 ( .A(n22225), .B(n22224), .Z(n22226) );
  AND U23236 ( .A(n22227), .B(n22226), .Z(n22247) );
  XOR U23237 ( .A(n22248), .B(n22247), .Z(c[1959]) );
  NANDN U23238 ( .A(n22229), .B(n22228), .Z(n22233) );
  NAND U23239 ( .A(n22231), .B(n22230), .Z(n22232) );
  NAND U23240 ( .A(n22233), .B(n22232), .Z(n22255) );
  AND U23241 ( .A(b[2]), .B(a[938]), .Z(n22261) );
  AND U23242 ( .A(a[939]), .B(b[1]), .Z(n22259) );
  AND U23243 ( .A(a[937]), .B(b[3]), .Z(n22258) );
  XOR U23244 ( .A(n22259), .B(n22258), .Z(n22260) );
  XOR U23245 ( .A(n22261), .B(n22260), .Z(n22264) );
  NAND U23246 ( .A(b[0]), .B(a[940]), .Z(n22265) );
  XOR U23247 ( .A(n22264), .B(n22265), .Z(n22267) );
  OR U23248 ( .A(n22235), .B(n22234), .Z(n22239) );
  NANDN U23249 ( .A(n22237), .B(n22236), .Z(n22238) );
  NAND U23250 ( .A(n22239), .B(n22238), .Z(n22266) );
  XNOR U23251 ( .A(n22267), .B(n22266), .Z(n22252) );
  NANDN U23252 ( .A(n22241), .B(n22240), .Z(n22245) );
  OR U23253 ( .A(n22243), .B(n22242), .Z(n22244) );
  NAND U23254 ( .A(n22245), .B(n22244), .Z(n22253) );
  XNOR U23255 ( .A(n22252), .B(n22253), .Z(n22254) );
  XOR U23256 ( .A(n22255), .B(n22254), .Z(n22271) );
  NAND U23257 ( .A(n22246), .B(sreg[1959]), .Z(n22250) );
  OR U23258 ( .A(n22248), .B(n22247), .Z(n22249) );
  NAND U23259 ( .A(n22250), .B(n22249), .Z(n22270) );
  XNOR U23260 ( .A(sreg[1960]), .B(n22270), .Z(n22251) );
  XOR U23261 ( .A(n22271), .B(n22251), .Z(c[1960]) );
  NANDN U23262 ( .A(n22253), .B(n22252), .Z(n22257) );
  NAND U23263 ( .A(n22255), .B(n22254), .Z(n22256) );
  NAND U23264 ( .A(n22257), .B(n22256), .Z(n22276) );
  AND U23265 ( .A(b[2]), .B(a[939]), .Z(n22282) );
  AND U23266 ( .A(a[940]), .B(b[1]), .Z(n22280) );
  AND U23267 ( .A(a[938]), .B(b[3]), .Z(n22279) );
  XOR U23268 ( .A(n22280), .B(n22279), .Z(n22281) );
  XOR U23269 ( .A(n22282), .B(n22281), .Z(n22285) );
  NAND U23270 ( .A(b[0]), .B(a[941]), .Z(n22286) );
  XOR U23271 ( .A(n22285), .B(n22286), .Z(n22288) );
  OR U23272 ( .A(n22259), .B(n22258), .Z(n22263) );
  NANDN U23273 ( .A(n22261), .B(n22260), .Z(n22262) );
  NAND U23274 ( .A(n22263), .B(n22262), .Z(n22287) );
  XNOR U23275 ( .A(n22288), .B(n22287), .Z(n22273) );
  NANDN U23276 ( .A(n22265), .B(n22264), .Z(n22269) );
  OR U23277 ( .A(n22267), .B(n22266), .Z(n22268) );
  NAND U23278 ( .A(n22269), .B(n22268), .Z(n22274) );
  XNOR U23279 ( .A(n22273), .B(n22274), .Z(n22275) );
  XOR U23280 ( .A(n22276), .B(n22275), .Z(n22292) );
  XNOR U23281 ( .A(sreg[1961]), .B(n22291), .Z(n22272) );
  XOR U23282 ( .A(n22292), .B(n22272), .Z(c[1961]) );
  NANDN U23283 ( .A(n22274), .B(n22273), .Z(n22278) );
  NAND U23284 ( .A(n22276), .B(n22275), .Z(n22277) );
  NAND U23285 ( .A(n22278), .B(n22277), .Z(n22299) );
  AND U23286 ( .A(b[2]), .B(a[940]), .Z(n22305) );
  AND U23287 ( .A(a[941]), .B(b[1]), .Z(n22303) );
  AND U23288 ( .A(a[939]), .B(b[3]), .Z(n22302) );
  XOR U23289 ( .A(n22303), .B(n22302), .Z(n22304) );
  XOR U23290 ( .A(n22305), .B(n22304), .Z(n22308) );
  NAND U23291 ( .A(b[0]), .B(a[942]), .Z(n22309) );
  XOR U23292 ( .A(n22308), .B(n22309), .Z(n22311) );
  OR U23293 ( .A(n22280), .B(n22279), .Z(n22284) );
  NANDN U23294 ( .A(n22282), .B(n22281), .Z(n22283) );
  NAND U23295 ( .A(n22284), .B(n22283), .Z(n22310) );
  XNOR U23296 ( .A(n22311), .B(n22310), .Z(n22296) );
  NANDN U23297 ( .A(n22286), .B(n22285), .Z(n22290) );
  OR U23298 ( .A(n22288), .B(n22287), .Z(n22289) );
  NAND U23299 ( .A(n22290), .B(n22289), .Z(n22297) );
  XNOR U23300 ( .A(n22296), .B(n22297), .Z(n22298) );
  XOR U23301 ( .A(n22299), .B(n22298), .Z(n22295) );
  XNOR U23302 ( .A(sreg[1962]), .B(n22294), .Z(n22293) );
  XOR U23303 ( .A(n22295), .B(n22293), .Z(c[1962]) );
  NANDN U23304 ( .A(n22297), .B(n22296), .Z(n22301) );
  NAND U23305 ( .A(n22299), .B(n22298), .Z(n22300) );
  NAND U23306 ( .A(n22301), .B(n22300), .Z(n22322) );
  AND U23307 ( .A(b[2]), .B(a[941]), .Z(n22328) );
  AND U23308 ( .A(a[942]), .B(b[1]), .Z(n22326) );
  AND U23309 ( .A(a[940]), .B(b[3]), .Z(n22325) );
  XOR U23310 ( .A(n22326), .B(n22325), .Z(n22327) );
  XOR U23311 ( .A(n22328), .B(n22327), .Z(n22331) );
  NAND U23312 ( .A(b[0]), .B(a[943]), .Z(n22332) );
  XOR U23313 ( .A(n22331), .B(n22332), .Z(n22334) );
  OR U23314 ( .A(n22303), .B(n22302), .Z(n22307) );
  NANDN U23315 ( .A(n22305), .B(n22304), .Z(n22306) );
  NAND U23316 ( .A(n22307), .B(n22306), .Z(n22333) );
  XNOR U23317 ( .A(n22334), .B(n22333), .Z(n22319) );
  NANDN U23318 ( .A(n22309), .B(n22308), .Z(n22313) );
  OR U23319 ( .A(n22311), .B(n22310), .Z(n22312) );
  NAND U23320 ( .A(n22313), .B(n22312), .Z(n22320) );
  XNOR U23321 ( .A(n22319), .B(n22320), .Z(n22321) );
  XNOR U23322 ( .A(n22322), .B(n22321), .Z(n22314) );
  XOR U23323 ( .A(sreg[1963]), .B(n22314), .Z(n22316) );
  XNOR U23324 ( .A(n22315), .B(n22316), .Z(c[1963]) );
  OR U23325 ( .A(n22314), .B(sreg[1963]), .Z(n22318) );
  NAND U23326 ( .A(n22316), .B(n22315), .Z(n22317) );
  NAND U23327 ( .A(n22318), .B(n22317), .Z(n22357) );
  NANDN U23328 ( .A(n22320), .B(n22319), .Z(n22324) );
  NAND U23329 ( .A(n22322), .B(n22321), .Z(n22323) );
  NAND U23330 ( .A(n22324), .B(n22323), .Z(n22340) );
  AND U23331 ( .A(b[2]), .B(a[942]), .Z(n22346) );
  AND U23332 ( .A(a[943]), .B(b[1]), .Z(n22344) );
  AND U23333 ( .A(a[941]), .B(b[3]), .Z(n22343) );
  XOR U23334 ( .A(n22344), .B(n22343), .Z(n22345) );
  XOR U23335 ( .A(n22346), .B(n22345), .Z(n22349) );
  NAND U23336 ( .A(b[0]), .B(a[944]), .Z(n22350) );
  XOR U23337 ( .A(n22349), .B(n22350), .Z(n22352) );
  OR U23338 ( .A(n22326), .B(n22325), .Z(n22330) );
  NANDN U23339 ( .A(n22328), .B(n22327), .Z(n22329) );
  NAND U23340 ( .A(n22330), .B(n22329), .Z(n22351) );
  XNOR U23341 ( .A(n22352), .B(n22351), .Z(n22337) );
  NANDN U23342 ( .A(n22332), .B(n22331), .Z(n22336) );
  OR U23343 ( .A(n22334), .B(n22333), .Z(n22335) );
  NAND U23344 ( .A(n22336), .B(n22335), .Z(n22338) );
  XNOR U23345 ( .A(n22337), .B(n22338), .Z(n22339) );
  XNOR U23346 ( .A(n22340), .B(n22339), .Z(n22355) );
  XNOR U23347 ( .A(n22355), .B(sreg[1964]), .Z(n22356) );
  XOR U23348 ( .A(n22357), .B(n22356), .Z(c[1964]) );
  NANDN U23349 ( .A(n22338), .B(n22337), .Z(n22342) );
  NAND U23350 ( .A(n22340), .B(n22339), .Z(n22341) );
  NAND U23351 ( .A(n22342), .B(n22341), .Z(n22368) );
  AND U23352 ( .A(b[2]), .B(a[943]), .Z(n22374) );
  AND U23353 ( .A(a[944]), .B(b[1]), .Z(n22372) );
  AND U23354 ( .A(a[942]), .B(b[3]), .Z(n22371) );
  XOR U23355 ( .A(n22372), .B(n22371), .Z(n22373) );
  XOR U23356 ( .A(n22374), .B(n22373), .Z(n22377) );
  NAND U23357 ( .A(b[0]), .B(a[945]), .Z(n22378) );
  XOR U23358 ( .A(n22377), .B(n22378), .Z(n22380) );
  OR U23359 ( .A(n22344), .B(n22343), .Z(n22348) );
  NANDN U23360 ( .A(n22346), .B(n22345), .Z(n22347) );
  NAND U23361 ( .A(n22348), .B(n22347), .Z(n22379) );
  XNOR U23362 ( .A(n22380), .B(n22379), .Z(n22365) );
  NANDN U23363 ( .A(n22350), .B(n22349), .Z(n22354) );
  OR U23364 ( .A(n22352), .B(n22351), .Z(n22353) );
  NAND U23365 ( .A(n22354), .B(n22353), .Z(n22366) );
  XNOR U23366 ( .A(n22365), .B(n22366), .Z(n22367) );
  XNOR U23367 ( .A(n22368), .B(n22367), .Z(n22360) );
  XNOR U23368 ( .A(n22360), .B(sreg[1965]), .Z(n22362) );
  NAND U23369 ( .A(n22355), .B(sreg[1964]), .Z(n22359) );
  OR U23370 ( .A(n22357), .B(n22356), .Z(n22358) );
  AND U23371 ( .A(n22359), .B(n22358), .Z(n22361) );
  XOR U23372 ( .A(n22362), .B(n22361), .Z(c[1965]) );
  NAND U23373 ( .A(n22360), .B(sreg[1965]), .Z(n22364) );
  OR U23374 ( .A(n22362), .B(n22361), .Z(n22363) );
  NAND U23375 ( .A(n22364), .B(n22363), .Z(n22403) );
  NANDN U23376 ( .A(n22366), .B(n22365), .Z(n22370) );
  NAND U23377 ( .A(n22368), .B(n22367), .Z(n22369) );
  NAND U23378 ( .A(n22370), .B(n22369), .Z(n22386) );
  AND U23379 ( .A(b[2]), .B(a[944]), .Z(n22392) );
  AND U23380 ( .A(a[945]), .B(b[1]), .Z(n22390) );
  AND U23381 ( .A(a[943]), .B(b[3]), .Z(n22389) );
  XOR U23382 ( .A(n22390), .B(n22389), .Z(n22391) );
  XOR U23383 ( .A(n22392), .B(n22391), .Z(n22395) );
  NAND U23384 ( .A(b[0]), .B(a[946]), .Z(n22396) );
  XOR U23385 ( .A(n22395), .B(n22396), .Z(n22398) );
  OR U23386 ( .A(n22372), .B(n22371), .Z(n22376) );
  NANDN U23387 ( .A(n22374), .B(n22373), .Z(n22375) );
  NAND U23388 ( .A(n22376), .B(n22375), .Z(n22397) );
  XNOR U23389 ( .A(n22398), .B(n22397), .Z(n22383) );
  NANDN U23390 ( .A(n22378), .B(n22377), .Z(n22382) );
  OR U23391 ( .A(n22380), .B(n22379), .Z(n22381) );
  NAND U23392 ( .A(n22382), .B(n22381), .Z(n22384) );
  XNOR U23393 ( .A(n22383), .B(n22384), .Z(n22385) );
  XNOR U23394 ( .A(n22386), .B(n22385), .Z(n22401) );
  XOR U23395 ( .A(sreg[1966]), .B(n22401), .Z(n22402) );
  XOR U23396 ( .A(n22403), .B(n22402), .Z(c[1966]) );
  NANDN U23397 ( .A(n22384), .B(n22383), .Z(n22388) );
  NAND U23398 ( .A(n22386), .B(n22385), .Z(n22387) );
  NAND U23399 ( .A(n22388), .B(n22387), .Z(n22412) );
  AND U23400 ( .A(b[2]), .B(a[945]), .Z(n22418) );
  AND U23401 ( .A(a[946]), .B(b[1]), .Z(n22416) );
  AND U23402 ( .A(a[944]), .B(b[3]), .Z(n22415) );
  XOR U23403 ( .A(n22416), .B(n22415), .Z(n22417) );
  XOR U23404 ( .A(n22418), .B(n22417), .Z(n22421) );
  NAND U23405 ( .A(b[0]), .B(a[947]), .Z(n22422) );
  XOR U23406 ( .A(n22421), .B(n22422), .Z(n22424) );
  OR U23407 ( .A(n22390), .B(n22389), .Z(n22394) );
  NANDN U23408 ( .A(n22392), .B(n22391), .Z(n22393) );
  NAND U23409 ( .A(n22394), .B(n22393), .Z(n22423) );
  XNOR U23410 ( .A(n22424), .B(n22423), .Z(n22409) );
  NANDN U23411 ( .A(n22396), .B(n22395), .Z(n22400) );
  OR U23412 ( .A(n22398), .B(n22397), .Z(n22399) );
  NAND U23413 ( .A(n22400), .B(n22399), .Z(n22410) );
  XNOR U23414 ( .A(n22409), .B(n22410), .Z(n22411) );
  XOR U23415 ( .A(n22412), .B(n22411), .Z(n22408) );
  OR U23416 ( .A(n22401), .B(sreg[1966]), .Z(n22405) );
  NANDN U23417 ( .A(n22403), .B(n22402), .Z(n22404) );
  AND U23418 ( .A(n22405), .B(n22404), .Z(n22407) );
  XNOR U23419 ( .A(sreg[1967]), .B(n22407), .Z(n22406) );
  XOR U23420 ( .A(n22408), .B(n22406), .Z(c[1967]) );
  NANDN U23421 ( .A(n22410), .B(n22409), .Z(n22414) );
  NAND U23422 ( .A(n22412), .B(n22411), .Z(n22413) );
  NAND U23423 ( .A(n22414), .B(n22413), .Z(n22430) );
  AND U23424 ( .A(b[2]), .B(a[946]), .Z(n22442) );
  AND U23425 ( .A(a[947]), .B(b[1]), .Z(n22440) );
  AND U23426 ( .A(a[945]), .B(b[3]), .Z(n22439) );
  XOR U23427 ( .A(n22440), .B(n22439), .Z(n22441) );
  XOR U23428 ( .A(n22442), .B(n22441), .Z(n22433) );
  NAND U23429 ( .A(b[0]), .B(a[948]), .Z(n22434) );
  XOR U23430 ( .A(n22433), .B(n22434), .Z(n22436) );
  OR U23431 ( .A(n22416), .B(n22415), .Z(n22420) );
  NANDN U23432 ( .A(n22418), .B(n22417), .Z(n22419) );
  NAND U23433 ( .A(n22420), .B(n22419), .Z(n22435) );
  XNOR U23434 ( .A(n22436), .B(n22435), .Z(n22427) );
  NANDN U23435 ( .A(n22422), .B(n22421), .Z(n22426) );
  OR U23436 ( .A(n22424), .B(n22423), .Z(n22425) );
  NAND U23437 ( .A(n22426), .B(n22425), .Z(n22428) );
  XNOR U23438 ( .A(n22427), .B(n22428), .Z(n22429) );
  XNOR U23439 ( .A(n22430), .B(n22429), .Z(n22445) );
  XNOR U23440 ( .A(n22445), .B(sreg[1968]), .Z(n22446) );
  XOR U23441 ( .A(n22447), .B(n22446), .Z(c[1968]) );
  NANDN U23442 ( .A(n22428), .B(n22427), .Z(n22432) );
  NAND U23443 ( .A(n22430), .B(n22429), .Z(n22431) );
  NAND U23444 ( .A(n22432), .B(n22431), .Z(n22470) );
  NANDN U23445 ( .A(n22434), .B(n22433), .Z(n22438) );
  OR U23446 ( .A(n22436), .B(n22435), .Z(n22437) );
  NAND U23447 ( .A(n22438), .B(n22437), .Z(n22467) );
  AND U23448 ( .A(b[2]), .B(a[947]), .Z(n22458) );
  AND U23449 ( .A(a[948]), .B(b[1]), .Z(n22456) );
  AND U23450 ( .A(a[946]), .B(b[3]), .Z(n22455) );
  XOR U23451 ( .A(n22456), .B(n22455), .Z(n22457) );
  XOR U23452 ( .A(n22458), .B(n22457), .Z(n22461) );
  NAND U23453 ( .A(b[0]), .B(a[949]), .Z(n22462) );
  XNOR U23454 ( .A(n22461), .B(n22462), .Z(n22463) );
  OR U23455 ( .A(n22440), .B(n22439), .Z(n22444) );
  NANDN U23456 ( .A(n22442), .B(n22441), .Z(n22443) );
  AND U23457 ( .A(n22444), .B(n22443), .Z(n22464) );
  XNOR U23458 ( .A(n22463), .B(n22464), .Z(n22468) );
  XNOR U23459 ( .A(n22467), .B(n22468), .Z(n22469) );
  XNOR U23460 ( .A(n22470), .B(n22469), .Z(n22450) );
  XOR U23461 ( .A(sreg[1969]), .B(n22450), .Z(n22451) );
  NAND U23462 ( .A(n22445), .B(sreg[1968]), .Z(n22449) );
  OR U23463 ( .A(n22447), .B(n22446), .Z(n22448) );
  NAND U23464 ( .A(n22449), .B(n22448), .Z(n22452) );
  XOR U23465 ( .A(n22451), .B(n22452), .Z(c[1969]) );
  OR U23466 ( .A(n22450), .B(sreg[1969]), .Z(n22454) );
  NANDN U23467 ( .A(n22452), .B(n22451), .Z(n22453) );
  AND U23468 ( .A(n22454), .B(n22453), .Z(n22475) );
  AND U23469 ( .A(b[2]), .B(a[948]), .Z(n22485) );
  AND U23470 ( .A(a[949]), .B(b[1]), .Z(n22483) );
  AND U23471 ( .A(a[947]), .B(b[3]), .Z(n22482) );
  XOR U23472 ( .A(n22483), .B(n22482), .Z(n22484) );
  XOR U23473 ( .A(n22485), .B(n22484), .Z(n22488) );
  NAND U23474 ( .A(b[0]), .B(a[950]), .Z(n22489) );
  XOR U23475 ( .A(n22488), .B(n22489), .Z(n22491) );
  OR U23476 ( .A(n22456), .B(n22455), .Z(n22460) );
  NANDN U23477 ( .A(n22458), .B(n22457), .Z(n22459) );
  NAND U23478 ( .A(n22460), .B(n22459), .Z(n22490) );
  XNOR U23479 ( .A(n22491), .B(n22490), .Z(n22476) );
  NANDN U23480 ( .A(n22462), .B(n22461), .Z(n22466) );
  NAND U23481 ( .A(n22464), .B(n22463), .Z(n22465) );
  NAND U23482 ( .A(n22466), .B(n22465), .Z(n22477) );
  XNOR U23483 ( .A(n22476), .B(n22477), .Z(n22478) );
  NANDN U23484 ( .A(n22468), .B(n22467), .Z(n22472) );
  NANDN U23485 ( .A(n22470), .B(n22469), .Z(n22471) );
  AND U23486 ( .A(n22472), .B(n22471), .Z(n22479) );
  XNOR U23487 ( .A(n22478), .B(n22479), .Z(n22474) );
  XOR U23488 ( .A(n22474), .B(sreg[1970]), .Z(n22473) );
  XOR U23489 ( .A(n22475), .B(n22473), .Z(c[1970]) );
  NANDN U23490 ( .A(n22477), .B(n22476), .Z(n22481) );
  NAND U23491 ( .A(n22479), .B(n22478), .Z(n22480) );
  NAND U23492 ( .A(n22481), .B(n22480), .Z(n22509) );
  AND U23493 ( .A(b[2]), .B(a[949]), .Z(n22503) );
  AND U23494 ( .A(a[950]), .B(b[1]), .Z(n22501) );
  AND U23495 ( .A(a[948]), .B(b[3]), .Z(n22500) );
  XOR U23496 ( .A(n22501), .B(n22500), .Z(n22502) );
  XOR U23497 ( .A(n22503), .B(n22502), .Z(n22494) );
  NAND U23498 ( .A(b[0]), .B(a[951]), .Z(n22495) );
  XOR U23499 ( .A(n22494), .B(n22495), .Z(n22497) );
  OR U23500 ( .A(n22483), .B(n22482), .Z(n22487) );
  NANDN U23501 ( .A(n22485), .B(n22484), .Z(n22486) );
  NAND U23502 ( .A(n22487), .B(n22486), .Z(n22496) );
  XNOR U23503 ( .A(n22497), .B(n22496), .Z(n22506) );
  NANDN U23504 ( .A(n22489), .B(n22488), .Z(n22493) );
  OR U23505 ( .A(n22491), .B(n22490), .Z(n22492) );
  NAND U23506 ( .A(n22493), .B(n22492), .Z(n22507) );
  XNOR U23507 ( .A(n22506), .B(n22507), .Z(n22508) );
  XOR U23508 ( .A(n22509), .B(n22508), .Z(n22512) );
  XOR U23509 ( .A(sreg[1971]), .B(n22512), .Z(n22514) );
  XNOR U23510 ( .A(n22513), .B(n22514), .Z(c[1971]) );
  NANDN U23511 ( .A(n22495), .B(n22494), .Z(n22499) );
  OR U23512 ( .A(n22497), .B(n22496), .Z(n22498) );
  NAND U23513 ( .A(n22499), .B(n22498), .Z(n22534) );
  AND U23514 ( .A(b[2]), .B(a[950]), .Z(n22525) );
  AND U23515 ( .A(a[951]), .B(b[1]), .Z(n22523) );
  AND U23516 ( .A(a[949]), .B(b[3]), .Z(n22522) );
  XOR U23517 ( .A(n22523), .B(n22522), .Z(n22524) );
  XOR U23518 ( .A(n22525), .B(n22524), .Z(n22528) );
  NAND U23519 ( .A(b[0]), .B(a[952]), .Z(n22529) );
  XNOR U23520 ( .A(n22528), .B(n22529), .Z(n22530) );
  OR U23521 ( .A(n22501), .B(n22500), .Z(n22505) );
  NANDN U23522 ( .A(n22503), .B(n22502), .Z(n22504) );
  AND U23523 ( .A(n22505), .B(n22504), .Z(n22531) );
  XNOR U23524 ( .A(n22530), .B(n22531), .Z(n22535) );
  XNOR U23525 ( .A(n22534), .B(n22535), .Z(n22536) );
  NANDN U23526 ( .A(n22507), .B(n22506), .Z(n22511) );
  NAND U23527 ( .A(n22509), .B(n22508), .Z(n22510) );
  NAND U23528 ( .A(n22511), .B(n22510), .Z(n22537) );
  XNOR U23529 ( .A(n22536), .B(n22537), .Z(n22517) );
  XOR U23530 ( .A(sreg[1972]), .B(n22517), .Z(n22518) );
  NANDN U23531 ( .A(n22512), .B(sreg[1971]), .Z(n22516) );
  NANDN U23532 ( .A(n22514), .B(n22513), .Z(n22515) );
  NAND U23533 ( .A(n22516), .B(n22515), .Z(n22519) );
  XOR U23534 ( .A(n22518), .B(n22519), .Z(c[1972]) );
  OR U23535 ( .A(n22517), .B(sreg[1972]), .Z(n22521) );
  NANDN U23536 ( .A(n22519), .B(n22518), .Z(n22520) );
  AND U23537 ( .A(n22521), .B(n22520), .Z(n22541) );
  AND U23538 ( .A(b[2]), .B(a[951]), .Z(n22552) );
  AND U23539 ( .A(a[952]), .B(b[1]), .Z(n22550) );
  AND U23540 ( .A(a[950]), .B(b[3]), .Z(n22549) );
  XOR U23541 ( .A(n22550), .B(n22549), .Z(n22551) );
  XOR U23542 ( .A(n22552), .B(n22551), .Z(n22555) );
  NAND U23543 ( .A(b[0]), .B(a[953]), .Z(n22556) );
  XOR U23544 ( .A(n22555), .B(n22556), .Z(n22558) );
  OR U23545 ( .A(n22523), .B(n22522), .Z(n22527) );
  NANDN U23546 ( .A(n22525), .B(n22524), .Z(n22526) );
  NAND U23547 ( .A(n22527), .B(n22526), .Z(n22557) );
  XNOR U23548 ( .A(n22558), .B(n22557), .Z(n22543) );
  NANDN U23549 ( .A(n22529), .B(n22528), .Z(n22533) );
  NAND U23550 ( .A(n22531), .B(n22530), .Z(n22532) );
  NAND U23551 ( .A(n22533), .B(n22532), .Z(n22544) );
  XNOR U23552 ( .A(n22543), .B(n22544), .Z(n22545) );
  NANDN U23553 ( .A(n22535), .B(n22534), .Z(n22539) );
  NANDN U23554 ( .A(n22537), .B(n22536), .Z(n22538) );
  AND U23555 ( .A(n22539), .B(n22538), .Z(n22546) );
  XNOR U23556 ( .A(n22545), .B(n22546), .Z(n22542) );
  XOR U23557 ( .A(sreg[1973]), .B(n22542), .Z(n22540) );
  XOR U23558 ( .A(n22541), .B(n22540), .Z(c[1973]) );
  NANDN U23559 ( .A(n22544), .B(n22543), .Z(n22548) );
  NAND U23560 ( .A(n22546), .B(n22545), .Z(n22547) );
  NAND U23561 ( .A(n22548), .B(n22547), .Z(n22564) );
  AND U23562 ( .A(b[2]), .B(a[952]), .Z(n22570) );
  AND U23563 ( .A(a[953]), .B(b[1]), .Z(n22568) );
  AND U23564 ( .A(a[951]), .B(b[3]), .Z(n22567) );
  XOR U23565 ( .A(n22568), .B(n22567), .Z(n22569) );
  XOR U23566 ( .A(n22570), .B(n22569), .Z(n22573) );
  NAND U23567 ( .A(b[0]), .B(a[954]), .Z(n22574) );
  XOR U23568 ( .A(n22573), .B(n22574), .Z(n22576) );
  OR U23569 ( .A(n22550), .B(n22549), .Z(n22554) );
  NANDN U23570 ( .A(n22552), .B(n22551), .Z(n22553) );
  NAND U23571 ( .A(n22554), .B(n22553), .Z(n22575) );
  XNOR U23572 ( .A(n22576), .B(n22575), .Z(n22561) );
  NANDN U23573 ( .A(n22556), .B(n22555), .Z(n22560) );
  OR U23574 ( .A(n22558), .B(n22557), .Z(n22559) );
  NAND U23575 ( .A(n22560), .B(n22559), .Z(n22562) );
  XNOR U23576 ( .A(n22561), .B(n22562), .Z(n22563) );
  XNOR U23577 ( .A(n22564), .B(n22563), .Z(n22579) );
  XNOR U23578 ( .A(n22579), .B(sreg[1974]), .Z(n22581) );
  XNOR U23579 ( .A(n22580), .B(n22581), .Z(c[1974]) );
  NANDN U23580 ( .A(n22562), .B(n22561), .Z(n22566) );
  NAND U23581 ( .A(n22564), .B(n22563), .Z(n22565) );
  NAND U23582 ( .A(n22566), .B(n22565), .Z(n22590) );
  AND U23583 ( .A(b[2]), .B(a[953]), .Z(n22596) );
  AND U23584 ( .A(a[954]), .B(b[1]), .Z(n22594) );
  AND U23585 ( .A(a[952]), .B(b[3]), .Z(n22593) );
  XOR U23586 ( .A(n22594), .B(n22593), .Z(n22595) );
  XOR U23587 ( .A(n22596), .B(n22595), .Z(n22599) );
  NAND U23588 ( .A(b[0]), .B(a[955]), .Z(n22600) );
  XOR U23589 ( .A(n22599), .B(n22600), .Z(n22602) );
  OR U23590 ( .A(n22568), .B(n22567), .Z(n22572) );
  NANDN U23591 ( .A(n22570), .B(n22569), .Z(n22571) );
  NAND U23592 ( .A(n22572), .B(n22571), .Z(n22601) );
  XNOR U23593 ( .A(n22602), .B(n22601), .Z(n22587) );
  NANDN U23594 ( .A(n22574), .B(n22573), .Z(n22578) );
  OR U23595 ( .A(n22576), .B(n22575), .Z(n22577) );
  NAND U23596 ( .A(n22578), .B(n22577), .Z(n22588) );
  XNOR U23597 ( .A(n22587), .B(n22588), .Z(n22589) );
  XOR U23598 ( .A(n22590), .B(n22589), .Z(n22586) );
  NAND U23599 ( .A(n22579), .B(sreg[1974]), .Z(n22583) );
  NANDN U23600 ( .A(n22581), .B(n22580), .Z(n22582) );
  NAND U23601 ( .A(n22583), .B(n22582), .Z(n22585) );
  XNOR U23602 ( .A(sreg[1975]), .B(n22585), .Z(n22584) );
  XOR U23603 ( .A(n22586), .B(n22584), .Z(c[1975]) );
  NANDN U23604 ( .A(n22588), .B(n22587), .Z(n22592) );
  NAND U23605 ( .A(n22590), .B(n22589), .Z(n22591) );
  NAND U23606 ( .A(n22592), .B(n22591), .Z(n22608) );
  AND U23607 ( .A(b[2]), .B(a[954]), .Z(n22614) );
  AND U23608 ( .A(a[955]), .B(b[1]), .Z(n22612) );
  AND U23609 ( .A(a[953]), .B(b[3]), .Z(n22611) );
  XOR U23610 ( .A(n22612), .B(n22611), .Z(n22613) );
  XOR U23611 ( .A(n22614), .B(n22613), .Z(n22617) );
  NAND U23612 ( .A(b[0]), .B(a[956]), .Z(n22618) );
  XOR U23613 ( .A(n22617), .B(n22618), .Z(n22620) );
  OR U23614 ( .A(n22594), .B(n22593), .Z(n22598) );
  NANDN U23615 ( .A(n22596), .B(n22595), .Z(n22597) );
  NAND U23616 ( .A(n22598), .B(n22597), .Z(n22619) );
  XNOR U23617 ( .A(n22620), .B(n22619), .Z(n22605) );
  NANDN U23618 ( .A(n22600), .B(n22599), .Z(n22604) );
  OR U23619 ( .A(n22602), .B(n22601), .Z(n22603) );
  NAND U23620 ( .A(n22604), .B(n22603), .Z(n22606) );
  XNOR U23621 ( .A(n22605), .B(n22606), .Z(n22607) );
  XNOR U23622 ( .A(n22608), .B(n22607), .Z(n22623) );
  XOR U23623 ( .A(sreg[1976]), .B(n22623), .Z(n22625) );
  XNOR U23624 ( .A(n22624), .B(n22625), .Z(c[1976]) );
  NANDN U23625 ( .A(n22606), .B(n22605), .Z(n22610) );
  NAND U23626 ( .A(n22608), .B(n22607), .Z(n22609) );
  NAND U23627 ( .A(n22610), .B(n22609), .Z(n22634) );
  AND U23628 ( .A(b[2]), .B(a[955]), .Z(n22640) );
  AND U23629 ( .A(a[956]), .B(b[1]), .Z(n22638) );
  AND U23630 ( .A(a[954]), .B(b[3]), .Z(n22637) );
  XOR U23631 ( .A(n22638), .B(n22637), .Z(n22639) );
  XOR U23632 ( .A(n22640), .B(n22639), .Z(n22643) );
  NAND U23633 ( .A(b[0]), .B(a[957]), .Z(n22644) );
  XOR U23634 ( .A(n22643), .B(n22644), .Z(n22646) );
  OR U23635 ( .A(n22612), .B(n22611), .Z(n22616) );
  NANDN U23636 ( .A(n22614), .B(n22613), .Z(n22615) );
  NAND U23637 ( .A(n22616), .B(n22615), .Z(n22645) );
  XNOR U23638 ( .A(n22646), .B(n22645), .Z(n22631) );
  NANDN U23639 ( .A(n22618), .B(n22617), .Z(n22622) );
  OR U23640 ( .A(n22620), .B(n22619), .Z(n22621) );
  NAND U23641 ( .A(n22622), .B(n22621), .Z(n22632) );
  XNOR U23642 ( .A(n22631), .B(n22632), .Z(n22633) );
  XOR U23643 ( .A(n22634), .B(n22633), .Z(n22630) );
  OR U23644 ( .A(n22623), .B(sreg[1976]), .Z(n22627) );
  NAND U23645 ( .A(n22625), .B(n22624), .Z(n22626) );
  AND U23646 ( .A(n22627), .B(n22626), .Z(n22629) );
  XNOR U23647 ( .A(sreg[1977]), .B(n22629), .Z(n22628) );
  XOR U23648 ( .A(n22630), .B(n22628), .Z(c[1977]) );
  NANDN U23649 ( .A(n22632), .B(n22631), .Z(n22636) );
  NAND U23650 ( .A(n22634), .B(n22633), .Z(n22635) );
  NAND U23651 ( .A(n22636), .B(n22635), .Z(n22652) );
  AND U23652 ( .A(b[2]), .B(a[956]), .Z(n22658) );
  AND U23653 ( .A(a[957]), .B(b[1]), .Z(n22656) );
  AND U23654 ( .A(a[955]), .B(b[3]), .Z(n22655) );
  XOR U23655 ( .A(n22656), .B(n22655), .Z(n22657) );
  XOR U23656 ( .A(n22658), .B(n22657), .Z(n22661) );
  NAND U23657 ( .A(b[0]), .B(a[958]), .Z(n22662) );
  XOR U23658 ( .A(n22661), .B(n22662), .Z(n22664) );
  OR U23659 ( .A(n22638), .B(n22637), .Z(n22642) );
  NANDN U23660 ( .A(n22640), .B(n22639), .Z(n22641) );
  NAND U23661 ( .A(n22642), .B(n22641), .Z(n22663) );
  XNOR U23662 ( .A(n22664), .B(n22663), .Z(n22649) );
  NANDN U23663 ( .A(n22644), .B(n22643), .Z(n22648) );
  OR U23664 ( .A(n22646), .B(n22645), .Z(n22647) );
  NAND U23665 ( .A(n22648), .B(n22647), .Z(n22650) );
  XNOR U23666 ( .A(n22649), .B(n22650), .Z(n22651) );
  XNOR U23667 ( .A(n22652), .B(n22651), .Z(n22667) );
  XNOR U23668 ( .A(n22667), .B(sreg[1978]), .Z(n22668) );
  XOR U23669 ( .A(n22669), .B(n22668), .Z(c[1978]) );
  NANDN U23670 ( .A(n22650), .B(n22649), .Z(n22654) );
  NAND U23671 ( .A(n22652), .B(n22651), .Z(n22653) );
  NAND U23672 ( .A(n22654), .B(n22653), .Z(n22675) );
  AND U23673 ( .A(b[2]), .B(a[957]), .Z(n22681) );
  AND U23674 ( .A(a[958]), .B(b[1]), .Z(n22679) );
  AND U23675 ( .A(a[956]), .B(b[3]), .Z(n22678) );
  XOR U23676 ( .A(n22679), .B(n22678), .Z(n22680) );
  XOR U23677 ( .A(n22681), .B(n22680), .Z(n22684) );
  NAND U23678 ( .A(b[0]), .B(a[959]), .Z(n22685) );
  XOR U23679 ( .A(n22684), .B(n22685), .Z(n22687) );
  OR U23680 ( .A(n22656), .B(n22655), .Z(n22660) );
  NANDN U23681 ( .A(n22658), .B(n22657), .Z(n22659) );
  NAND U23682 ( .A(n22660), .B(n22659), .Z(n22686) );
  XNOR U23683 ( .A(n22687), .B(n22686), .Z(n22672) );
  NANDN U23684 ( .A(n22662), .B(n22661), .Z(n22666) );
  OR U23685 ( .A(n22664), .B(n22663), .Z(n22665) );
  NAND U23686 ( .A(n22666), .B(n22665), .Z(n22673) );
  XNOR U23687 ( .A(n22672), .B(n22673), .Z(n22674) );
  XNOR U23688 ( .A(n22675), .B(n22674), .Z(n22690) );
  XOR U23689 ( .A(sreg[1979]), .B(n22690), .Z(n22691) );
  NAND U23690 ( .A(n22667), .B(sreg[1978]), .Z(n22671) );
  OR U23691 ( .A(n22669), .B(n22668), .Z(n22670) );
  NAND U23692 ( .A(n22671), .B(n22670), .Z(n22692) );
  XOR U23693 ( .A(n22691), .B(n22692), .Z(c[1979]) );
  NANDN U23694 ( .A(n22673), .B(n22672), .Z(n22677) );
  NAND U23695 ( .A(n22675), .B(n22674), .Z(n22676) );
  NAND U23696 ( .A(n22677), .B(n22676), .Z(n22701) );
  AND U23697 ( .A(b[2]), .B(a[958]), .Z(n22707) );
  AND U23698 ( .A(a[959]), .B(b[1]), .Z(n22705) );
  AND U23699 ( .A(a[957]), .B(b[3]), .Z(n22704) );
  XOR U23700 ( .A(n22705), .B(n22704), .Z(n22706) );
  XOR U23701 ( .A(n22707), .B(n22706), .Z(n22710) );
  NAND U23702 ( .A(b[0]), .B(a[960]), .Z(n22711) );
  XOR U23703 ( .A(n22710), .B(n22711), .Z(n22713) );
  OR U23704 ( .A(n22679), .B(n22678), .Z(n22683) );
  NANDN U23705 ( .A(n22681), .B(n22680), .Z(n22682) );
  NAND U23706 ( .A(n22683), .B(n22682), .Z(n22712) );
  XNOR U23707 ( .A(n22713), .B(n22712), .Z(n22698) );
  NANDN U23708 ( .A(n22685), .B(n22684), .Z(n22689) );
  OR U23709 ( .A(n22687), .B(n22686), .Z(n22688) );
  NAND U23710 ( .A(n22689), .B(n22688), .Z(n22699) );
  XNOR U23711 ( .A(n22698), .B(n22699), .Z(n22700) );
  XOR U23712 ( .A(n22701), .B(n22700), .Z(n22697) );
  OR U23713 ( .A(n22690), .B(sreg[1979]), .Z(n22694) );
  NANDN U23714 ( .A(n22692), .B(n22691), .Z(n22693) );
  AND U23715 ( .A(n22694), .B(n22693), .Z(n22696) );
  XNOR U23716 ( .A(sreg[1980]), .B(n22696), .Z(n22695) );
  XOR U23717 ( .A(n22697), .B(n22695), .Z(c[1980]) );
  NANDN U23718 ( .A(n22699), .B(n22698), .Z(n22703) );
  NAND U23719 ( .A(n22701), .B(n22700), .Z(n22702) );
  NAND U23720 ( .A(n22703), .B(n22702), .Z(n22719) );
  AND U23721 ( .A(b[2]), .B(a[959]), .Z(n22725) );
  AND U23722 ( .A(a[960]), .B(b[1]), .Z(n22723) );
  AND U23723 ( .A(a[958]), .B(b[3]), .Z(n22722) );
  XOR U23724 ( .A(n22723), .B(n22722), .Z(n22724) );
  XOR U23725 ( .A(n22725), .B(n22724), .Z(n22728) );
  NAND U23726 ( .A(b[0]), .B(a[961]), .Z(n22729) );
  XOR U23727 ( .A(n22728), .B(n22729), .Z(n22731) );
  OR U23728 ( .A(n22705), .B(n22704), .Z(n22709) );
  NANDN U23729 ( .A(n22707), .B(n22706), .Z(n22708) );
  NAND U23730 ( .A(n22709), .B(n22708), .Z(n22730) );
  XNOR U23731 ( .A(n22731), .B(n22730), .Z(n22716) );
  NANDN U23732 ( .A(n22711), .B(n22710), .Z(n22715) );
  OR U23733 ( .A(n22713), .B(n22712), .Z(n22714) );
  NAND U23734 ( .A(n22715), .B(n22714), .Z(n22717) );
  XNOR U23735 ( .A(n22716), .B(n22717), .Z(n22718) );
  XNOR U23736 ( .A(n22719), .B(n22718), .Z(n22734) );
  XNOR U23737 ( .A(n22734), .B(sreg[1981]), .Z(n22735) );
  XOR U23738 ( .A(n22736), .B(n22735), .Z(c[1981]) );
  NANDN U23739 ( .A(n22717), .B(n22716), .Z(n22721) );
  NAND U23740 ( .A(n22719), .B(n22718), .Z(n22720) );
  NAND U23741 ( .A(n22721), .B(n22720), .Z(n22745) );
  AND U23742 ( .A(b[2]), .B(a[960]), .Z(n22751) );
  AND U23743 ( .A(a[961]), .B(b[1]), .Z(n22749) );
  AND U23744 ( .A(a[959]), .B(b[3]), .Z(n22748) );
  XOR U23745 ( .A(n22749), .B(n22748), .Z(n22750) );
  XOR U23746 ( .A(n22751), .B(n22750), .Z(n22754) );
  NAND U23747 ( .A(b[0]), .B(a[962]), .Z(n22755) );
  XOR U23748 ( .A(n22754), .B(n22755), .Z(n22757) );
  OR U23749 ( .A(n22723), .B(n22722), .Z(n22727) );
  NANDN U23750 ( .A(n22725), .B(n22724), .Z(n22726) );
  NAND U23751 ( .A(n22727), .B(n22726), .Z(n22756) );
  XNOR U23752 ( .A(n22757), .B(n22756), .Z(n22742) );
  NANDN U23753 ( .A(n22729), .B(n22728), .Z(n22733) );
  OR U23754 ( .A(n22731), .B(n22730), .Z(n22732) );
  NAND U23755 ( .A(n22733), .B(n22732), .Z(n22743) );
  XNOR U23756 ( .A(n22742), .B(n22743), .Z(n22744) );
  XOR U23757 ( .A(n22745), .B(n22744), .Z(n22741) );
  NAND U23758 ( .A(n22734), .B(sreg[1981]), .Z(n22738) );
  OR U23759 ( .A(n22736), .B(n22735), .Z(n22737) );
  NAND U23760 ( .A(n22738), .B(n22737), .Z(n22740) );
  XNOR U23761 ( .A(sreg[1982]), .B(n22740), .Z(n22739) );
  XOR U23762 ( .A(n22741), .B(n22739), .Z(c[1982]) );
  NANDN U23763 ( .A(n22743), .B(n22742), .Z(n22747) );
  NAND U23764 ( .A(n22745), .B(n22744), .Z(n22746) );
  NAND U23765 ( .A(n22747), .B(n22746), .Z(n22763) );
  AND U23766 ( .A(b[2]), .B(a[961]), .Z(n22769) );
  AND U23767 ( .A(a[962]), .B(b[1]), .Z(n22767) );
  AND U23768 ( .A(a[960]), .B(b[3]), .Z(n22766) );
  XOR U23769 ( .A(n22767), .B(n22766), .Z(n22768) );
  XOR U23770 ( .A(n22769), .B(n22768), .Z(n22772) );
  NAND U23771 ( .A(b[0]), .B(a[963]), .Z(n22773) );
  XOR U23772 ( .A(n22772), .B(n22773), .Z(n22775) );
  OR U23773 ( .A(n22749), .B(n22748), .Z(n22753) );
  NANDN U23774 ( .A(n22751), .B(n22750), .Z(n22752) );
  NAND U23775 ( .A(n22753), .B(n22752), .Z(n22774) );
  XNOR U23776 ( .A(n22775), .B(n22774), .Z(n22760) );
  NANDN U23777 ( .A(n22755), .B(n22754), .Z(n22759) );
  OR U23778 ( .A(n22757), .B(n22756), .Z(n22758) );
  NAND U23779 ( .A(n22759), .B(n22758), .Z(n22761) );
  XNOR U23780 ( .A(n22760), .B(n22761), .Z(n22762) );
  XNOR U23781 ( .A(n22763), .B(n22762), .Z(n22778) );
  XNOR U23782 ( .A(n22778), .B(sreg[1983]), .Z(n22779) );
  XOR U23783 ( .A(n22780), .B(n22779), .Z(c[1983]) );
  NANDN U23784 ( .A(n22761), .B(n22760), .Z(n22765) );
  NAND U23785 ( .A(n22763), .B(n22762), .Z(n22764) );
  NAND U23786 ( .A(n22765), .B(n22764), .Z(n22789) );
  AND U23787 ( .A(b[2]), .B(a[962]), .Z(n22801) );
  AND U23788 ( .A(a[963]), .B(b[1]), .Z(n22799) );
  AND U23789 ( .A(a[961]), .B(b[3]), .Z(n22798) );
  XOR U23790 ( .A(n22799), .B(n22798), .Z(n22800) );
  XOR U23791 ( .A(n22801), .B(n22800), .Z(n22792) );
  NAND U23792 ( .A(b[0]), .B(a[964]), .Z(n22793) );
  XOR U23793 ( .A(n22792), .B(n22793), .Z(n22795) );
  OR U23794 ( .A(n22767), .B(n22766), .Z(n22771) );
  NANDN U23795 ( .A(n22769), .B(n22768), .Z(n22770) );
  NAND U23796 ( .A(n22771), .B(n22770), .Z(n22794) );
  XNOR U23797 ( .A(n22795), .B(n22794), .Z(n22786) );
  NANDN U23798 ( .A(n22773), .B(n22772), .Z(n22777) );
  OR U23799 ( .A(n22775), .B(n22774), .Z(n22776) );
  NAND U23800 ( .A(n22777), .B(n22776), .Z(n22787) );
  XNOR U23801 ( .A(n22786), .B(n22787), .Z(n22788) );
  XNOR U23802 ( .A(n22789), .B(n22788), .Z(n22785) );
  NAND U23803 ( .A(n22778), .B(sreg[1983]), .Z(n22782) );
  OR U23804 ( .A(n22780), .B(n22779), .Z(n22781) );
  AND U23805 ( .A(n22782), .B(n22781), .Z(n22784) );
  XNOR U23806 ( .A(n22784), .B(sreg[1984]), .Z(n22783) );
  XOR U23807 ( .A(n22785), .B(n22783), .Z(c[1984]) );
  NANDN U23808 ( .A(n22787), .B(n22786), .Z(n22791) );
  NAND U23809 ( .A(n22789), .B(n22788), .Z(n22790) );
  NAND U23810 ( .A(n22791), .B(n22790), .Z(n22819) );
  NANDN U23811 ( .A(n22793), .B(n22792), .Z(n22797) );
  OR U23812 ( .A(n22795), .B(n22794), .Z(n22796) );
  NAND U23813 ( .A(n22797), .B(n22796), .Z(n22816) );
  AND U23814 ( .A(b[2]), .B(a[963]), .Z(n22807) );
  AND U23815 ( .A(a[964]), .B(b[1]), .Z(n22805) );
  AND U23816 ( .A(a[962]), .B(b[3]), .Z(n22804) );
  XOR U23817 ( .A(n22805), .B(n22804), .Z(n22806) );
  XOR U23818 ( .A(n22807), .B(n22806), .Z(n22810) );
  NAND U23819 ( .A(b[0]), .B(a[965]), .Z(n22811) );
  XNOR U23820 ( .A(n22810), .B(n22811), .Z(n22812) );
  OR U23821 ( .A(n22799), .B(n22798), .Z(n22803) );
  NANDN U23822 ( .A(n22801), .B(n22800), .Z(n22802) );
  AND U23823 ( .A(n22803), .B(n22802), .Z(n22813) );
  XNOR U23824 ( .A(n22812), .B(n22813), .Z(n22817) );
  XNOR U23825 ( .A(n22816), .B(n22817), .Z(n22818) );
  XNOR U23826 ( .A(n22819), .B(n22818), .Z(n22822) );
  XNOR U23827 ( .A(sreg[1985]), .B(n22822), .Z(n22824) );
  XNOR U23828 ( .A(n22823), .B(n22824), .Z(c[1985]) );
  AND U23829 ( .A(b[2]), .B(a[964]), .Z(n22839) );
  AND U23830 ( .A(a[965]), .B(b[1]), .Z(n22837) );
  AND U23831 ( .A(a[963]), .B(b[3]), .Z(n22836) );
  XOR U23832 ( .A(n22837), .B(n22836), .Z(n22838) );
  XOR U23833 ( .A(n22839), .B(n22838), .Z(n22842) );
  NAND U23834 ( .A(b[0]), .B(a[966]), .Z(n22843) );
  XOR U23835 ( .A(n22842), .B(n22843), .Z(n22845) );
  OR U23836 ( .A(n22805), .B(n22804), .Z(n22809) );
  NANDN U23837 ( .A(n22807), .B(n22806), .Z(n22808) );
  NAND U23838 ( .A(n22809), .B(n22808), .Z(n22844) );
  XNOR U23839 ( .A(n22845), .B(n22844), .Z(n22830) );
  NANDN U23840 ( .A(n22811), .B(n22810), .Z(n22815) );
  NAND U23841 ( .A(n22813), .B(n22812), .Z(n22814) );
  NAND U23842 ( .A(n22815), .B(n22814), .Z(n22831) );
  XNOR U23843 ( .A(n22830), .B(n22831), .Z(n22832) );
  NANDN U23844 ( .A(n22817), .B(n22816), .Z(n22821) );
  NANDN U23845 ( .A(n22819), .B(n22818), .Z(n22820) );
  NAND U23846 ( .A(n22821), .B(n22820), .Z(n22833) );
  XOR U23847 ( .A(n22832), .B(n22833), .Z(n22829) );
  NAND U23848 ( .A(sreg[1985]), .B(n22822), .Z(n22826) );
  NANDN U23849 ( .A(n22824), .B(n22823), .Z(n22825) );
  NAND U23850 ( .A(n22826), .B(n22825), .Z(n22828) );
  XNOR U23851 ( .A(sreg[1986]), .B(n22828), .Z(n22827) );
  XNOR U23852 ( .A(n22829), .B(n22827), .Z(c[1986]) );
  NANDN U23853 ( .A(n22831), .B(n22830), .Z(n22835) );
  NANDN U23854 ( .A(n22833), .B(n22832), .Z(n22834) );
  NAND U23855 ( .A(n22835), .B(n22834), .Z(n22868) );
  AND U23856 ( .A(b[2]), .B(a[965]), .Z(n22862) );
  AND U23857 ( .A(a[966]), .B(b[1]), .Z(n22860) );
  AND U23858 ( .A(a[964]), .B(b[3]), .Z(n22859) );
  XOR U23859 ( .A(n22860), .B(n22859), .Z(n22861) );
  XOR U23860 ( .A(n22862), .B(n22861), .Z(n22853) );
  NAND U23861 ( .A(b[0]), .B(a[967]), .Z(n22854) );
  XOR U23862 ( .A(n22853), .B(n22854), .Z(n22856) );
  OR U23863 ( .A(n22837), .B(n22836), .Z(n22841) );
  NANDN U23864 ( .A(n22839), .B(n22838), .Z(n22840) );
  NAND U23865 ( .A(n22841), .B(n22840), .Z(n22855) );
  XNOR U23866 ( .A(n22856), .B(n22855), .Z(n22865) );
  NANDN U23867 ( .A(n22843), .B(n22842), .Z(n22847) );
  OR U23868 ( .A(n22845), .B(n22844), .Z(n22846) );
  NAND U23869 ( .A(n22847), .B(n22846), .Z(n22866) );
  XNOR U23870 ( .A(n22865), .B(n22866), .Z(n22867) );
  XNOR U23871 ( .A(n22868), .B(n22867), .Z(n22848) );
  XOR U23872 ( .A(sreg[1987]), .B(n22848), .Z(n22850) );
  XNOR U23873 ( .A(n22849), .B(n22850), .Z(c[1987]) );
  OR U23874 ( .A(n22848), .B(sreg[1987]), .Z(n22852) );
  NAND U23875 ( .A(n22850), .B(n22849), .Z(n22851) );
  NAND U23876 ( .A(n22852), .B(n22851), .Z(n22891) );
  NANDN U23877 ( .A(n22854), .B(n22853), .Z(n22858) );
  OR U23878 ( .A(n22856), .B(n22855), .Z(n22857) );
  NAND U23879 ( .A(n22858), .B(n22857), .Z(n22871) );
  AND U23880 ( .A(b[2]), .B(a[966]), .Z(n22880) );
  AND U23881 ( .A(a[967]), .B(b[1]), .Z(n22878) );
  AND U23882 ( .A(a[965]), .B(b[3]), .Z(n22877) );
  XOR U23883 ( .A(n22878), .B(n22877), .Z(n22879) );
  XOR U23884 ( .A(n22880), .B(n22879), .Z(n22883) );
  NAND U23885 ( .A(b[0]), .B(a[968]), .Z(n22884) );
  XNOR U23886 ( .A(n22883), .B(n22884), .Z(n22885) );
  OR U23887 ( .A(n22860), .B(n22859), .Z(n22864) );
  NANDN U23888 ( .A(n22862), .B(n22861), .Z(n22863) );
  AND U23889 ( .A(n22864), .B(n22863), .Z(n22886) );
  XNOR U23890 ( .A(n22885), .B(n22886), .Z(n22872) );
  XNOR U23891 ( .A(n22871), .B(n22872), .Z(n22873) );
  NANDN U23892 ( .A(n22866), .B(n22865), .Z(n22870) );
  NAND U23893 ( .A(n22868), .B(n22867), .Z(n22869) );
  AND U23894 ( .A(n22870), .B(n22869), .Z(n22874) );
  XOR U23895 ( .A(n22873), .B(n22874), .Z(n22889) );
  XNOR U23896 ( .A(sreg[1988]), .B(n22889), .Z(n22890) );
  XOR U23897 ( .A(n22891), .B(n22890), .Z(c[1988]) );
  NANDN U23898 ( .A(n22872), .B(n22871), .Z(n22876) );
  NAND U23899 ( .A(n22874), .B(n22873), .Z(n22875) );
  NAND U23900 ( .A(n22876), .B(n22875), .Z(n22898) );
  AND U23901 ( .A(b[2]), .B(a[967]), .Z(n22904) );
  AND U23902 ( .A(a[968]), .B(b[1]), .Z(n22902) );
  AND U23903 ( .A(a[966]), .B(b[3]), .Z(n22901) );
  XOR U23904 ( .A(n22902), .B(n22901), .Z(n22903) );
  XOR U23905 ( .A(n22904), .B(n22903), .Z(n22907) );
  NAND U23906 ( .A(b[0]), .B(a[969]), .Z(n22908) );
  XOR U23907 ( .A(n22907), .B(n22908), .Z(n22910) );
  OR U23908 ( .A(n22878), .B(n22877), .Z(n22882) );
  NANDN U23909 ( .A(n22880), .B(n22879), .Z(n22881) );
  NAND U23910 ( .A(n22882), .B(n22881), .Z(n22909) );
  XNOR U23911 ( .A(n22910), .B(n22909), .Z(n22895) );
  NANDN U23912 ( .A(n22884), .B(n22883), .Z(n22888) );
  NAND U23913 ( .A(n22886), .B(n22885), .Z(n22887) );
  NAND U23914 ( .A(n22888), .B(n22887), .Z(n22896) );
  XNOR U23915 ( .A(n22895), .B(n22896), .Z(n22897) );
  XOR U23916 ( .A(n22898), .B(n22897), .Z(n22914) );
  NAND U23917 ( .A(sreg[1988]), .B(n22889), .Z(n22893) );
  OR U23918 ( .A(n22891), .B(n22890), .Z(n22892) );
  NAND U23919 ( .A(n22893), .B(n22892), .Z(n22913) );
  XNOR U23920 ( .A(sreg[1989]), .B(n22913), .Z(n22894) );
  XNOR U23921 ( .A(n22914), .B(n22894), .Z(c[1989]) );
  NANDN U23922 ( .A(n22896), .B(n22895), .Z(n22900) );
  NANDN U23923 ( .A(n22898), .B(n22897), .Z(n22899) );
  NAND U23924 ( .A(n22900), .B(n22899), .Z(n22931) );
  AND U23925 ( .A(b[2]), .B(a[968]), .Z(n22925) );
  AND U23926 ( .A(a[969]), .B(b[1]), .Z(n22923) );
  AND U23927 ( .A(a[967]), .B(b[3]), .Z(n22922) );
  XOR U23928 ( .A(n22923), .B(n22922), .Z(n22924) );
  XOR U23929 ( .A(n22925), .B(n22924), .Z(n22916) );
  NAND U23930 ( .A(b[0]), .B(a[970]), .Z(n22917) );
  XOR U23931 ( .A(n22916), .B(n22917), .Z(n22919) );
  OR U23932 ( .A(n22902), .B(n22901), .Z(n22906) );
  NANDN U23933 ( .A(n22904), .B(n22903), .Z(n22905) );
  NAND U23934 ( .A(n22906), .B(n22905), .Z(n22918) );
  XNOR U23935 ( .A(n22919), .B(n22918), .Z(n22928) );
  NANDN U23936 ( .A(n22908), .B(n22907), .Z(n22912) );
  OR U23937 ( .A(n22910), .B(n22909), .Z(n22911) );
  NAND U23938 ( .A(n22912), .B(n22911), .Z(n22929) );
  XNOR U23939 ( .A(n22928), .B(n22929), .Z(n22930) );
  XNOR U23940 ( .A(n22931), .B(n22930), .Z(n22935) );
  XOR U23941 ( .A(n22934), .B(sreg[1990]), .Z(n22915) );
  XOR U23942 ( .A(n22935), .B(n22915), .Z(c[1990]) );
  NANDN U23943 ( .A(n22917), .B(n22916), .Z(n22921) );
  OR U23944 ( .A(n22919), .B(n22918), .Z(n22920) );
  NAND U23945 ( .A(n22921), .B(n22920), .Z(n22937) );
  AND U23946 ( .A(b[2]), .B(a[969]), .Z(n22946) );
  AND U23947 ( .A(a[970]), .B(b[1]), .Z(n22944) );
  AND U23948 ( .A(a[968]), .B(b[3]), .Z(n22943) );
  XOR U23949 ( .A(n22944), .B(n22943), .Z(n22945) );
  XOR U23950 ( .A(n22946), .B(n22945), .Z(n22949) );
  NAND U23951 ( .A(b[0]), .B(a[971]), .Z(n22950) );
  XNOR U23952 ( .A(n22949), .B(n22950), .Z(n22951) );
  OR U23953 ( .A(n22923), .B(n22922), .Z(n22927) );
  NANDN U23954 ( .A(n22925), .B(n22924), .Z(n22926) );
  AND U23955 ( .A(n22927), .B(n22926), .Z(n22952) );
  XNOR U23956 ( .A(n22951), .B(n22952), .Z(n22938) );
  XNOR U23957 ( .A(n22937), .B(n22938), .Z(n22939) );
  NANDN U23958 ( .A(n22929), .B(n22928), .Z(n22933) );
  NAND U23959 ( .A(n22931), .B(n22930), .Z(n22932) );
  NAND U23960 ( .A(n22933), .B(n22932), .Z(n22940) );
  XOR U23961 ( .A(n22939), .B(n22940), .Z(n22956) );
  XOR U23962 ( .A(n22955), .B(sreg[1991]), .Z(n22936) );
  XNOR U23963 ( .A(n22956), .B(n22936), .Z(c[1991]) );
  NANDN U23964 ( .A(n22938), .B(n22937), .Z(n22942) );
  NANDN U23965 ( .A(n22940), .B(n22939), .Z(n22941) );
  NAND U23966 ( .A(n22942), .B(n22941), .Z(n22963) );
  AND U23967 ( .A(b[2]), .B(a[970]), .Z(n22969) );
  AND U23968 ( .A(a[971]), .B(b[1]), .Z(n22967) );
  AND U23969 ( .A(a[969]), .B(b[3]), .Z(n22966) );
  XOR U23970 ( .A(n22967), .B(n22966), .Z(n22968) );
  XOR U23971 ( .A(n22969), .B(n22968), .Z(n22972) );
  NAND U23972 ( .A(b[0]), .B(a[972]), .Z(n22973) );
  XOR U23973 ( .A(n22972), .B(n22973), .Z(n22975) );
  OR U23974 ( .A(n22944), .B(n22943), .Z(n22948) );
  NANDN U23975 ( .A(n22946), .B(n22945), .Z(n22947) );
  NAND U23976 ( .A(n22948), .B(n22947), .Z(n22974) );
  XNOR U23977 ( .A(n22975), .B(n22974), .Z(n22960) );
  NANDN U23978 ( .A(n22950), .B(n22949), .Z(n22954) );
  NAND U23979 ( .A(n22952), .B(n22951), .Z(n22953) );
  NAND U23980 ( .A(n22954), .B(n22953), .Z(n22961) );
  XNOR U23981 ( .A(n22960), .B(n22961), .Z(n22962) );
  XNOR U23982 ( .A(n22963), .B(n22962), .Z(n22959) );
  XOR U23983 ( .A(n22958), .B(sreg[1992]), .Z(n22957) );
  XNOR U23984 ( .A(n22959), .B(n22957), .Z(c[1992]) );
  NANDN U23985 ( .A(n22961), .B(n22960), .Z(n22965) );
  NANDN U23986 ( .A(n22963), .B(n22962), .Z(n22964) );
  NAND U23987 ( .A(n22965), .B(n22964), .Z(n22998) );
  AND U23988 ( .A(b[2]), .B(a[971]), .Z(n22992) );
  AND U23989 ( .A(a[972]), .B(b[1]), .Z(n22990) );
  AND U23990 ( .A(a[970]), .B(b[3]), .Z(n22989) );
  XOR U23991 ( .A(n22990), .B(n22989), .Z(n22991) );
  XOR U23992 ( .A(n22992), .B(n22991), .Z(n22983) );
  NAND U23993 ( .A(b[0]), .B(a[973]), .Z(n22984) );
  XOR U23994 ( .A(n22983), .B(n22984), .Z(n22986) );
  OR U23995 ( .A(n22967), .B(n22966), .Z(n22971) );
  NANDN U23996 ( .A(n22969), .B(n22968), .Z(n22970) );
  NAND U23997 ( .A(n22971), .B(n22970), .Z(n22985) );
  XNOR U23998 ( .A(n22986), .B(n22985), .Z(n22995) );
  NANDN U23999 ( .A(n22973), .B(n22972), .Z(n22977) );
  OR U24000 ( .A(n22975), .B(n22974), .Z(n22976) );
  NAND U24001 ( .A(n22977), .B(n22976), .Z(n22996) );
  XNOR U24002 ( .A(n22995), .B(n22996), .Z(n22997) );
  XNOR U24003 ( .A(n22998), .B(n22997), .Z(n22978) );
  XNOR U24004 ( .A(n22978), .B(sreg[1993]), .Z(n22980) );
  XNOR U24005 ( .A(n22979), .B(n22980), .Z(c[1993]) );
  NAND U24006 ( .A(n22978), .B(sreg[1993]), .Z(n22982) );
  NANDN U24007 ( .A(n22980), .B(n22979), .Z(n22981) );
  NAND U24008 ( .A(n22982), .B(n22981), .Z(n23020) );
  NANDN U24009 ( .A(n22984), .B(n22983), .Z(n22988) );
  OR U24010 ( .A(n22986), .B(n22985), .Z(n22987) );
  NAND U24011 ( .A(n22988), .B(n22987), .Z(n23002) );
  AND U24012 ( .A(b[2]), .B(a[972]), .Z(n23011) );
  AND U24013 ( .A(a[973]), .B(b[1]), .Z(n23009) );
  AND U24014 ( .A(a[971]), .B(b[3]), .Z(n23008) );
  XOR U24015 ( .A(n23009), .B(n23008), .Z(n23010) );
  XOR U24016 ( .A(n23011), .B(n23010), .Z(n23014) );
  NAND U24017 ( .A(b[0]), .B(a[974]), .Z(n23015) );
  XNOR U24018 ( .A(n23014), .B(n23015), .Z(n23016) );
  OR U24019 ( .A(n22990), .B(n22989), .Z(n22994) );
  NANDN U24020 ( .A(n22992), .B(n22991), .Z(n22993) );
  AND U24021 ( .A(n22994), .B(n22993), .Z(n23017) );
  XNOR U24022 ( .A(n23016), .B(n23017), .Z(n23003) );
  XNOR U24023 ( .A(n23002), .B(n23003), .Z(n23004) );
  NANDN U24024 ( .A(n22996), .B(n22995), .Z(n23000) );
  NAND U24025 ( .A(n22998), .B(n22997), .Z(n22999) );
  AND U24026 ( .A(n23000), .B(n22999), .Z(n23005) );
  XNOR U24027 ( .A(n23004), .B(n23005), .Z(n23021) );
  XOR U24028 ( .A(sreg[1994]), .B(n23021), .Z(n23001) );
  XNOR U24029 ( .A(n23020), .B(n23001), .Z(c[1994]) );
  NANDN U24030 ( .A(n23003), .B(n23002), .Z(n23007) );
  NAND U24031 ( .A(n23005), .B(n23004), .Z(n23006) );
  NAND U24032 ( .A(n23007), .B(n23006), .Z(n23028) );
  AND U24033 ( .A(b[2]), .B(a[973]), .Z(n23034) );
  AND U24034 ( .A(a[974]), .B(b[1]), .Z(n23032) );
  AND U24035 ( .A(a[972]), .B(b[3]), .Z(n23031) );
  XOR U24036 ( .A(n23032), .B(n23031), .Z(n23033) );
  XOR U24037 ( .A(n23034), .B(n23033), .Z(n23037) );
  NAND U24038 ( .A(b[0]), .B(a[975]), .Z(n23038) );
  XOR U24039 ( .A(n23037), .B(n23038), .Z(n23040) );
  OR U24040 ( .A(n23009), .B(n23008), .Z(n23013) );
  NANDN U24041 ( .A(n23011), .B(n23010), .Z(n23012) );
  NAND U24042 ( .A(n23013), .B(n23012), .Z(n23039) );
  XNOR U24043 ( .A(n23040), .B(n23039), .Z(n23025) );
  NANDN U24044 ( .A(n23015), .B(n23014), .Z(n23019) );
  NAND U24045 ( .A(n23017), .B(n23016), .Z(n23018) );
  NAND U24046 ( .A(n23019), .B(n23018), .Z(n23026) );
  XNOR U24047 ( .A(n23025), .B(n23026), .Z(n23027) );
  XNOR U24048 ( .A(n23028), .B(n23027), .Z(n23024) );
  XOR U24049 ( .A(n23023), .B(sreg[1995]), .Z(n23022) );
  XNOR U24050 ( .A(n23024), .B(n23022), .Z(c[1995]) );
  NANDN U24051 ( .A(n23026), .B(n23025), .Z(n23030) );
  NANDN U24052 ( .A(n23028), .B(n23027), .Z(n23029) );
  NAND U24053 ( .A(n23030), .B(n23029), .Z(n23063) );
  AND U24054 ( .A(b[2]), .B(a[974]), .Z(n23057) );
  AND U24055 ( .A(a[975]), .B(b[1]), .Z(n23055) );
  AND U24056 ( .A(a[973]), .B(b[3]), .Z(n23054) );
  XOR U24057 ( .A(n23055), .B(n23054), .Z(n23056) );
  XOR U24058 ( .A(n23057), .B(n23056), .Z(n23048) );
  NAND U24059 ( .A(b[0]), .B(a[976]), .Z(n23049) );
  XOR U24060 ( .A(n23048), .B(n23049), .Z(n23051) );
  OR U24061 ( .A(n23032), .B(n23031), .Z(n23036) );
  NANDN U24062 ( .A(n23034), .B(n23033), .Z(n23035) );
  NAND U24063 ( .A(n23036), .B(n23035), .Z(n23050) );
  XNOR U24064 ( .A(n23051), .B(n23050), .Z(n23060) );
  NANDN U24065 ( .A(n23038), .B(n23037), .Z(n23042) );
  OR U24066 ( .A(n23040), .B(n23039), .Z(n23041) );
  NAND U24067 ( .A(n23042), .B(n23041), .Z(n23061) );
  XNOR U24068 ( .A(n23060), .B(n23061), .Z(n23062) );
  XNOR U24069 ( .A(n23063), .B(n23062), .Z(n23043) );
  XNOR U24070 ( .A(n23043), .B(sreg[1996]), .Z(n23045) );
  XNOR U24071 ( .A(n23044), .B(n23045), .Z(c[1996]) );
  NAND U24072 ( .A(n23043), .B(sreg[1996]), .Z(n23047) );
  NANDN U24073 ( .A(n23045), .B(n23044), .Z(n23046) );
  NAND U24074 ( .A(n23047), .B(n23046), .Z(n23085) );
  NANDN U24075 ( .A(n23049), .B(n23048), .Z(n23053) );
  OR U24076 ( .A(n23051), .B(n23050), .Z(n23052) );
  NAND U24077 ( .A(n23053), .B(n23052), .Z(n23067) );
  AND U24078 ( .A(b[2]), .B(a[975]), .Z(n23076) );
  AND U24079 ( .A(a[976]), .B(b[1]), .Z(n23074) );
  AND U24080 ( .A(a[974]), .B(b[3]), .Z(n23073) );
  XOR U24081 ( .A(n23074), .B(n23073), .Z(n23075) );
  XOR U24082 ( .A(n23076), .B(n23075), .Z(n23079) );
  NAND U24083 ( .A(b[0]), .B(a[977]), .Z(n23080) );
  XNOR U24084 ( .A(n23079), .B(n23080), .Z(n23081) );
  OR U24085 ( .A(n23055), .B(n23054), .Z(n23059) );
  NANDN U24086 ( .A(n23057), .B(n23056), .Z(n23058) );
  AND U24087 ( .A(n23059), .B(n23058), .Z(n23082) );
  XNOR U24088 ( .A(n23081), .B(n23082), .Z(n23068) );
  XNOR U24089 ( .A(n23067), .B(n23068), .Z(n23069) );
  NANDN U24090 ( .A(n23061), .B(n23060), .Z(n23065) );
  NAND U24091 ( .A(n23063), .B(n23062), .Z(n23064) );
  AND U24092 ( .A(n23065), .B(n23064), .Z(n23070) );
  XNOR U24093 ( .A(n23069), .B(n23070), .Z(n23086) );
  XOR U24094 ( .A(sreg[1997]), .B(n23086), .Z(n23066) );
  XNOR U24095 ( .A(n23085), .B(n23066), .Z(c[1997]) );
  NANDN U24096 ( .A(n23068), .B(n23067), .Z(n23072) );
  NAND U24097 ( .A(n23070), .B(n23069), .Z(n23071) );
  NAND U24098 ( .A(n23072), .B(n23071), .Z(n23093) );
  AND U24099 ( .A(b[2]), .B(a[976]), .Z(n23099) );
  AND U24100 ( .A(a[977]), .B(b[1]), .Z(n23097) );
  AND U24101 ( .A(a[975]), .B(b[3]), .Z(n23096) );
  XOR U24102 ( .A(n23097), .B(n23096), .Z(n23098) );
  XOR U24103 ( .A(n23099), .B(n23098), .Z(n23102) );
  NAND U24104 ( .A(b[0]), .B(a[978]), .Z(n23103) );
  XOR U24105 ( .A(n23102), .B(n23103), .Z(n23105) );
  OR U24106 ( .A(n23074), .B(n23073), .Z(n23078) );
  NANDN U24107 ( .A(n23076), .B(n23075), .Z(n23077) );
  NAND U24108 ( .A(n23078), .B(n23077), .Z(n23104) );
  XNOR U24109 ( .A(n23105), .B(n23104), .Z(n23090) );
  NANDN U24110 ( .A(n23080), .B(n23079), .Z(n23084) );
  NAND U24111 ( .A(n23082), .B(n23081), .Z(n23083) );
  NAND U24112 ( .A(n23084), .B(n23083), .Z(n23091) );
  XNOR U24113 ( .A(n23090), .B(n23091), .Z(n23092) );
  XOR U24114 ( .A(n23093), .B(n23092), .Z(n23089) );
  XNOR U24115 ( .A(sreg[1998]), .B(n23088), .Z(n23087) );
  XNOR U24116 ( .A(n23089), .B(n23087), .Z(c[1998]) );
  NANDN U24117 ( .A(n23091), .B(n23090), .Z(n23095) );
  NANDN U24118 ( .A(n23093), .B(n23092), .Z(n23094) );
  NAND U24119 ( .A(n23095), .B(n23094), .Z(n23111) );
  AND U24120 ( .A(b[2]), .B(a[977]), .Z(n23117) );
  AND U24121 ( .A(a[978]), .B(b[1]), .Z(n23115) );
  AND U24122 ( .A(a[976]), .B(b[3]), .Z(n23114) );
  XOR U24123 ( .A(n23115), .B(n23114), .Z(n23116) );
  XOR U24124 ( .A(n23117), .B(n23116), .Z(n23120) );
  NAND U24125 ( .A(b[0]), .B(a[979]), .Z(n23121) );
  XOR U24126 ( .A(n23120), .B(n23121), .Z(n23123) );
  OR U24127 ( .A(n23097), .B(n23096), .Z(n23101) );
  NANDN U24128 ( .A(n23099), .B(n23098), .Z(n23100) );
  NAND U24129 ( .A(n23101), .B(n23100), .Z(n23122) );
  XNOR U24130 ( .A(n23123), .B(n23122), .Z(n23108) );
  NANDN U24131 ( .A(n23103), .B(n23102), .Z(n23107) );
  OR U24132 ( .A(n23105), .B(n23104), .Z(n23106) );
  NAND U24133 ( .A(n23107), .B(n23106), .Z(n23109) );
  XNOR U24134 ( .A(n23108), .B(n23109), .Z(n23110) );
  XNOR U24135 ( .A(n23111), .B(n23110), .Z(n23127) );
  XNOR U24136 ( .A(n23127), .B(sreg[1999]), .Z(n23128) );
  XOR U24137 ( .A(n23129), .B(n23128), .Z(c[1999]) );
  NANDN U24138 ( .A(n23109), .B(n23108), .Z(n23113) );
  NAND U24139 ( .A(n23111), .B(n23110), .Z(n23112) );
  AND U24140 ( .A(n23113), .B(n23112), .Z(n23134) );
  AND U24141 ( .A(b[2]), .B(a[978]), .Z(n23142) );
  AND U24142 ( .A(a[979]), .B(b[1]), .Z(n23140) );
  AND U24143 ( .A(a[977]), .B(b[3]), .Z(n23139) );
  XOR U24144 ( .A(n23140), .B(n23139), .Z(n23141) );
  XOR U24145 ( .A(n23142), .B(n23141), .Z(n23135) );
  NAND U24146 ( .A(b[0]), .B(a[980]), .Z(n23136) );
  XOR U24147 ( .A(n23135), .B(n23136), .Z(n23137) );
  OR U24148 ( .A(n23115), .B(n23114), .Z(n23119) );
  NANDN U24149 ( .A(n23117), .B(n23116), .Z(n23118) );
  AND U24150 ( .A(n23119), .B(n23118), .Z(n23138) );
  XOR U24151 ( .A(n23137), .B(n23138), .Z(n23132) );
  NANDN U24152 ( .A(n23121), .B(n23120), .Z(n23125) );
  OR U24153 ( .A(n23123), .B(n23122), .Z(n23124) );
  AND U24154 ( .A(n23125), .B(n23124), .Z(n23133) );
  XOR U24155 ( .A(n23132), .B(n23133), .Z(n23126) );
  XOR U24156 ( .A(n23134), .B(n23126), .Z(n23145) );
  XNOR U24157 ( .A(sreg[2000]), .B(n23145), .Z(n23147) );
  NAND U24158 ( .A(n23127), .B(sreg[1999]), .Z(n23131) );
  OR U24159 ( .A(n23129), .B(n23128), .Z(n23130) );
  AND U24160 ( .A(n23131), .B(n23130), .Z(n23146) );
  XOR U24161 ( .A(n23147), .B(n23146), .Z(c[2000]) );
  AND U24162 ( .A(b[2]), .B(a[979]), .Z(n23154) );
  AND U24163 ( .A(a[980]), .B(b[1]), .Z(n23152) );
  AND U24164 ( .A(a[978]), .B(b[3]), .Z(n23151) );
  XOR U24165 ( .A(n23152), .B(n23151), .Z(n23153) );
  XOR U24166 ( .A(n23154), .B(n23153), .Z(n23157) );
  NAND U24167 ( .A(b[0]), .B(a[981]), .Z(n23158) );
  XNOR U24168 ( .A(n23157), .B(n23158), .Z(n23159) );
  OR U24169 ( .A(n23140), .B(n23139), .Z(n23144) );
  NANDN U24170 ( .A(n23142), .B(n23141), .Z(n23143) );
  AND U24171 ( .A(n23144), .B(n23143), .Z(n23160) );
  XNOR U24172 ( .A(n23159), .B(n23160), .Z(n23164) );
  XNOR U24173 ( .A(n23163), .B(n23164), .Z(n23165) );
  XOR U24174 ( .A(n23166), .B(n23165), .Z(n23170) );
  NAND U24175 ( .A(sreg[2000]), .B(n23145), .Z(n23149) );
  OR U24176 ( .A(n23147), .B(n23146), .Z(n23148) );
  AND U24177 ( .A(n23149), .B(n23148), .Z(n23169) );
  XNOR U24178 ( .A(n23169), .B(sreg[2001]), .Z(n23150) );
  XNOR U24179 ( .A(n23170), .B(n23150), .Z(c[2001]) );
  AND U24180 ( .A(b[2]), .B(a[980]), .Z(n23183) );
  AND U24181 ( .A(a[981]), .B(b[1]), .Z(n23181) );
  AND U24182 ( .A(a[979]), .B(b[3]), .Z(n23180) );
  XOR U24183 ( .A(n23181), .B(n23180), .Z(n23182) );
  XOR U24184 ( .A(n23183), .B(n23182), .Z(n23186) );
  NAND U24185 ( .A(b[0]), .B(a[982]), .Z(n23187) );
  XOR U24186 ( .A(n23186), .B(n23187), .Z(n23189) );
  OR U24187 ( .A(n23152), .B(n23151), .Z(n23156) );
  NANDN U24188 ( .A(n23154), .B(n23153), .Z(n23155) );
  NAND U24189 ( .A(n23156), .B(n23155), .Z(n23188) );
  XNOR U24190 ( .A(n23189), .B(n23188), .Z(n23174) );
  NANDN U24191 ( .A(n23158), .B(n23157), .Z(n23162) );
  NAND U24192 ( .A(n23160), .B(n23159), .Z(n23161) );
  NAND U24193 ( .A(n23162), .B(n23161), .Z(n23175) );
  XNOR U24194 ( .A(n23174), .B(n23175), .Z(n23176) );
  NANDN U24195 ( .A(n23164), .B(n23163), .Z(n23168) );
  NANDN U24196 ( .A(n23166), .B(n23165), .Z(n23167) );
  NAND U24197 ( .A(n23168), .B(n23167), .Z(n23177) );
  XOR U24198 ( .A(n23176), .B(n23177), .Z(n23173) );
  XOR U24199 ( .A(sreg[2002]), .B(n23172), .Z(n23171) );
  XNOR U24200 ( .A(n23173), .B(n23171), .Z(c[2002]) );
  NANDN U24201 ( .A(n23175), .B(n23174), .Z(n23179) );
  NANDN U24202 ( .A(n23177), .B(n23176), .Z(n23178) );
  NAND U24203 ( .A(n23179), .B(n23178), .Z(n23212) );
  AND U24204 ( .A(b[2]), .B(a[981]), .Z(n23206) );
  AND U24205 ( .A(a[982]), .B(b[1]), .Z(n23204) );
  AND U24206 ( .A(a[980]), .B(b[3]), .Z(n23203) );
  XOR U24207 ( .A(n23204), .B(n23203), .Z(n23205) );
  XOR U24208 ( .A(n23206), .B(n23205), .Z(n23197) );
  NAND U24209 ( .A(b[0]), .B(a[983]), .Z(n23198) );
  XOR U24210 ( .A(n23197), .B(n23198), .Z(n23200) );
  OR U24211 ( .A(n23181), .B(n23180), .Z(n23185) );
  NANDN U24212 ( .A(n23183), .B(n23182), .Z(n23184) );
  NAND U24213 ( .A(n23185), .B(n23184), .Z(n23199) );
  XNOR U24214 ( .A(n23200), .B(n23199), .Z(n23209) );
  NANDN U24215 ( .A(n23187), .B(n23186), .Z(n23191) );
  OR U24216 ( .A(n23189), .B(n23188), .Z(n23190) );
  NAND U24217 ( .A(n23191), .B(n23190), .Z(n23210) );
  XNOR U24218 ( .A(n23209), .B(n23210), .Z(n23211) );
  XNOR U24219 ( .A(n23212), .B(n23211), .Z(n23192) );
  XNOR U24220 ( .A(n23192), .B(sreg[2003]), .Z(n23193) );
  XOR U24221 ( .A(n23194), .B(n23193), .Z(c[2003]) );
  NAND U24222 ( .A(n23192), .B(sreg[2003]), .Z(n23196) );
  OR U24223 ( .A(n23194), .B(n23193), .Z(n23195) );
  AND U24224 ( .A(n23196), .B(n23195), .Z(n23235) );
  NANDN U24225 ( .A(n23198), .B(n23197), .Z(n23202) );
  OR U24226 ( .A(n23200), .B(n23199), .Z(n23201) );
  NAND U24227 ( .A(n23202), .B(n23201), .Z(n23228) );
  AND U24228 ( .A(b[2]), .B(a[982]), .Z(n23219) );
  AND U24229 ( .A(a[983]), .B(b[1]), .Z(n23217) );
  AND U24230 ( .A(a[981]), .B(b[3]), .Z(n23216) );
  XOR U24231 ( .A(n23217), .B(n23216), .Z(n23218) );
  XOR U24232 ( .A(n23219), .B(n23218), .Z(n23222) );
  NAND U24233 ( .A(b[0]), .B(a[984]), .Z(n23223) );
  XNOR U24234 ( .A(n23222), .B(n23223), .Z(n23224) );
  OR U24235 ( .A(n23204), .B(n23203), .Z(n23208) );
  NANDN U24236 ( .A(n23206), .B(n23205), .Z(n23207) );
  AND U24237 ( .A(n23208), .B(n23207), .Z(n23225) );
  XNOR U24238 ( .A(n23224), .B(n23225), .Z(n23229) );
  XNOR U24239 ( .A(n23228), .B(n23229), .Z(n23230) );
  NANDN U24240 ( .A(n23210), .B(n23209), .Z(n23214) );
  NAND U24241 ( .A(n23212), .B(n23211), .Z(n23213) );
  AND U24242 ( .A(n23214), .B(n23213), .Z(n23231) );
  XOR U24243 ( .A(n23230), .B(n23231), .Z(n23234) );
  XNOR U24244 ( .A(sreg[2004]), .B(n23234), .Z(n23215) );
  XOR U24245 ( .A(n23235), .B(n23215), .Z(c[2004]) );
  AND U24246 ( .A(b[2]), .B(a[983]), .Z(n23248) );
  AND U24247 ( .A(a[984]), .B(b[1]), .Z(n23246) );
  AND U24248 ( .A(a[982]), .B(b[3]), .Z(n23245) );
  XOR U24249 ( .A(n23246), .B(n23245), .Z(n23247) );
  XOR U24250 ( .A(n23248), .B(n23247), .Z(n23251) );
  NAND U24251 ( .A(b[0]), .B(a[985]), .Z(n23252) );
  XOR U24252 ( .A(n23251), .B(n23252), .Z(n23254) );
  OR U24253 ( .A(n23217), .B(n23216), .Z(n23221) );
  NANDN U24254 ( .A(n23219), .B(n23218), .Z(n23220) );
  NAND U24255 ( .A(n23221), .B(n23220), .Z(n23253) );
  XNOR U24256 ( .A(n23254), .B(n23253), .Z(n23239) );
  NANDN U24257 ( .A(n23223), .B(n23222), .Z(n23227) );
  NAND U24258 ( .A(n23225), .B(n23224), .Z(n23226) );
  NAND U24259 ( .A(n23227), .B(n23226), .Z(n23240) );
  XNOR U24260 ( .A(n23239), .B(n23240), .Z(n23241) );
  NANDN U24261 ( .A(n23229), .B(n23228), .Z(n23233) );
  NAND U24262 ( .A(n23231), .B(n23230), .Z(n23232) );
  AND U24263 ( .A(n23233), .B(n23232), .Z(n23242) );
  XNOR U24264 ( .A(n23241), .B(n23242), .Z(n23238) );
  XOR U24265 ( .A(n23237), .B(sreg[2005]), .Z(n23236) );
  XOR U24266 ( .A(n23238), .B(n23236), .Z(c[2005]) );
  NANDN U24267 ( .A(n23240), .B(n23239), .Z(n23244) );
  NAND U24268 ( .A(n23242), .B(n23241), .Z(n23243) );
  NAND U24269 ( .A(n23244), .B(n23243), .Z(n23260) );
  AND U24270 ( .A(b[2]), .B(a[984]), .Z(n23266) );
  AND U24271 ( .A(a[985]), .B(b[1]), .Z(n23264) );
  AND U24272 ( .A(a[983]), .B(b[3]), .Z(n23263) );
  XOR U24273 ( .A(n23264), .B(n23263), .Z(n23265) );
  XOR U24274 ( .A(n23266), .B(n23265), .Z(n23269) );
  NAND U24275 ( .A(b[0]), .B(a[986]), .Z(n23270) );
  XOR U24276 ( .A(n23269), .B(n23270), .Z(n23272) );
  OR U24277 ( .A(n23246), .B(n23245), .Z(n23250) );
  NANDN U24278 ( .A(n23248), .B(n23247), .Z(n23249) );
  NAND U24279 ( .A(n23250), .B(n23249), .Z(n23271) );
  XNOR U24280 ( .A(n23272), .B(n23271), .Z(n23257) );
  NANDN U24281 ( .A(n23252), .B(n23251), .Z(n23256) );
  OR U24282 ( .A(n23254), .B(n23253), .Z(n23255) );
  NAND U24283 ( .A(n23256), .B(n23255), .Z(n23258) );
  XNOR U24284 ( .A(n23257), .B(n23258), .Z(n23259) );
  XNOR U24285 ( .A(n23260), .B(n23259), .Z(n23275) );
  XNOR U24286 ( .A(n23275), .B(sreg[2006]), .Z(n23277) );
  XNOR U24287 ( .A(n23276), .B(n23277), .Z(c[2006]) );
  NANDN U24288 ( .A(n23258), .B(n23257), .Z(n23262) );
  NAND U24289 ( .A(n23260), .B(n23259), .Z(n23261) );
  NAND U24290 ( .A(n23262), .B(n23261), .Z(n23286) );
  AND U24291 ( .A(b[2]), .B(a[985]), .Z(n23292) );
  AND U24292 ( .A(a[986]), .B(b[1]), .Z(n23290) );
  AND U24293 ( .A(a[984]), .B(b[3]), .Z(n23289) );
  XOR U24294 ( .A(n23290), .B(n23289), .Z(n23291) );
  XOR U24295 ( .A(n23292), .B(n23291), .Z(n23295) );
  NAND U24296 ( .A(b[0]), .B(a[987]), .Z(n23296) );
  XOR U24297 ( .A(n23295), .B(n23296), .Z(n23298) );
  OR U24298 ( .A(n23264), .B(n23263), .Z(n23268) );
  NANDN U24299 ( .A(n23266), .B(n23265), .Z(n23267) );
  NAND U24300 ( .A(n23268), .B(n23267), .Z(n23297) );
  XNOR U24301 ( .A(n23298), .B(n23297), .Z(n23283) );
  NANDN U24302 ( .A(n23270), .B(n23269), .Z(n23274) );
  OR U24303 ( .A(n23272), .B(n23271), .Z(n23273) );
  NAND U24304 ( .A(n23274), .B(n23273), .Z(n23284) );
  XNOR U24305 ( .A(n23283), .B(n23284), .Z(n23285) );
  XOR U24306 ( .A(n23286), .B(n23285), .Z(n23282) );
  NAND U24307 ( .A(n23275), .B(sreg[2006]), .Z(n23279) );
  NANDN U24308 ( .A(n23277), .B(n23276), .Z(n23278) );
  NAND U24309 ( .A(n23279), .B(n23278), .Z(n23281) );
  XNOR U24310 ( .A(sreg[2007]), .B(n23281), .Z(n23280) );
  XOR U24311 ( .A(n23282), .B(n23280), .Z(c[2007]) );
  NANDN U24312 ( .A(n23284), .B(n23283), .Z(n23288) );
  NAND U24313 ( .A(n23286), .B(n23285), .Z(n23287) );
  NAND U24314 ( .A(n23288), .B(n23287), .Z(n23304) );
  AND U24315 ( .A(b[2]), .B(a[986]), .Z(n23310) );
  AND U24316 ( .A(a[987]), .B(b[1]), .Z(n23308) );
  AND U24317 ( .A(a[985]), .B(b[3]), .Z(n23307) );
  XOR U24318 ( .A(n23308), .B(n23307), .Z(n23309) );
  XOR U24319 ( .A(n23310), .B(n23309), .Z(n23313) );
  NAND U24320 ( .A(b[0]), .B(a[988]), .Z(n23314) );
  XOR U24321 ( .A(n23313), .B(n23314), .Z(n23316) );
  OR U24322 ( .A(n23290), .B(n23289), .Z(n23294) );
  NANDN U24323 ( .A(n23292), .B(n23291), .Z(n23293) );
  NAND U24324 ( .A(n23294), .B(n23293), .Z(n23315) );
  XNOR U24325 ( .A(n23316), .B(n23315), .Z(n23301) );
  NANDN U24326 ( .A(n23296), .B(n23295), .Z(n23300) );
  OR U24327 ( .A(n23298), .B(n23297), .Z(n23299) );
  NAND U24328 ( .A(n23300), .B(n23299), .Z(n23302) );
  XNOR U24329 ( .A(n23301), .B(n23302), .Z(n23303) );
  XNOR U24330 ( .A(n23304), .B(n23303), .Z(n23319) );
  XNOR U24331 ( .A(n23319), .B(sreg[2008]), .Z(n23320) );
  XOR U24332 ( .A(n23321), .B(n23320), .Z(c[2008]) );
  NANDN U24333 ( .A(n23302), .B(n23301), .Z(n23306) );
  NAND U24334 ( .A(n23304), .B(n23303), .Z(n23305) );
  NAND U24335 ( .A(n23306), .B(n23305), .Z(n23327) );
  AND U24336 ( .A(b[2]), .B(a[987]), .Z(n23333) );
  AND U24337 ( .A(a[988]), .B(b[1]), .Z(n23331) );
  AND U24338 ( .A(a[986]), .B(b[3]), .Z(n23330) );
  XOR U24339 ( .A(n23331), .B(n23330), .Z(n23332) );
  XOR U24340 ( .A(n23333), .B(n23332), .Z(n23336) );
  NAND U24341 ( .A(b[0]), .B(a[989]), .Z(n23337) );
  XOR U24342 ( .A(n23336), .B(n23337), .Z(n23339) );
  OR U24343 ( .A(n23308), .B(n23307), .Z(n23312) );
  NANDN U24344 ( .A(n23310), .B(n23309), .Z(n23311) );
  NAND U24345 ( .A(n23312), .B(n23311), .Z(n23338) );
  XNOR U24346 ( .A(n23339), .B(n23338), .Z(n23324) );
  NANDN U24347 ( .A(n23314), .B(n23313), .Z(n23318) );
  OR U24348 ( .A(n23316), .B(n23315), .Z(n23317) );
  NAND U24349 ( .A(n23318), .B(n23317), .Z(n23325) );
  XNOR U24350 ( .A(n23324), .B(n23325), .Z(n23326) );
  XNOR U24351 ( .A(n23327), .B(n23326), .Z(n23342) );
  XNOR U24352 ( .A(n23342), .B(sreg[2009]), .Z(n23344) );
  NAND U24353 ( .A(n23319), .B(sreg[2008]), .Z(n23323) );
  OR U24354 ( .A(n23321), .B(n23320), .Z(n23322) );
  AND U24355 ( .A(n23323), .B(n23322), .Z(n23343) );
  XOR U24356 ( .A(n23344), .B(n23343), .Z(c[2009]) );
  NANDN U24357 ( .A(n23325), .B(n23324), .Z(n23329) );
  NAND U24358 ( .A(n23327), .B(n23326), .Z(n23328) );
  NAND U24359 ( .A(n23329), .B(n23328), .Z(n23353) );
  AND U24360 ( .A(b[2]), .B(a[988]), .Z(n23359) );
  AND U24361 ( .A(a[989]), .B(b[1]), .Z(n23357) );
  AND U24362 ( .A(a[987]), .B(b[3]), .Z(n23356) );
  XOR U24363 ( .A(n23357), .B(n23356), .Z(n23358) );
  XOR U24364 ( .A(n23359), .B(n23358), .Z(n23362) );
  NAND U24365 ( .A(b[0]), .B(a[990]), .Z(n23363) );
  XOR U24366 ( .A(n23362), .B(n23363), .Z(n23365) );
  OR U24367 ( .A(n23331), .B(n23330), .Z(n23335) );
  NANDN U24368 ( .A(n23333), .B(n23332), .Z(n23334) );
  NAND U24369 ( .A(n23335), .B(n23334), .Z(n23364) );
  XNOR U24370 ( .A(n23365), .B(n23364), .Z(n23350) );
  NANDN U24371 ( .A(n23337), .B(n23336), .Z(n23341) );
  OR U24372 ( .A(n23339), .B(n23338), .Z(n23340) );
  NAND U24373 ( .A(n23341), .B(n23340), .Z(n23351) );
  XNOR U24374 ( .A(n23350), .B(n23351), .Z(n23352) );
  XOR U24375 ( .A(n23353), .B(n23352), .Z(n23349) );
  NAND U24376 ( .A(n23342), .B(sreg[2009]), .Z(n23346) );
  OR U24377 ( .A(n23344), .B(n23343), .Z(n23345) );
  NAND U24378 ( .A(n23346), .B(n23345), .Z(n23348) );
  XNOR U24379 ( .A(sreg[2010]), .B(n23348), .Z(n23347) );
  XOR U24380 ( .A(n23349), .B(n23347), .Z(c[2010]) );
  NANDN U24381 ( .A(n23351), .B(n23350), .Z(n23355) );
  NAND U24382 ( .A(n23353), .B(n23352), .Z(n23354) );
  NAND U24383 ( .A(n23355), .B(n23354), .Z(n23371) );
  AND U24384 ( .A(b[2]), .B(a[989]), .Z(n23377) );
  AND U24385 ( .A(a[990]), .B(b[1]), .Z(n23375) );
  AND U24386 ( .A(a[988]), .B(b[3]), .Z(n23374) );
  XOR U24387 ( .A(n23375), .B(n23374), .Z(n23376) );
  XOR U24388 ( .A(n23377), .B(n23376), .Z(n23380) );
  NAND U24389 ( .A(b[0]), .B(a[991]), .Z(n23381) );
  XOR U24390 ( .A(n23380), .B(n23381), .Z(n23383) );
  OR U24391 ( .A(n23357), .B(n23356), .Z(n23361) );
  NANDN U24392 ( .A(n23359), .B(n23358), .Z(n23360) );
  NAND U24393 ( .A(n23361), .B(n23360), .Z(n23382) );
  XNOR U24394 ( .A(n23383), .B(n23382), .Z(n23368) );
  NANDN U24395 ( .A(n23363), .B(n23362), .Z(n23367) );
  OR U24396 ( .A(n23365), .B(n23364), .Z(n23366) );
  NAND U24397 ( .A(n23367), .B(n23366), .Z(n23369) );
  XNOR U24398 ( .A(n23368), .B(n23369), .Z(n23370) );
  XNOR U24399 ( .A(n23371), .B(n23370), .Z(n23386) );
  XNOR U24400 ( .A(n23386), .B(sreg[2011]), .Z(n23387) );
  XOR U24401 ( .A(n23388), .B(n23387), .Z(c[2011]) );
  NANDN U24402 ( .A(n23369), .B(n23368), .Z(n23373) );
  NAND U24403 ( .A(n23371), .B(n23370), .Z(n23372) );
  NAND U24404 ( .A(n23373), .B(n23372), .Z(n23397) );
  AND U24405 ( .A(b[2]), .B(a[990]), .Z(n23403) );
  AND U24406 ( .A(a[991]), .B(b[1]), .Z(n23401) );
  AND U24407 ( .A(a[989]), .B(b[3]), .Z(n23400) );
  XOR U24408 ( .A(n23401), .B(n23400), .Z(n23402) );
  XOR U24409 ( .A(n23403), .B(n23402), .Z(n23406) );
  NAND U24410 ( .A(b[0]), .B(a[992]), .Z(n23407) );
  XOR U24411 ( .A(n23406), .B(n23407), .Z(n23409) );
  OR U24412 ( .A(n23375), .B(n23374), .Z(n23379) );
  NANDN U24413 ( .A(n23377), .B(n23376), .Z(n23378) );
  NAND U24414 ( .A(n23379), .B(n23378), .Z(n23408) );
  XNOR U24415 ( .A(n23409), .B(n23408), .Z(n23394) );
  NANDN U24416 ( .A(n23381), .B(n23380), .Z(n23385) );
  OR U24417 ( .A(n23383), .B(n23382), .Z(n23384) );
  NAND U24418 ( .A(n23385), .B(n23384), .Z(n23395) );
  XNOR U24419 ( .A(n23394), .B(n23395), .Z(n23396) );
  XOR U24420 ( .A(n23397), .B(n23396), .Z(n23393) );
  NAND U24421 ( .A(n23386), .B(sreg[2011]), .Z(n23390) );
  OR U24422 ( .A(n23388), .B(n23387), .Z(n23389) );
  NAND U24423 ( .A(n23390), .B(n23389), .Z(n23392) );
  XNOR U24424 ( .A(sreg[2012]), .B(n23392), .Z(n23391) );
  XOR U24425 ( .A(n23393), .B(n23391), .Z(c[2012]) );
  NANDN U24426 ( .A(n23395), .B(n23394), .Z(n23399) );
  NAND U24427 ( .A(n23397), .B(n23396), .Z(n23398) );
  NAND U24428 ( .A(n23399), .B(n23398), .Z(n23420) );
  AND U24429 ( .A(b[2]), .B(a[991]), .Z(n23426) );
  AND U24430 ( .A(a[992]), .B(b[1]), .Z(n23424) );
  AND U24431 ( .A(a[990]), .B(b[3]), .Z(n23423) );
  XOR U24432 ( .A(n23424), .B(n23423), .Z(n23425) );
  XOR U24433 ( .A(n23426), .B(n23425), .Z(n23429) );
  NAND U24434 ( .A(b[0]), .B(a[993]), .Z(n23430) );
  XOR U24435 ( .A(n23429), .B(n23430), .Z(n23432) );
  OR U24436 ( .A(n23401), .B(n23400), .Z(n23405) );
  NANDN U24437 ( .A(n23403), .B(n23402), .Z(n23404) );
  NAND U24438 ( .A(n23405), .B(n23404), .Z(n23431) );
  XNOR U24439 ( .A(n23432), .B(n23431), .Z(n23417) );
  NANDN U24440 ( .A(n23407), .B(n23406), .Z(n23411) );
  OR U24441 ( .A(n23409), .B(n23408), .Z(n23410) );
  NAND U24442 ( .A(n23411), .B(n23410), .Z(n23418) );
  XNOR U24443 ( .A(n23417), .B(n23418), .Z(n23419) );
  XNOR U24444 ( .A(n23420), .B(n23419), .Z(n23412) );
  XOR U24445 ( .A(sreg[2013]), .B(n23412), .Z(n23414) );
  XNOR U24446 ( .A(n23413), .B(n23414), .Z(c[2013]) );
  OR U24447 ( .A(n23412), .B(sreg[2013]), .Z(n23416) );
  NAND U24448 ( .A(n23414), .B(n23413), .Z(n23415) );
  AND U24449 ( .A(n23416), .B(n23415), .Z(n23436) );
  NANDN U24450 ( .A(n23418), .B(n23417), .Z(n23422) );
  NAND U24451 ( .A(n23420), .B(n23419), .Z(n23421) );
  NAND U24452 ( .A(n23422), .B(n23421), .Z(n23441) );
  AND U24453 ( .A(b[2]), .B(a[992]), .Z(n23447) );
  AND U24454 ( .A(a[993]), .B(b[1]), .Z(n23445) );
  AND U24455 ( .A(a[991]), .B(b[3]), .Z(n23444) );
  XOR U24456 ( .A(n23445), .B(n23444), .Z(n23446) );
  XOR U24457 ( .A(n23447), .B(n23446), .Z(n23450) );
  NAND U24458 ( .A(b[0]), .B(a[994]), .Z(n23451) );
  XOR U24459 ( .A(n23450), .B(n23451), .Z(n23453) );
  OR U24460 ( .A(n23424), .B(n23423), .Z(n23428) );
  NANDN U24461 ( .A(n23426), .B(n23425), .Z(n23427) );
  NAND U24462 ( .A(n23428), .B(n23427), .Z(n23452) );
  XNOR U24463 ( .A(n23453), .B(n23452), .Z(n23438) );
  NANDN U24464 ( .A(n23430), .B(n23429), .Z(n23434) );
  OR U24465 ( .A(n23432), .B(n23431), .Z(n23433) );
  NAND U24466 ( .A(n23434), .B(n23433), .Z(n23439) );
  XNOR U24467 ( .A(n23438), .B(n23439), .Z(n23440) );
  XNOR U24468 ( .A(n23441), .B(n23440), .Z(n23437) );
  XOR U24469 ( .A(sreg[2014]), .B(n23437), .Z(n23435) );
  XOR U24470 ( .A(n23436), .B(n23435), .Z(c[2014]) );
  NANDN U24471 ( .A(n23439), .B(n23438), .Z(n23443) );
  NAND U24472 ( .A(n23441), .B(n23440), .Z(n23442) );
  NAND U24473 ( .A(n23443), .B(n23442), .Z(n23459) );
  AND U24474 ( .A(b[2]), .B(a[993]), .Z(n23465) );
  AND U24475 ( .A(a[994]), .B(b[1]), .Z(n23463) );
  AND U24476 ( .A(a[992]), .B(b[3]), .Z(n23462) );
  XOR U24477 ( .A(n23463), .B(n23462), .Z(n23464) );
  XOR U24478 ( .A(n23465), .B(n23464), .Z(n23468) );
  NAND U24479 ( .A(b[0]), .B(a[995]), .Z(n23469) );
  XOR U24480 ( .A(n23468), .B(n23469), .Z(n23471) );
  OR U24481 ( .A(n23445), .B(n23444), .Z(n23449) );
  NANDN U24482 ( .A(n23447), .B(n23446), .Z(n23448) );
  NAND U24483 ( .A(n23449), .B(n23448), .Z(n23470) );
  XNOR U24484 ( .A(n23471), .B(n23470), .Z(n23456) );
  NANDN U24485 ( .A(n23451), .B(n23450), .Z(n23455) );
  OR U24486 ( .A(n23453), .B(n23452), .Z(n23454) );
  NAND U24487 ( .A(n23455), .B(n23454), .Z(n23457) );
  XNOR U24488 ( .A(n23456), .B(n23457), .Z(n23458) );
  XNOR U24489 ( .A(n23459), .B(n23458), .Z(n23474) );
  XNOR U24490 ( .A(n23474), .B(sreg[2015]), .Z(n23476) );
  XNOR U24491 ( .A(n23475), .B(n23476), .Z(c[2015]) );
  NANDN U24492 ( .A(n23457), .B(n23456), .Z(n23461) );
  NAND U24493 ( .A(n23459), .B(n23458), .Z(n23460) );
  NAND U24494 ( .A(n23461), .B(n23460), .Z(n23487) );
  AND U24495 ( .A(b[2]), .B(a[994]), .Z(n23493) );
  AND U24496 ( .A(a[995]), .B(b[1]), .Z(n23491) );
  AND U24497 ( .A(a[993]), .B(b[3]), .Z(n23490) );
  XOR U24498 ( .A(n23491), .B(n23490), .Z(n23492) );
  XOR U24499 ( .A(n23493), .B(n23492), .Z(n23496) );
  NAND U24500 ( .A(b[0]), .B(a[996]), .Z(n23497) );
  XOR U24501 ( .A(n23496), .B(n23497), .Z(n23499) );
  OR U24502 ( .A(n23463), .B(n23462), .Z(n23467) );
  NANDN U24503 ( .A(n23465), .B(n23464), .Z(n23466) );
  NAND U24504 ( .A(n23467), .B(n23466), .Z(n23498) );
  XNOR U24505 ( .A(n23499), .B(n23498), .Z(n23484) );
  NANDN U24506 ( .A(n23469), .B(n23468), .Z(n23473) );
  OR U24507 ( .A(n23471), .B(n23470), .Z(n23472) );
  NAND U24508 ( .A(n23473), .B(n23472), .Z(n23485) );
  XNOR U24509 ( .A(n23484), .B(n23485), .Z(n23486) );
  XNOR U24510 ( .A(n23487), .B(n23486), .Z(n23479) );
  XOR U24511 ( .A(sreg[2016]), .B(n23479), .Z(n23480) );
  NAND U24512 ( .A(n23474), .B(sreg[2015]), .Z(n23478) );
  NANDN U24513 ( .A(n23476), .B(n23475), .Z(n23477) );
  NAND U24514 ( .A(n23478), .B(n23477), .Z(n23481) );
  XOR U24515 ( .A(n23480), .B(n23481), .Z(c[2016]) );
  OR U24516 ( .A(n23479), .B(sreg[2016]), .Z(n23483) );
  NANDN U24517 ( .A(n23481), .B(n23480), .Z(n23482) );
  AND U24518 ( .A(n23483), .B(n23482), .Z(n23521) );
  NANDN U24519 ( .A(n23485), .B(n23484), .Z(n23489) );
  NAND U24520 ( .A(n23487), .B(n23486), .Z(n23488) );
  NAND U24521 ( .A(n23489), .B(n23488), .Z(n23506) );
  AND U24522 ( .A(b[2]), .B(a[995]), .Z(n23512) );
  AND U24523 ( .A(a[996]), .B(b[1]), .Z(n23510) );
  AND U24524 ( .A(a[994]), .B(b[3]), .Z(n23509) );
  XOR U24525 ( .A(n23510), .B(n23509), .Z(n23511) );
  XOR U24526 ( .A(n23512), .B(n23511), .Z(n23515) );
  NAND U24527 ( .A(b[0]), .B(a[997]), .Z(n23516) );
  XOR U24528 ( .A(n23515), .B(n23516), .Z(n23518) );
  OR U24529 ( .A(n23491), .B(n23490), .Z(n23495) );
  NANDN U24530 ( .A(n23493), .B(n23492), .Z(n23494) );
  NAND U24531 ( .A(n23495), .B(n23494), .Z(n23517) );
  XNOR U24532 ( .A(n23518), .B(n23517), .Z(n23503) );
  NANDN U24533 ( .A(n23497), .B(n23496), .Z(n23501) );
  OR U24534 ( .A(n23499), .B(n23498), .Z(n23500) );
  NAND U24535 ( .A(n23501), .B(n23500), .Z(n23504) );
  XNOR U24536 ( .A(n23503), .B(n23504), .Z(n23505) );
  XNOR U24537 ( .A(n23506), .B(n23505), .Z(n23522) );
  XOR U24538 ( .A(sreg[2017]), .B(n23522), .Z(n23502) );
  XOR U24539 ( .A(n23521), .B(n23502), .Z(c[2017]) );
  NANDN U24540 ( .A(n23504), .B(n23503), .Z(n23508) );
  NAND U24541 ( .A(n23506), .B(n23505), .Z(n23507) );
  NAND U24542 ( .A(n23508), .B(n23507), .Z(n23529) );
  AND U24543 ( .A(b[2]), .B(a[996]), .Z(n23535) );
  AND U24544 ( .A(a[997]), .B(b[1]), .Z(n23533) );
  AND U24545 ( .A(a[995]), .B(b[3]), .Z(n23532) );
  XOR U24546 ( .A(n23533), .B(n23532), .Z(n23534) );
  XOR U24547 ( .A(n23535), .B(n23534), .Z(n23538) );
  NAND U24548 ( .A(b[0]), .B(a[998]), .Z(n23539) );
  XOR U24549 ( .A(n23538), .B(n23539), .Z(n23541) );
  OR U24550 ( .A(n23510), .B(n23509), .Z(n23514) );
  NANDN U24551 ( .A(n23512), .B(n23511), .Z(n23513) );
  NAND U24552 ( .A(n23514), .B(n23513), .Z(n23540) );
  XNOR U24553 ( .A(n23541), .B(n23540), .Z(n23526) );
  NANDN U24554 ( .A(n23516), .B(n23515), .Z(n23520) );
  OR U24555 ( .A(n23518), .B(n23517), .Z(n23519) );
  NAND U24556 ( .A(n23520), .B(n23519), .Z(n23527) );
  XNOR U24557 ( .A(n23526), .B(n23527), .Z(n23528) );
  XNOR U24558 ( .A(n23529), .B(n23528), .Z(n23525) );
  XOR U24559 ( .A(n23524), .B(sreg[2018]), .Z(n23523) );
  XOR U24560 ( .A(n23525), .B(n23523), .Z(c[2018]) );
  NANDN U24561 ( .A(n23527), .B(n23526), .Z(n23531) );
  NAND U24562 ( .A(n23529), .B(n23528), .Z(n23530) );
  NAND U24563 ( .A(n23531), .B(n23530), .Z(n23547) );
  AND U24564 ( .A(b[2]), .B(a[997]), .Z(n23553) );
  AND U24565 ( .A(a[998]), .B(b[1]), .Z(n23551) );
  AND U24566 ( .A(a[996]), .B(b[3]), .Z(n23550) );
  XOR U24567 ( .A(n23551), .B(n23550), .Z(n23552) );
  XOR U24568 ( .A(n23553), .B(n23552), .Z(n23556) );
  NAND U24569 ( .A(b[0]), .B(a[999]), .Z(n23557) );
  XOR U24570 ( .A(n23556), .B(n23557), .Z(n23559) );
  OR U24571 ( .A(n23533), .B(n23532), .Z(n23537) );
  NANDN U24572 ( .A(n23535), .B(n23534), .Z(n23536) );
  NAND U24573 ( .A(n23537), .B(n23536), .Z(n23558) );
  XNOR U24574 ( .A(n23559), .B(n23558), .Z(n23544) );
  NANDN U24575 ( .A(n23539), .B(n23538), .Z(n23543) );
  OR U24576 ( .A(n23541), .B(n23540), .Z(n23542) );
  NAND U24577 ( .A(n23543), .B(n23542), .Z(n23545) );
  XNOR U24578 ( .A(n23544), .B(n23545), .Z(n23546) );
  XNOR U24579 ( .A(n23547), .B(n23546), .Z(n23562) );
  XNOR U24580 ( .A(n23562), .B(sreg[2019]), .Z(n23564) );
  XNOR U24581 ( .A(n23563), .B(n23564), .Z(c[2019]) );
  NANDN U24582 ( .A(n23545), .B(n23544), .Z(n23549) );
  NAND U24583 ( .A(n23547), .B(n23546), .Z(n23548) );
  NAND U24584 ( .A(n23549), .B(n23548), .Z(n23571) );
  AND U24585 ( .A(b[2]), .B(a[998]), .Z(n23577) );
  AND U24586 ( .A(a[999]), .B(b[1]), .Z(n23575) );
  AND U24587 ( .A(a[997]), .B(b[3]), .Z(n23574) );
  XOR U24588 ( .A(n23575), .B(n23574), .Z(n23576) );
  XOR U24589 ( .A(n23577), .B(n23576), .Z(n23580) );
  NAND U24590 ( .A(b[0]), .B(a[1000]), .Z(n23581) );
  XOR U24591 ( .A(n23580), .B(n23581), .Z(n23583) );
  OR U24592 ( .A(n23551), .B(n23550), .Z(n23555) );
  NANDN U24593 ( .A(n23553), .B(n23552), .Z(n23554) );
  NAND U24594 ( .A(n23555), .B(n23554), .Z(n23582) );
  XNOR U24595 ( .A(n23583), .B(n23582), .Z(n23568) );
  NANDN U24596 ( .A(n23557), .B(n23556), .Z(n23561) );
  OR U24597 ( .A(n23559), .B(n23558), .Z(n23560) );
  NAND U24598 ( .A(n23561), .B(n23560), .Z(n23569) );
  XNOR U24599 ( .A(n23568), .B(n23569), .Z(n23570) );
  XNOR U24600 ( .A(n23571), .B(n23570), .Z(n23587) );
  NAND U24601 ( .A(n23562), .B(sreg[2019]), .Z(n23566) );
  NANDN U24602 ( .A(n23564), .B(n23563), .Z(n23565) );
  AND U24603 ( .A(n23566), .B(n23565), .Z(n23586) );
  XNOR U24604 ( .A(n23586), .B(sreg[2020]), .Z(n23567) );
  XOR U24605 ( .A(n23587), .B(n23567), .Z(c[2020]) );
  NANDN U24606 ( .A(n23569), .B(n23568), .Z(n23573) );
  NAND U24607 ( .A(n23571), .B(n23570), .Z(n23572) );
  NAND U24608 ( .A(n23573), .B(n23572), .Z(n23592) );
  AND U24609 ( .A(b[2]), .B(a[999]), .Z(n23598) );
  AND U24610 ( .A(a[1000]), .B(b[1]), .Z(n23596) );
  AND U24611 ( .A(a[998]), .B(b[3]), .Z(n23595) );
  XOR U24612 ( .A(n23596), .B(n23595), .Z(n23597) );
  XOR U24613 ( .A(n23598), .B(n23597), .Z(n23601) );
  NAND U24614 ( .A(b[0]), .B(a[1001]), .Z(n23602) );
  XOR U24615 ( .A(n23601), .B(n23602), .Z(n23604) );
  OR U24616 ( .A(n23575), .B(n23574), .Z(n23579) );
  NANDN U24617 ( .A(n23577), .B(n23576), .Z(n23578) );
  NAND U24618 ( .A(n23579), .B(n23578), .Z(n23603) );
  XNOR U24619 ( .A(n23604), .B(n23603), .Z(n23589) );
  NANDN U24620 ( .A(n23581), .B(n23580), .Z(n23585) );
  OR U24621 ( .A(n23583), .B(n23582), .Z(n23584) );
  NAND U24622 ( .A(n23585), .B(n23584), .Z(n23590) );
  XNOR U24623 ( .A(n23589), .B(n23590), .Z(n23591) );
  XOR U24624 ( .A(n23592), .B(n23591), .Z(n23608) );
  XOR U24625 ( .A(sreg[2021]), .B(n23607), .Z(n23588) );
  XOR U24626 ( .A(n23608), .B(n23588), .Z(c[2021]) );
  NANDN U24627 ( .A(n23590), .B(n23589), .Z(n23594) );
  NAND U24628 ( .A(n23592), .B(n23591), .Z(n23593) );
  NAND U24629 ( .A(n23594), .B(n23593), .Z(n23615) );
  AND U24630 ( .A(b[2]), .B(a[1000]), .Z(n23621) );
  AND U24631 ( .A(a[1001]), .B(b[1]), .Z(n23619) );
  AND U24632 ( .A(a[999]), .B(b[3]), .Z(n23618) );
  XOR U24633 ( .A(n23619), .B(n23618), .Z(n23620) );
  XOR U24634 ( .A(n23621), .B(n23620), .Z(n23624) );
  NAND U24635 ( .A(b[0]), .B(a[1002]), .Z(n23625) );
  XOR U24636 ( .A(n23624), .B(n23625), .Z(n23627) );
  OR U24637 ( .A(n23596), .B(n23595), .Z(n23600) );
  NANDN U24638 ( .A(n23598), .B(n23597), .Z(n23599) );
  NAND U24639 ( .A(n23600), .B(n23599), .Z(n23626) );
  XNOR U24640 ( .A(n23627), .B(n23626), .Z(n23612) );
  NANDN U24641 ( .A(n23602), .B(n23601), .Z(n23606) );
  OR U24642 ( .A(n23604), .B(n23603), .Z(n23605) );
  NAND U24643 ( .A(n23606), .B(n23605), .Z(n23613) );
  XNOR U24644 ( .A(n23612), .B(n23613), .Z(n23614) );
  XOR U24645 ( .A(n23615), .B(n23614), .Z(n23611) );
  XNOR U24646 ( .A(sreg[2022]), .B(n23610), .Z(n23609) );
  XOR U24647 ( .A(n23611), .B(n23609), .Z(c[2022]) );
  NANDN U24648 ( .A(n23613), .B(n23612), .Z(n23617) );
  NAND U24649 ( .A(n23615), .B(n23614), .Z(n23616) );
  NAND U24650 ( .A(n23617), .B(n23616), .Z(n23633) );
  AND U24651 ( .A(b[2]), .B(a[1001]), .Z(n23639) );
  AND U24652 ( .A(a[1002]), .B(b[1]), .Z(n23637) );
  AND U24653 ( .A(a[1000]), .B(b[3]), .Z(n23636) );
  XOR U24654 ( .A(n23637), .B(n23636), .Z(n23638) );
  XOR U24655 ( .A(n23639), .B(n23638), .Z(n23642) );
  NAND U24656 ( .A(b[0]), .B(a[1003]), .Z(n23643) );
  XOR U24657 ( .A(n23642), .B(n23643), .Z(n23645) );
  OR U24658 ( .A(n23619), .B(n23618), .Z(n23623) );
  NANDN U24659 ( .A(n23621), .B(n23620), .Z(n23622) );
  NAND U24660 ( .A(n23623), .B(n23622), .Z(n23644) );
  XNOR U24661 ( .A(n23645), .B(n23644), .Z(n23630) );
  NANDN U24662 ( .A(n23625), .B(n23624), .Z(n23629) );
  OR U24663 ( .A(n23627), .B(n23626), .Z(n23628) );
  NAND U24664 ( .A(n23629), .B(n23628), .Z(n23631) );
  XNOR U24665 ( .A(n23630), .B(n23631), .Z(n23632) );
  XNOR U24666 ( .A(n23633), .B(n23632), .Z(n23648) );
  XNOR U24667 ( .A(n23648), .B(sreg[2023]), .Z(n23649) );
  XOR U24668 ( .A(n23650), .B(n23649), .Z(c[2023]) );
  NANDN U24669 ( .A(n23631), .B(n23630), .Z(n23635) );
  NAND U24670 ( .A(n23633), .B(n23632), .Z(n23634) );
  NAND U24671 ( .A(n23635), .B(n23634), .Z(n23657) );
  AND U24672 ( .A(b[2]), .B(a[1002]), .Z(n23663) );
  AND U24673 ( .A(a[1003]), .B(b[1]), .Z(n23661) );
  AND U24674 ( .A(a[1001]), .B(b[3]), .Z(n23660) );
  XOR U24675 ( .A(n23661), .B(n23660), .Z(n23662) );
  XOR U24676 ( .A(n23663), .B(n23662), .Z(n23666) );
  NAND U24677 ( .A(b[0]), .B(a[1004]), .Z(n23667) );
  XOR U24678 ( .A(n23666), .B(n23667), .Z(n23669) );
  OR U24679 ( .A(n23637), .B(n23636), .Z(n23641) );
  NANDN U24680 ( .A(n23639), .B(n23638), .Z(n23640) );
  NAND U24681 ( .A(n23641), .B(n23640), .Z(n23668) );
  XNOR U24682 ( .A(n23669), .B(n23668), .Z(n23654) );
  NANDN U24683 ( .A(n23643), .B(n23642), .Z(n23647) );
  OR U24684 ( .A(n23645), .B(n23644), .Z(n23646) );
  NAND U24685 ( .A(n23647), .B(n23646), .Z(n23655) );
  XNOR U24686 ( .A(n23654), .B(n23655), .Z(n23656) );
  XOR U24687 ( .A(n23657), .B(n23656), .Z(n23673) );
  NAND U24688 ( .A(n23648), .B(sreg[2023]), .Z(n23652) );
  OR U24689 ( .A(n23650), .B(n23649), .Z(n23651) );
  NAND U24690 ( .A(n23652), .B(n23651), .Z(n23672) );
  XNOR U24691 ( .A(sreg[2024]), .B(n23672), .Z(n23653) );
  XOR U24692 ( .A(n23673), .B(n23653), .Z(c[2024]) );
  NANDN U24693 ( .A(n23655), .B(n23654), .Z(n23659) );
  NAND U24694 ( .A(n23657), .B(n23656), .Z(n23658) );
  NAND U24695 ( .A(n23659), .B(n23658), .Z(n23678) );
  AND U24696 ( .A(b[2]), .B(a[1003]), .Z(n23684) );
  AND U24697 ( .A(a[1004]), .B(b[1]), .Z(n23682) );
  AND U24698 ( .A(a[1002]), .B(b[3]), .Z(n23681) );
  XOR U24699 ( .A(n23682), .B(n23681), .Z(n23683) );
  XOR U24700 ( .A(n23684), .B(n23683), .Z(n23687) );
  NAND U24701 ( .A(b[0]), .B(a[1005]), .Z(n23688) );
  XOR U24702 ( .A(n23687), .B(n23688), .Z(n23690) );
  OR U24703 ( .A(n23661), .B(n23660), .Z(n23665) );
  NANDN U24704 ( .A(n23663), .B(n23662), .Z(n23664) );
  NAND U24705 ( .A(n23665), .B(n23664), .Z(n23689) );
  XNOR U24706 ( .A(n23690), .B(n23689), .Z(n23675) );
  NANDN U24707 ( .A(n23667), .B(n23666), .Z(n23671) );
  OR U24708 ( .A(n23669), .B(n23668), .Z(n23670) );
  NAND U24709 ( .A(n23671), .B(n23670), .Z(n23676) );
  XNOR U24710 ( .A(n23675), .B(n23676), .Z(n23677) );
  XOR U24711 ( .A(n23678), .B(n23677), .Z(n23694) );
  XNOR U24712 ( .A(sreg[2025]), .B(n23693), .Z(n23674) );
  XOR U24713 ( .A(n23694), .B(n23674), .Z(c[2025]) );
  NANDN U24714 ( .A(n23676), .B(n23675), .Z(n23680) );
  NAND U24715 ( .A(n23678), .B(n23677), .Z(n23679) );
  NAND U24716 ( .A(n23680), .B(n23679), .Z(n23701) );
  AND U24717 ( .A(b[2]), .B(a[1004]), .Z(n23707) );
  AND U24718 ( .A(a[1005]), .B(b[1]), .Z(n23705) );
  AND U24719 ( .A(a[1003]), .B(b[3]), .Z(n23704) );
  XOR U24720 ( .A(n23705), .B(n23704), .Z(n23706) );
  XOR U24721 ( .A(n23707), .B(n23706), .Z(n23710) );
  NAND U24722 ( .A(b[0]), .B(a[1006]), .Z(n23711) );
  XOR U24723 ( .A(n23710), .B(n23711), .Z(n23713) );
  OR U24724 ( .A(n23682), .B(n23681), .Z(n23686) );
  NANDN U24725 ( .A(n23684), .B(n23683), .Z(n23685) );
  NAND U24726 ( .A(n23686), .B(n23685), .Z(n23712) );
  XNOR U24727 ( .A(n23713), .B(n23712), .Z(n23698) );
  NANDN U24728 ( .A(n23688), .B(n23687), .Z(n23692) );
  OR U24729 ( .A(n23690), .B(n23689), .Z(n23691) );
  NAND U24730 ( .A(n23692), .B(n23691), .Z(n23699) );
  XNOR U24731 ( .A(n23698), .B(n23699), .Z(n23700) );
  XOR U24732 ( .A(n23701), .B(n23700), .Z(n23697) );
  XNOR U24733 ( .A(sreg[2026]), .B(n23696), .Z(n23695) );
  XOR U24734 ( .A(n23697), .B(n23695), .Z(c[2026]) );
  NANDN U24735 ( .A(n23699), .B(n23698), .Z(n23703) );
  NAND U24736 ( .A(n23701), .B(n23700), .Z(n23702) );
  NAND U24737 ( .A(n23703), .B(n23702), .Z(n23719) );
  AND U24738 ( .A(b[2]), .B(a[1005]), .Z(n23725) );
  AND U24739 ( .A(a[1006]), .B(b[1]), .Z(n23723) );
  AND U24740 ( .A(a[1004]), .B(b[3]), .Z(n23722) );
  XOR U24741 ( .A(n23723), .B(n23722), .Z(n23724) );
  XOR U24742 ( .A(n23725), .B(n23724), .Z(n23728) );
  NAND U24743 ( .A(b[0]), .B(a[1007]), .Z(n23729) );
  XOR U24744 ( .A(n23728), .B(n23729), .Z(n23731) );
  OR U24745 ( .A(n23705), .B(n23704), .Z(n23709) );
  NANDN U24746 ( .A(n23707), .B(n23706), .Z(n23708) );
  NAND U24747 ( .A(n23709), .B(n23708), .Z(n23730) );
  XNOR U24748 ( .A(n23731), .B(n23730), .Z(n23716) );
  NANDN U24749 ( .A(n23711), .B(n23710), .Z(n23715) );
  OR U24750 ( .A(n23713), .B(n23712), .Z(n23714) );
  NAND U24751 ( .A(n23715), .B(n23714), .Z(n23717) );
  XNOR U24752 ( .A(n23716), .B(n23717), .Z(n23718) );
  XNOR U24753 ( .A(n23719), .B(n23718), .Z(n23734) );
  XNOR U24754 ( .A(n23734), .B(sreg[2027]), .Z(n23735) );
  XOR U24755 ( .A(n23736), .B(n23735), .Z(c[2027]) );
  NANDN U24756 ( .A(n23717), .B(n23716), .Z(n23721) );
  NAND U24757 ( .A(n23719), .B(n23718), .Z(n23720) );
  NAND U24758 ( .A(n23721), .B(n23720), .Z(n23742) );
  AND U24759 ( .A(b[2]), .B(a[1006]), .Z(n23748) );
  AND U24760 ( .A(a[1007]), .B(b[1]), .Z(n23746) );
  AND U24761 ( .A(a[1005]), .B(b[3]), .Z(n23745) );
  XOR U24762 ( .A(n23746), .B(n23745), .Z(n23747) );
  XOR U24763 ( .A(n23748), .B(n23747), .Z(n23751) );
  NAND U24764 ( .A(b[0]), .B(a[1008]), .Z(n23752) );
  XOR U24765 ( .A(n23751), .B(n23752), .Z(n23754) );
  OR U24766 ( .A(n23723), .B(n23722), .Z(n23727) );
  NANDN U24767 ( .A(n23725), .B(n23724), .Z(n23726) );
  NAND U24768 ( .A(n23727), .B(n23726), .Z(n23753) );
  XNOR U24769 ( .A(n23754), .B(n23753), .Z(n23739) );
  NANDN U24770 ( .A(n23729), .B(n23728), .Z(n23733) );
  OR U24771 ( .A(n23731), .B(n23730), .Z(n23732) );
  NAND U24772 ( .A(n23733), .B(n23732), .Z(n23740) );
  XNOR U24773 ( .A(n23739), .B(n23740), .Z(n23741) );
  XNOR U24774 ( .A(n23742), .B(n23741), .Z(n23757) );
  XOR U24775 ( .A(sreg[2028]), .B(n23757), .Z(n23758) );
  NAND U24776 ( .A(n23734), .B(sreg[2027]), .Z(n23738) );
  OR U24777 ( .A(n23736), .B(n23735), .Z(n23737) );
  NAND U24778 ( .A(n23738), .B(n23737), .Z(n23759) );
  XOR U24779 ( .A(n23758), .B(n23759), .Z(c[2028]) );
  NANDN U24780 ( .A(n23740), .B(n23739), .Z(n23744) );
  NAND U24781 ( .A(n23742), .B(n23741), .Z(n23743) );
  NAND U24782 ( .A(n23744), .B(n23743), .Z(n23768) );
  AND U24783 ( .A(b[2]), .B(a[1007]), .Z(n23774) );
  AND U24784 ( .A(a[1008]), .B(b[1]), .Z(n23772) );
  AND U24785 ( .A(a[1006]), .B(b[3]), .Z(n23771) );
  XOR U24786 ( .A(n23772), .B(n23771), .Z(n23773) );
  XOR U24787 ( .A(n23774), .B(n23773), .Z(n23777) );
  NAND U24788 ( .A(b[0]), .B(a[1009]), .Z(n23778) );
  XOR U24789 ( .A(n23777), .B(n23778), .Z(n23780) );
  OR U24790 ( .A(n23746), .B(n23745), .Z(n23750) );
  NANDN U24791 ( .A(n23748), .B(n23747), .Z(n23749) );
  NAND U24792 ( .A(n23750), .B(n23749), .Z(n23779) );
  XNOR U24793 ( .A(n23780), .B(n23779), .Z(n23765) );
  NANDN U24794 ( .A(n23752), .B(n23751), .Z(n23756) );
  OR U24795 ( .A(n23754), .B(n23753), .Z(n23755) );
  NAND U24796 ( .A(n23756), .B(n23755), .Z(n23766) );
  XNOR U24797 ( .A(n23765), .B(n23766), .Z(n23767) );
  XOR U24798 ( .A(n23768), .B(n23767), .Z(n23764) );
  OR U24799 ( .A(n23757), .B(sreg[2028]), .Z(n23761) );
  NANDN U24800 ( .A(n23759), .B(n23758), .Z(n23760) );
  AND U24801 ( .A(n23761), .B(n23760), .Z(n23763) );
  XNOR U24802 ( .A(sreg[2029]), .B(n23763), .Z(n23762) );
  XOR U24803 ( .A(n23764), .B(n23762), .Z(c[2029]) );
  NANDN U24804 ( .A(n23766), .B(n23765), .Z(n23770) );
  NAND U24805 ( .A(n23768), .B(n23767), .Z(n23769) );
  NAND U24806 ( .A(n23770), .B(n23769), .Z(n23786) );
  AND U24807 ( .A(b[2]), .B(a[1008]), .Z(n23792) );
  AND U24808 ( .A(a[1009]), .B(b[1]), .Z(n23790) );
  AND U24809 ( .A(a[1007]), .B(b[3]), .Z(n23789) );
  XOR U24810 ( .A(n23790), .B(n23789), .Z(n23791) );
  XOR U24811 ( .A(n23792), .B(n23791), .Z(n23795) );
  NAND U24812 ( .A(b[0]), .B(a[1010]), .Z(n23796) );
  XOR U24813 ( .A(n23795), .B(n23796), .Z(n23798) );
  OR U24814 ( .A(n23772), .B(n23771), .Z(n23776) );
  NANDN U24815 ( .A(n23774), .B(n23773), .Z(n23775) );
  NAND U24816 ( .A(n23776), .B(n23775), .Z(n23797) );
  XNOR U24817 ( .A(n23798), .B(n23797), .Z(n23783) );
  NANDN U24818 ( .A(n23778), .B(n23777), .Z(n23782) );
  OR U24819 ( .A(n23780), .B(n23779), .Z(n23781) );
  NAND U24820 ( .A(n23782), .B(n23781), .Z(n23784) );
  XNOR U24821 ( .A(n23783), .B(n23784), .Z(n23785) );
  XNOR U24822 ( .A(n23786), .B(n23785), .Z(n23801) );
  XNOR U24823 ( .A(n23801), .B(sreg[2030]), .Z(n23802) );
  XOR U24824 ( .A(n23803), .B(n23802), .Z(c[2030]) );
  NANDN U24825 ( .A(n23784), .B(n23783), .Z(n23788) );
  NAND U24826 ( .A(n23786), .B(n23785), .Z(n23787) );
  NAND U24827 ( .A(n23788), .B(n23787), .Z(n23812) );
  AND U24828 ( .A(b[2]), .B(a[1009]), .Z(n23818) );
  AND U24829 ( .A(a[1010]), .B(b[1]), .Z(n23816) );
  AND U24830 ( .A(a[1008]), .B(b[3]), .Z(n23815) );
  XOR U24831 ( .A(n23816), .B(n23815), .Z(n23817) );
  XOR U24832 ( .A(n23818), .B(n23817), .Z(n23821) );
  NAND U24833 ( .A(b[0]), .B(a[1011]), .Z(n23822) );
  XOR U24834 ( .A(n23821), .B(n23822), .Z(n23824) );
  OR U24835 ( .A(n23790), .B(n23789), .Z(n23794) );
  NANDN U24836 ( .A(n23792), .B(n23791), .Z(n23793) );
  NAND U24837 ( .A(n23794), .B(n23793), .Z(n23823) );
  XNOR U24838 ( .A(n23824), .B(n23823), .Z(n23809) );
  NANDN U24839 ( .A(n23796), .B(n23795), .Z(n23800) );
  OR U24840 ( .A(n23798), .B(n23797), .Z(n23799) );
  NAND U24841 ( .A(n23800), .B(n23799), .Z(n23810) );
  XNOR U24842 ( .A(n23809), .B(n23810), .Z(n23811) );
  XNOR U24843 ( .A(n23812), .B(n23811), .Z(n23808) );
  NAND U24844 ( .A(n23801), .B(sreg[2030]), .Z(n23805) );
  OR U24845 ( .A(n23803), .B(n23802), .Z(n23804) );
  AND U24846 ( .A(n23805), .B(n23804), .Z(n23807) );
  XNOR U24847 ( .A(n23807), .B(sreg[2031]), .Z(n23806) );
  XOR U24848 ( .A(n23808), .B(n23806), .Z(c[2031]) );
  NANDN U24849 ( .A(n23810), .B(n23809), .Z(n23814) );
  NAND U24850 ( .A(n23812), .B(n23811), .Z(n23813) );
  NAND U24851 ( .A(n23814), .B(n23813), .Z(n23830) );
  AND U24852 ( .A(b[2]), .B(a[1010]), .Z(n23836) );
  AND U24853 ( .A(a[1011]), .B(b[1]), .Z(n23834) );
  AND U24854 ( .A(a[1009]), .B(b[3]), .Z(n23833) );
  XOR U24855 ( .A(n23834), .B(n23833), .Z(n23835) );
  XOR U24856 ( .A(n23836), .B(n23835), .Z(n23839) );
  NAND U24857 ( .A(b[0]), .B(a[1012]), .Z(n23840) );
  XOR U24858 ( .A(n23839), .B(n23840), .Z(n23842) );
  OR U24859 ( .A(n23816), .B(n23815), .Z(n23820) );
  NANDN U24860 ( .A(n23818), .B(n23817), .Z(n23819) );
  NAND U24861 ( .A(n23820), .B(n23819), .Z(n23841) );
  XNOR U24862 ( .A(n23842), .B(n23841), .Z(n23827) );
  NANDN U24863 ( .A(n23822), .B(n23821), .Z(n23826) );
  OR U24864 ( .A(n23824), .B(n23823), .Z(n23825) );
  NAND U24865 ( .A(n23826), .B(n23825), .Z(n23828) );
  XNOR U24866 ( .A(n23827), .B(n23828), .Z(n23829) );
  XNOR U24867 ( .A(n23830), .B(n23829), .Z(n23845) );
  XNOR U24868 ( .A(n23845), .B(sreg[2032]), .Z(n23847) );
  XNOR U24869 ( .A(n23846), .B(n23847), .Z(c[2032]) );
  NANDN U24870 ( .A(n23828), .B(n23827), .Z(n23832) );
  NAND U24871 ( .A(n23830), .B(n23829), .Z(n23831) );
  NAND U24872 ( .A(n23832), .B(n23831), .Z(n23853) );
  AND U24873 ( .A(b[2]), .B(a[1011]), .Z(n23859) );
  AND U24874 ( .A(a[1012]), .B(b[1]), .Z(n23857) );
  AND U24875 ( .A(a[1010]), .B(b[3]), .Z(n23856) );
  XOR U24876 ( .A(n23857), .B(n23856), .Z(n23858) );
  XOR U24877 ( .A(n23859), .B(n23858), .Z(n23862) );
  NAND U24878 ( .A(b[0]), .B(a[1013]), .Z(n23863) );
  XOR U24879 ( .A(n23862), .B(n23863), .Z(n23865) );
  OR U24880 ( .A(n23834), .B(n23833), .Z(n23838) );
  NANDN U24881 ( .A(n23836), .B(n23835), .Z(n23837) );
  NAND U24882 ( .A(n23838), .B(n23837), .Z(n23864) );
  XNOR U24883 ( .A(n23865), .B(n23864), .Z(n23850) );
  NANDN U24884 ( .A(n23840), .B(n23839), .Z(n23844) );
  OR U24885 ( .A(n23842), .B(n23841), .Z(n23843) );
  NAND U24886 ( .A(n23844), .B(n23843), .Z(n23851) );
  XNOR U24887 ( .A(n23850), .B(n23851), .Z(n23852) );
  XNOR U24888 ( .A(n23853), .B(n23852), .Z(n23868) );
  XNOR U24889 ( .A(n23868), .B(sreg[2033]), .Z(n23870) );
  NAND U24890 ( .A(n23845), .B(sreg[2032]), .Z(n23849) );
  NANDN U24891 ( .A(n23847), .B(n23846), .Z(n23848) );
  AND U24892 ( .A(n23849), .B(n23848), .Z(n23869) );
  XOR U24893 ( .A(n23870), .B(n23869), .Z(c[2033]) );
  NANDN U24894 ( .A(n23851), .B(n23850), .Z(n23855) );
  NAND U24895 ( .A(n23853), .B(n23852), .Z(n23854) );
  NAND U24896 ( .A(n23855), .B(n23854), .Z(n23879) );
  AND U24897 ( .A(b[2]), .B(a[1012]), .Z(n23885) );
  AND U24898 ( .A(a[1013]), .B(b[1]), .Z(n23883) );
  AND U24899 ( .A(a[1011]), .B(b[3]), .Z(n23882) );
  XOR U24900 ( .A(n23883), .B(n23882), .Z(n23884) );
  XOR U24901 ( .A(n23885), .B(n23884), .Z(n23888) );
  NAND U24902 ( .A(b[0]), .B(a[1014]), .Z(n23889) );
  XOR U24903 ( .A(n23888), .B(n23889), .Z(n23891) );
  OR U24904 ( .A(n23857), .B(n23856), .Z(n23861) );
  NANDN U24905 ( .A(n23859), .B(n23858), .Z(n23860) );
  NAND U24906 ( .A(n23861), .B(n23860), .Z(n23890) );
  XNOR U24907 ( .A(n23891), .B(n23890), .Z(n23876) );
  NANDN U24908 ( .A(n23863), .B(n23862), .Z(n23867) );
  OR U24909 ( .A(n23865), .B(n23864), .Z(n23866) );
  NAND U24910 ( .A(n23867), .B(n23866), .Z(n23877) );
  XNOR U24911 ( .A(n23876), .B(n23877), .Z(n23878) );
  XOR U24912 ( .A(n23879), .B(n23878), .Z(n23875) );
  NAND U24913 ( .A(n23868), .B(sreg[2033]), .Z(n23872) );
  OR U24914 ( .A(n23870), .B(n23869), .Z(n23871) );
  NAND U24915 ( .A(n23872), .B(n23871), .Z(n23874) );
  XNOR U24916 ( .A(sreg[2034]), .B(n23874), .Z(n23873) );
  XOR U24917 ( .A(n23875), .B(n23873), .Z(c[2034]) );
  NANDN U24918 ( .A(n23877), .B(n23876), .Z(n23881) );
  NAND U24919 ( .A(n23879), .B(n23878), .Z(n23880) );
  NAND U24920 ( .A(n23881), .B(n23880), .Z(n23897) );
  AND U24921 ( .A(b[2]), .B(a[1013]), .Z(n23903) );
  AND U24922 ( .A(a[1014]), .B(b[1]), .Z(n23901) );
  AND U24923 ( .A(a[1012]), .B(b[3]), .Z(n23900) );
  XOR U24924 ( .A(n23901), .B(n23900), .Z(n23902) );
  XOR U24925 ( .A(n23903), .B(n23902), .Z(n23906) );
  NAND U24926 ( .A(b[0]), .B(a[1015]), .Z(n23907) );
  XOR U24927 ( .A(n23906), .B(n23907), .Z(n23909) );
  OR U24928 ( .A(n23883), .B(n23882), .Z(n23887) );
  NANDN U24929 ( .A(n23885), .B(n23884), .Z(n23886) );
  NAND U24930 ( .A(n23887), .B(n23886), .Z(n23908) );
  XNOR U24931 ( .A(n23909), .B(n23908), .Z(n23894) );
  NANDN U24932 ( .A(n23889), .B(n23888), .Z(n23893) );
  OR U24933 ( .A(n23891), .B(n23890), .Z(n23892) );
  NAND U24934 ( .A(n23893), .B(n23892), .Z(n23895) );
  XNOR U24935 ( .A(n23894), .B(n23895), .Z(n23896) );
  XNOR U24936 ( .A(n23897), .B(n23896), .Z(n23912) );
  XNOR U24937 ( .A(n23912), .B(sreg[2035]), .Z(n23913) );
  XOR U24938 ( .A(n23914), .B(n23913), .Z(c[2035]) );
  NANDN U24939 ( .A(n23895), .B(n23894), .Z(n23899) );
  NAND U24940 ( .A(n23897), .B(n23896), .Z(n23898) );
  NAND U24941 ( .A(n23899), .B(n23898), .Z(n23920) );
  AND U24942 ( .A(b[2]), .B(a[1014]), .Z(n23926) );
  AND U24943 ( .A(a[1015]), .B(b[1]), .Z(n23924) );
  AND U24944 ( .A(a[1013]), .B(b[3]), .Z(n23923) );
  XOR U24945 ( .A(n23924), .B(n23923), .Z(n23925) );
  XOR U24946 ( .A(n23926), .B(n23925), .Z(n23929) );
  NAND U24947 ( .A(b[0]), .B(a[1016]), .Z(n23930) );
  XOR U24948 ( .A(n23929), .B(n23930), .Z(n23932) );
  OR U24949 ( .A(n23901), .B(n23900), .Z(n23905) );
  NANDN U24950 ( .A(n23903), .B(n23902), .Z(n23904) );
  NAND U24951 ( .A(n23905), .B(n23904), .Z(n23931) );
  XNOR U24952 ( .A(n23932), .B(n23931), .Z(n23917) );
  NANDN U24953 ( .A(n23907), .B(n23906), .Z(n23911) );
  OR U24954 ( .A(n23909), .B(n23908), .Z(n23910) );
  NAND U24955 ( .A(n23911), .B(n23910), .Z(n23918) );
  XNOR U24956 ( .A(n23917), .B(n23918), .Z(n23919) );
  XNOR U24957 ( .A(n23920), .B(n23919), .Z(n23935) );
  XNOR U24958 ( .A(n23935), .B(sreg[2036]), .Z(n23937) );
  NAND U24959 ( .A(n23912), .B(sreg[2035]), .Z(n23916) );
  OR U24960 ( .A(n23914), .B(n23913), .Z(n23915) );
  AND U24961 ( .A(n23916), .B(n23915), .Z(n23936) );
  XOR U24962 ( .A(n23937), .B(n23936), .Z(c[2036]) );
  NANDN U24963 ( .A(n23918), .B(n23917), .Z(n23922) );
  NAND U24964 ( .A(n23920), .B(n23919), .Z(n23921) );
  NAND U24965 ( .A(n23922), .B(n23921), .Z(n23948) );
  AND U24966 ( .A(b[2]), .B(a[1015]), .Z(n23954) );
  AND U24967 ( .A(a[1016]), .B(b[1]), .Z(n23952) );
  AND U24968 ( .A(a[1014]), .B(b[3]), .Z(n23951) );
  XOR U24969 ( .A(n23952), .B(n23951), .Z(n23953) );
  XOR U24970 ( .A(n23954), .B(n23953), .Z(n23957) );
  NAND U24971 ( .A(b[0]), .B(a[1017]), .Z(n23958) );
  XOR U24972 ( .A(n23957), .B(n23958), .Z(n23960) );
  OR U24973 ( .A(n23924), .B(n23923), .Z(n23928) );
  NANDN U24974 ( .A(n23926), .B(n23925), .Z(n23927) );
  NAND U24975 ( .A(n23928), .B(n23927), .Z(n23959) );
  XNOR U24976 ( .A(n23960), .B(n23959), .Z(n23945) );
  NANDN U24977 ( .A(n23930), .B(n23929), .Z(n23934) );
  OR U24978 ( .A(n23932), .B(n23931), .Z(n23933) );
  NAND U24979 ( .A(n23934), .B(n23933), .Z(n23946) );
  XNOR U24980 ( .A(n23945), .B(n23946), .Z(n23947) );
  XNOR U24981 ( .A(n23948), .B(n23947), .Z(n23940) );
  XOR U24982 ( .A(sreg[2037]), .B(n23940), .Z(n23941) );
  NAND U24983 ( .A(n23935), .B(sreg[2036]), .Z(n23939) );
  OR U24984 ( .A(n23937), .B(n23936), .Z(n23938) );
  NAND U24985 ( .A(n23939), .B(n23938), .Z(n23942) );
  XOR U24986 ( .A(n23941), .B(n23942), .Z(c[2037]) );
  OR U24987 ( .A(n23940), .B(sreg[2037]), .Z(n23944) );
  NANDN U24988 ( .A(n23942), .B(n23941), .Z(n23943) );
  AND U24989 ( .A(n23944), .B(n23943), .Z(n23964) );
  NANDN U24990 ( .A(n23946), .B(n23945), .Z(n23950) );
  NAND U24991 ( .A(n23948), .B(n23947), .Z(n23949) );
  NAND U24992 ( .A(n23950), .B(n23949), .Z(n23969) );
  AND U24993 ( .A(b[2]), .B(a[1016]), .Z(n23975) );
  AND U24994 ( .A(a[1017]), .B(b[1]), .Z(n23973) );
  AND U24995 ( .A(a[1015]), .B(b[3]), .Z(n23972) );
  XOR U24996 ( .A(n23973), .B(n23972), .Z(n23974) );
  XOR U24997 ( .A(n23975), .B(n23974), .Z(n23978) );
  NAND U24998 ( .A(b[0]), .B(a[1018]), .Z(n23979) );
  XOR U24999 ( .A(n23978), .B(n23979), .Z(n23981) );
  OR U25000 ( .A(n23952), .B(n23951), .Z(n23956) );
  NANDN U25001 ( .A(n23954), .B(n23953), .Z(n23955) );
  NAND U25002 ( .A(n23956), .B(n23955), .Z(n23980) );
  XNOR U25003 ( .A(n23981), .B(n23980), .Z(n23966) );
  NANDN U25004 ( .A(n23958), .B(n23957), .Z(n23962) );
  OR U25005 ( .A(n23960), .B(n23959), .Z(n23961) );
  NAND U25006 ( .A(n23962), .B(n23961), .Z(n23967) );
  XNOR U25007 ( .A(n23966), .B(n23967), .Z(n23968) );
  XNOR U25008 ( .A(n23969), .B(n23968), .Z(n23965) );
  XOR U25009 ( .A(sreg[2038]), .B(n23965), .Z(n23963) );
  XOR U25010 ( .A(n23964), .B(n23963), .Z(c[2038]) );
  NANDN U25011 ( .A(n23967), .B(n23966), .Z(n23971) );
  NAND U25012 ( .A(n23969), .B(n23968), .Z(n23970) );
  NAND U25013 ( .A(n23971), .B(n23970), .Z(n23992) );
  AND U25014 ( .A(b[2]), .B(a[1017]), .Z(n23998) );
  AND U25015 ( .A(a[1018]), .B(b[1]), .Z(n23996) );
  AND U25016 ( .A(a[1016]), .B(b[3]), .Z(n23995) );
  XOR U25017 ( .A(n23996), .B(n23995), .Z(n23997) );
  XOR U25018 ( .A(n23998), .B(n23997), .Z(n24001) );
  NAND U25019 ( .A(b[0]), .B(a[1019]), .Z(n24002) );
  XOR U25020 ( .A(n24001), .B(n24002), .Z(n24004) );
  OR U25021 ( .A(n23973), .B(n23972), .Z(n23977) );
  NANDN U25022 ( .A(n23975), .B(n23974), .Z(n23976) );
  NAND U25023 ( .A(n23977), .B(n23976), .Z(n24003) );
  XNOR U25024 ( .A(n24004), .B(n24003), .Z(n23989) );
  NANDN U25025 ( .A(n23979), .B(n23978), .Z(n23983) );
  OR U25026 ( .A(n23981), .B(n23980), .Z(n23982) );
  NAND U25027 ( .A(n23983), .B(n23982), .Z(n23990) );
  XNOR U25028 ( .A(n23989), .B(n23990), .Z(n23991) );
  XNOR U25029 ( .A(n23992), .B(n23991), .Z(n23984) );
  XNOR U25030 ( .A(n23984), .B(sreg[2039]), .Z(n23986) );
  XNOR U25031 ( .A(n23985), .B(n23986), .Z(c[2039]) );
  NAND U25032 ( .A(n23984), .B(sreg[2039]), .Z(n23988) );
  NANDN U25033 ( .A(n23986), .B(n23985), .Z(n23987) );
  NAND U25034 ( .A(n23988), .B(n23987), .Z(n24009) );
  NANDN U25035 ( .A(n23990), .B(n23989), .Z(n23994) );
  NAND U25036 ( .A(n23992), .B(n23991), .Z(n23993) );
  NAND U25037 ( .A(n23994), .B(n23993), .Z(n24015) );
  AND U25038 ( .A(b[2]), .B(a[1018]), .Z(n24021) );
  AND U25039 ( .A(a[1019]), .B(b[1]), .Z(n24019) );
  AND U25040 ( .A(a[1017]), .B(b[3]), .Z(n24018) );
  XOR U25041 ( .A(n24019), .B(n24018), .Z(n24020) );
  XOR U25042 ( .A(n24021), .B(n24020), .Z(n24024) );
  NAND U25043 ( .A(b[0]), .B(a[1020]), .Z(n24025) );
  XOR U25044 ( .A(n24024), .B(n24025), .Z(n24027) );
  OR U25045 ( .A(n23996), .B(n23995), .Z(n24000) );
  NANDN U25046 ( .A(n23998), .B(n23997), .Z(n23999) );
  NAND U25047 ( .A(n24000), .B(n23999), .Z(n24026) );
  XNOR U25048 ( .A(n24027), .B(n24026), .Z(n24012) );
  NANDN U25049 ( .A(n24002), .B(n24001), .Z(n24006) );
  OR U25050 ( .A(n24004), .B(n24003), .Z(n24005) );
  NAND U25051 ( .A(n24006), .B(n24005), .Z(n24013) );
  XNOR U25052 ( .A(n24012), .B(n24013), .Z(n24014) );
  XNOR U25053 ( .A(n24015), .B(n24014), .Z(n24007) );
  XOR U25054 ( .A(sreg[2040]), .B(n24007), .Z(n24008) );
  XOR U25055 ( .A(n24009), .B(n24008), .Z(c[2040]) );
  OR U25056 ( .A(n24007), .B(sreg[2040]), .Z(n24011) );
  NANDN U25057 ( .A(n24009), .B(n24008), .Z(n24010) );
  AND U25058 ( .A(n24011), .B(n24010), .Z(n24031) );
  NANDN U25059 ( .A(n24013), .B(n24012), .Z(n24017) );
  NAND U25060 ( .A(n24015), .B(n24014), .Z(n24016) );
  NAND U25061 ( .A(n24017), .B(n24016), .Z(n24036) );
  AND U25062 ( .A(b[2]), .B(a[1019]), .Z(n24041) );
  AND U25063 ( .A(a[1020]), .B(b[1]), .Z(n24079) );
  ANDN U25064 ( .B(a[1018]), .A(n1796), .Z(n24039) );
  XOR U25065 ( .A(n24079), .B(n24039), .Z(n24040) );
  XOR U25066 ( .A(n24041), .B(n24040), .Z(n24042) );
  NAND U25067 ( .A(a[1021]), .B(b[0]), .Z(n24043) );
  XNOR U25068 ( .A(n24042), .B(n24043), .Z(n24044) );
  OR U25069 ( .A(n24019), .B(n24018), .Z(n24023) );
  NANDN U25070 ( .A(n24021), .B(n24020), .Z(n24022) );
  NAND U25071 ( .A(n24023), .B(n24022), .Z(n24045) );
  XOR U25072 ( .A(n24044), .B(n24045), .Z(n24033) );
  NANDN U25073 ( .A(n24025), .B(n24024), .Z(n24029) );
  OR U25074 ( .A(n24027), .B(n24026), .Z(n24028) );
  NAND U25075 ( .A(n24029), .B(n24028), .Z(n24034) );
  XNOR U25076 ( .A(n24033), .B(n24034), .Z(n24035) );
  XNOR U25077 ( .A(n24036), .B(n24035), .Z(n24032) );
  XOR U25078 ( .A(sreg[2041]), .B(n24032), .Z(n24030) );
  XOR U25079 ( .A(n24031), .B(n24030), .Z(c[2041]) );
  NANDN U25080 ( .A(n24034), .B(n24033), .Z(n24038) );
  NAND U25081 ( .A(n24036), .B(n24035), .Z(n24037) );
  NAND U25082 ( .A(n24038), .B(n24037), .Z(n24056) );
  AND U25083 ( .A(b[2]), .B(a[1020]), .Z(n24060) );
  NANDN U25084 ( .A(n1796), .B(a[1019]), .Z(n24058) );
  XNOR U25085 ( .A(n24059), .B(n24058), .Z(n24061) );
  XOR U25086 ( .A(n24060), .B(n24061), .Z(n24064) );
  NAND U25087 ( .A(b[0]), .B(a[1022]), .Z(n24065) );
  XOR U25088 ( .A(n24064), .B(n24065), .Z(n24066) );
  XOR U25089 ( .A(n24066), .B(n24067), .Z(n24053) );
  NANDN U25090 ( .A(n24043), .B(n24042), .Z(n24047) );
  NANDN U25091 ( .A(n24045), .B(n24044), .Z(n24046) );
  AND U25092 ( .A(n24047), .B(n24046), .Z(n24054) );
  XOR U25093 ( .A(n24053), .B(n24054), .Z(n24055) );
  XOR U25094 ( .A(n24056), .B(n24055), .Z(n24048) );
  XNOR U25095 ( .A(n24048), .B(sreg[2042]), .Z(n24050) );
  XNOR U25096 ( .A(n24049), .B(n24050), .Z(c[2042]) );
  NAND U25097 ( .A(n24048), .B(sreg[2042]), .Z(n24052) );
  NANDN U25098 ( .A(n24050), .B(n24049), .Z(n24051) );
  NAND U25099 ( .A(n24052), .B(n24051), .Z(n24068) );
  XNOR U25100 ( .A(n24068), .B(sreg[2043]), .Z(n24070) );
  AND U25101 ( .A(a[1020]), .B(b[3]), .Z(n24057) );
  NAND U25102 ( .A(b[1]), .B(a[1022]), .Z(n24100) );
  XOR U25103 ( .A(n24057), .B(n24100), .Z(n24081) );
  NAND U25104 ( .A(a[1021]), .B(b[2]), .Z(n24080) );
  XOR U25105 ( .A(n24081), .B(n24080), .Z(n24084) );
  NAND U25106 ( .A(b[0]), .B(a[1023]), .Z(n24085) );
  XOR U25107 ( .A(n24084), .B(n24085), .Z(n24086) );
  NAND U25108 ( .A(n24059), .B(n24058), .Z(n24063) );
  OR U25109 ( .A(n24061), .B(n24060), .Z(n24062) );
  AND U25110 ( .A(n24063), .B(n24062), .Z(n24087) );
  XNOR U25111 ( .A(n24086), .B(n24087), .Z(n24074) );
  XNOR U25112 ( .A(n24074), .B(n24073), .Z(n24076) );
  XOR U25113 ( .A(n24075), .B(n24076), .Z(n24069) );
  XOR U25114 ( .A(n24070), .B(n24069), .Z(c[2043]) );
  NAND U25115 ( .A(n24068), .B(sreg[2043]), .Z(n24072) );
  OR U25116 ( .A(n24070), .B(n24069), .Z(n24071) );
  AND U25117 ( .A(n24072), .B(n24071), .Z(n24089) );
  NANDN U25118 ( .A(n24074), .B(n24073), .Z(n24078) );
  NAND U25119 ( .A(n24076), .B(n24075), .Z(n24077) );
  NAND U25120 ( .A(n24078), .B(n24077), .Z(n24092) );
  AND U25121 ( .A(a[1022]), .B(b[3]), .Z(n24110) );
  NAND U25122 ( .A(n24079), .B(n24110), .Z(n24083) );
  OR U25123 ( .A(n24081), .B(n24080), .Z(n24082) );
  NAND U25124 ( .A(n24083), .B(n24082), .Z(n24099) );
  NAND U25125 ( .A(b[1]), .B(a[1023]), .Z(n24109) );
  AND U25126 ( .A(b[2]), .B(a[1022]), .Z(n24108) );
  XNOR U25127 ( .A(n24109), .B(n24108), .Z(n24096) );
  NAND U25128 ( .A(a[1021]), .B(b[3]), .Z(n24097) );
  XOR U25129 ( .A(n24096), .B(n24097), .Z(n24098) );
  XNOR U25130 ( .A(n24099), .B(n24098), .Z(n24091) );
  XNOR U25131 ( .A(n24091), .B(n24090), .Z(n24093) );
  XOR U25132 ( .A(n24092), .B(n24093), .Z(n24088) );
  XOR U25133 ( .A(n24089), .B(n24088), .Z(c[2044]) );
  OR U25134 ( .A(n24089), .B(n24088), .Z(n24114) );
  NANDN U25135 ( .A(n24091), .B(n24090), .Z(n24095) );
  NAND U25136 ( .A(n24093), .B(n24092), .Z(n24094) );
  NAND U25137 ( .A(n24095), .B(n24094), .Z(n24105) );
  AND U25138 ( .A(n24100), .B(b[2]), .Z(n24101) );
  NAND U25139 ( .A(n24101), .B(a[1023]), .Z(n24111) );
  XNOR U25140 ( .A(n24110), .B(n24111), .Z(n24103) );
  XOR U25141 ( .A(n24102), .B(n24103), .Z(n24104) );
  XOR U25142 ( .A(n24105), .B(n24104), .Z(n24115) );
  XOR U25143 ( .A(n24114), .B(n24115), .Z(c[2045]) );
  NAND U25144 ( .A(n24103), .B(n24102), .Z(n24107) );
  NANDN U25145 ( .A(n24105), .B(n24104), .Z(n24106) );
  NAND U25146 ( .A(n24107), .B(n24106), .Z(n24122) );
  NAND U25147 ( .A(b[3]), .B(a[1023]), .Z(n24119) );
  XOR U25148 ( .A(n24122), .B(n24119), .Z(n24117) );
  NANDN U25149 ( .A(n24109), .B(n24108), .Z(n24113) );
  NANDN U25150 ( .A(n24111), .B(n24110), .Z(n24112) );
  NAND U25151 ( .A(n24113), .B(n24112), .Z(n24120) );
  NOR U25152 ( .A(n24115), .B(n24114), .Z(n24121) );
  XOR U25153 ( .A(n24120), .B(n24121), .Z(n24116) );
  XNOR U25154 ( .A(n24117), .B(n24116), .Z(c[2046]) );
  XNOR U25155 ( .A(n24121), .B(n24120), .Z(n24123) );
  XNOR U25156 ( .A(n24122), .B(n24123), .Z(n24118) );
  NANDN U25157 ( .A(n24119), .B(n24118), .Z(n24127) );
  OR U25158 ( .A(n24121), .B(n24120), .Z(n24125) );
  OR U25159 ( .A(n24123), .B(n24122), .Z(n24124) );
  NAND U25160 ( .A(n24125), .B(n24124), .Z(n24126) );
  NAND U25161 ( .A(n24127), .B(n24126), .Z(c[2047]) );
endmodule

